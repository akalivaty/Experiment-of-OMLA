//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0010(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0011(.A1(new_n206), .A2(new_n207), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT66), .Z(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR3_X1   g0018(.A1(new_n217), .A2(new_n218), .A3(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n213), .A2(new_n215), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n203), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n225), .B(new_n230), .C1(G58), .C2(G232), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(G1), .B2(G20), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT1), .Z(new_n233));
  AOI211_X1 g0033(.A(new_n221), .B(new_n233), .C1(new_n216), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  INV_X1    g0038(.A(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n224), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G107), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n223), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  AND2_X1   g0053(.A1(KEYINPUT77), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(KEYINPUT77), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT3), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n229), .A2(G1698), .ZN(new_n259));
  OR2_X1    g0059(.A1(G250), .A2(G1698), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n256), .A2(new_n258), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n254), .A2(new_n255), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G294), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n265), .B1(G33), .B2(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT5), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n217), .B(G45), .C1(new_n268), .C2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT68), .A2(G41), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT68), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(new_n273), .A3(G274), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n266), .B1(new_n270), .B2(new_n273), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G264), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n267), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G200), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n261), .B2(new_n263), .ZN(new_n282));
  INV_X1    g0082(.A(G264), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n283), .B(new_n266), .C1(new_n270), .C2(new_n273), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G190), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(new_n274), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT22), .ZN(new_n290));
  INV_X1    g0090(.A(G87), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n290), .A2(new_n291), .A3(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n256), .A2(new_n258), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n291), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT3), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n258), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n290), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n262), .A2(new_n218), .A3(G116), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n218), .B2(G107), .ZN(new_n301));
  INV_X1    g0101(.A(G107), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT23), .A3(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n293), .A2(new_n298), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT88), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n254), .A2(new_n255), .A3(new_n223), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n218), .A2(new_n307), .B1(new_n297), .B2(new_n290), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT88), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n304), .A4(new_n293), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n310), .A3(KEYINPUT24), .ZN(new_n311));
  NAND3_X1  g0111(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n265), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT24), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n305), .A2(KEYINPUT88), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n313), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(G1), .C2(new_n295), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT25), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n318), .B2(G107), .ZN(new_n322));
  INV_X1    g0122(.A(new_n318), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n302), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n320), .A2(G107), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT89), .B1(new_n289), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT89), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n288), .A2(new_n328), .A3(new_n316), .A4(new_n325), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n218), .A2(G33), .A3(G77), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n218), .A2(new_n295), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n332), .B1(new_n218), .B2(G68), .C1(new_n333), .C2(new_n207), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n313), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT11), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n323), .A2(new_n203), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n317), .A2(KEYINPUT70), .A3(new_n318), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n323), .B2(new_n313), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G1), .B2(new_n218), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n336), .B(new_n338), .C1(new_n203), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n343), .A2(new_n203), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(new_n338), .A4(new_n336), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT3), .B(G33), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G226), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n258), .A2(new_n296), .A3(G232), .A4(G1698), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n266), .ZN(new_n357));
  INV_X1    g0157(.A(G45), .ZN(new_n358));
  AND2_X1   g0158(.A1(KEYINPUT68), .A2(G41), .ZN(new_n359));
  NOR2_X1   g0159(.A1(KEYINPUT68), .A2(G41), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n217), .A3(G274), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n281), .A2(G238), .A3(new_n363), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n362), .A2(KEYINPUT72), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT72), .B1(new_n362), .B2(new_n364), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n357), .B(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n350), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT14), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(KEYINPUT74), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n362), .A2(new_n364), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n362), .A2(KEYINPUT72), .A3(new_n364), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n369), .A4(new_n357), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n367), .B2(KEYINPUT13), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n367), .A2(new_n382), .A3(KEYINPUT13), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n381), .B(G179), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n349), .B1(new_n372), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n381), .B(G190), .C1(new_n383), .C2(new_n384), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n369), .B1(new_n378), .B2(new_n357), .ZN(new_n388));
  INV_X1    g0188(.A(new_n370), .ZN(new_n389));
  OAI21_X1  g0189(.A(G200), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n387), .A2(new_n349), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n331), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(G169), .B1(new_n388), .B2(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT14), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n371), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n385), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n349), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n387), .A2(new_n349), .A3(new_n390), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n351), .A2(G222), .A3(new_n352), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n351), .A2(G1698), .ZN(new_n404));
  INV_X1    g0204(.A(G223), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n403), .B1(new_n251), .B2(new_n351), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n266), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n281), .A2(new_n363), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n362), .C1(new_n239), .C2(new_n408), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n409), .A2(G179), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT8), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G58), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n218), .B(G33), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n208), .A2(G20), .ZN(new_n418));
  INV_X1    g0218(.A(new_n333), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G150), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n313), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n318), .A2(G50), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n313), .B1(new_n217), .B2(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G50), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n409), .A2(new_n350), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n410), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n404), .A2(new_n227), .B1(new_n302), .B2(new_n351), .ZN(new_n430));
  INV_X1    g0230(.A(new_n351), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n431), .A2(new_n236), .A3(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n266), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G244), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n433), .B(new_n362), .C1(new_n434), .C2(new_n408), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n323), .A2(new_n251), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G20), .A2(G77), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT15), .B(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n218), .A2(G33), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n411), .A2(new_n413), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n438), .B1(new_n439), .B2(new_n440), .C1(new_n441), .C2(new_n333), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n313), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n437), .B(new_n443), .C1(new_n343), .C2(new_n251), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n435), .A2(new_n350), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n436), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT9), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT71), .ZN(new_n449));
  AND4_X1   g0249(.A1(new_n449), .A2(new_n422), .A3(new_n424), .A4(new_n426), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n423), .B1(new_n421), .B2(new_n313), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(new_n426), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n448), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n449), .A3(new_n426), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(KEYINPUT9), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n409), .A2(new_n286), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n409), .A2(G200), .ZN(new_n459));
  AND4_X1   g0259(.A1(new_n447), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n459), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n453), .B2(new_n456), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n447), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n429), .B(new_n446), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n281), .A2(G232), .A3(new_n363), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n362), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT81), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n362), .A2(KEYINPUT81), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G87), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT80), .Z(new_n472));
  NAND2_X1  g0272(.A1(new_n405), .A2(new_n352), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n256), .A2(new_n258), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n352), .A2(G226), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n266), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n286), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n468), .A2(new_n469), .B1(new_n476), .B2(new_n266), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(G200), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n415), .A2(new_n416), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n425), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n318), .B2(new_n481), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n257), .B1(new_n254), .B2(new_n255), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(KEYINPUT7), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT79), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n485), .A2(new_n489), .A3(KEYINPUT7), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT7), .B1(new_n431), .B2(new_n218), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G68), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n202), .A2(new_n203), .ZN(new_n496));
  OAI21_X1  g0296(.A(G20), .B1(new_n206), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n419), .A2(G159), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT16), .B1(new_n495), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g0301(.A1(KEYINPUT77), .A2(G33), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT77), .A2(G33), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n257), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n258), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT78), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT78), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n256), .A2(new_n507), .A3(new_n258), .ZN(new_n508));
  NOR2_X1   g0308(.A1(KEYINPUT7), .A2(G20), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(G20), .B1(new_n256), .B2(new_n258), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT7), .ZN(new_n512));
  OAI21_X1  g0312(.A(G68), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(KEYINPUT16), .B(new_n500), .C1(new_n510), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n313), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n480), .B(new_n484), .C1(new_n501), .C2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT17), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(KEYINPUT82), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(KEYINPUT82), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n492), .B1(new_n488), .B2(new_n490), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n500), .B1(new_n522), .B2(new_n203), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT16), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n218), .B1(new_n504), .B2(new_n505), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n203), .B1(new_n526), .B2(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n499), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n317), .B1(new_n529), .B2(KEYINPUT16), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n483), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n521), .B1(new_n531), .B2(new_n480), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n519), .B1(new_n532), .B2(new_n518), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n484), .B1(new_n501), .B2(new_n515), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n470), .A2(G179), .A3(new_n477), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n350), .B1(new_n470), .B2(new_n477), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n534), .A2(new_n538), .A3(KEYINPUT18), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT18), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n531), .B2(new_n537), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n435), .A2(new_n286), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n444), .B1(G200), .B2(new_n435), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n533), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n402), .A2(new_n464), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(KEYINPUT6), .A2(G97), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT83), .B1(new_n548), .B2(G107), .ZN(new_n549));
  OR3_X1    g0349(.A1(new_n548), .A2(KEYINPUT83), .A3(G107), .ZN(new_n550));
  XOR2_X1   g0350(.A(G97), .B(G107), .Z(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(KEYINPUT6), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n419), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n522), .B2(new_n302), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n313), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n318), .A2(G97), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n556), .B1(new_n320), .B2(G97), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n258), .A2(new_n296), .A3(G250), .A4(G1698), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G283), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(KEYINPUT4), .A2(G244), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n258), .A2(new_n296), .A3(new_n561), .A4(new_n352), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT84), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT84), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n351), .A2(new_n564), .A3(new_n352), .A4(new_n561), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n256), .A2(G244), .A3(new_n352), .A4(new_n258), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n281), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n275), .A2(G257), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n274), .ZN(new_n572));
  OAI21_X1  g0372(.A(G200), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n555), .A2(new_n557), .A3(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n560), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n563), .A2(new_n565), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n266), .ZN(new_n578));
  INV_X1    g0378(.A(new_n572), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT85), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n570), .A2(new_n581), .A3(new_n572), .ZN(new_n582));
  OAI21_X1  g0382(.A(G190), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n570), .A2(G179), .A3(new_n572), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n555), .B2(new_n557), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n581), .B1(new_n570), .B2(new_n572), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n578), .A2(KEYINPUT85), .A3(new_n579), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n350), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(new_n218), .A3(G33), .A4(G97), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n291), .B1(new_n354), .B2(new_n218), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n591), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n256), .A2(new_n218), .A3(G68), .A4(new_n258), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n317), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n319), .A2(new_n439), .ZN(new_n598));
  INV_X1    g0398(.A(new_n439), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n318), .ZN(new_n600));
  OR3_X1    g0400(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n227), .A2(new_n352), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n434), .A2(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n256), .A2(new_n258), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n307), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n266), .ZN(new_n607));
  INV_X1    g0407(.A(G179), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n217), .A2(G45), .ZN(new_n609));
  INV_X1    g0409(.A(G274), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n281), .A2(G250), .A3(new_n609), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n607), .A2(new_n608), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n607), .A2(new_n612), .A3(new_n613), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n601), .B(new_n614), .C1(new_n615), .C2(G169), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n319), .A2(new_n291), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n597), .A2(new_n617), .A3(new_n600), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n607), .A2(G190), .A3(new_n612), .A4(new_n613), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n615), .C2(new_n278), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n584), .A2(new_n590), .A3(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n312), .A2(new_n265), .B1(G20), .B2(new_n223), .ZN(new_n623));
  AOI21_X1  g0423(.A(G20), .B1(G33), .B2(G283), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n295), .A2(G97), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT87), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT87), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(KEYINPUT20), .B(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n223), .B1(new_n217), .B2(G33), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n342), .A2(new_n633), .B1(new_n223), .B2(new_n323), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n350), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT5), .ZN(new_n636));
  OAI211_X1 g0436(.A(G270), .B(new_n281), .C1(new_n636), .C2(new_n269), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n274), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT86), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n283), .A2(G1698), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n229), .A2(new_n352), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n256), .A2(new_n258), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G303), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n642), .B1(new_n643), .B2(new_n351), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n266), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT86), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n274), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n639), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n635), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n647), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n637), .B2(new_n274), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n632), .A2(new_n634), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(G179), .A4(new_n645), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n635), .A2(KEYINPUT21), .A3(new_n648), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n651), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n274), .ZN(new_n659));
  NOR4_X1   g0459(.A1(new_n282), .A2(new_n284), .A3(new_n659), .A4(G179), .ZN(new_n660));
  AOI21_X1  g0460(.A(G169), .B1(new_n285), .B2(new_n274), .ZN(new_n661));
  AOI211_X1 g0461(.A(new_n660), .B(new_n661), .C1(new_n316), .C2(new_n325), .ZN(new_n662));
  INV_X1    g0462(.A(new_n655), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n639), .A2(new_n645), .A3(G190), .A4(new_n647), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n639), .A2(new_n645), .A3(new_n647), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n278), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n658), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n330), .A2(new_n547), .A3(new_n622), .A4(new_n668), .ZN(G372));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n656), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT21), .B1(new_n635), .B2(new_n648), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT90), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n661), .B1(new_n316), .B2(new_n325), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(G179), .B2(new_n277), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n651), .A2(new_n675), .A3(new_n656), .A4(new_n657), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n622), .A2(new_n330), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n616), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n616), .A2(new_n620), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n590), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n621), .A2(KEYINPUT26), .A3(new_n589), .A4(new_n586), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n547), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n429), .ZN(new_n687));
  INV_X1    g0487(.A(new_n446), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n533), .B(new_n400), .C1(new_n386), .C2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n542), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n460), .A2(new_n463), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(G330), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n672), .A2(new_n676), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n217), .A2(new_n218), .A3(G13), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(KEYINPUT91), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n698), .A2(G213), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n663), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n695), .A2(new_n705), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n658), .A2(new_n667), .A3(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n706), .A2(new_n710), .A3(new_n707), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n694), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n662), .A2(new_n704), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n327), .A2(new_n329), .B1(new_n326), .B2(new_n703), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n662), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n658), .A3(new_n674), .A4(new_n704), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n713), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n219), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n359), .A2(new_n360), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n593), .A2(new_n291), .A3(new_n223), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n724), .A2(new_n217), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  INV_X1    g0529(.A(new_n724), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(new_n729), .C1(new_n213), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT28), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n584), .A2(new_n590), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  INV_X1    g0535(.A(new_n658), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n674), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT96), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n584), .A2(new_n590), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n681), .B1(new_n327), .B2(new_n329), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n735), .A2(new_n737), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n684), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n733), .B1(new_n742), .B2(new_n704), .ZN(new_n743));
  AOI211_X1 g0543(.A(KEYINPUT29), .B(new_n703), .C1(new_n678), .C2(new_n684), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n580), .A2(new_n582), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n665), .A2(G179), .A3(new_n285), .A4(new_n615), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n277), .B1(new_n570), .B2(new_n572), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT94), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n615), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n277), .B(KEYINPUT94), .C1(new_n570), .C2(new_n572), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n752), .A2(new_n608), .A3(new_n648), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n587), .A2(new_n588), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n615), .A2(new_n285), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n648), .A2(new_n608), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT30), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n749), .A2(new_n754), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n703), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT95), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n622), .A2(new_n668), .A3(new_n330), .A4(new_n704), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n759), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(KEYINPUT95), .A3(new_n761), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G330), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n745), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n732), .B1(new_n770), .B2(G1), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT97), .Z(G364));
  INV_X1    g0572(.A(G13), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n217), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n724), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n712), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n709), .A2(new_n711), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(G330), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n506), .A2(new_n508), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n722), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n212), .A2(new_n358), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n783), .C1(new_n252), .C2(new_n358), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n351), .A2(new_n219), .A3(G355), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(G116), .C2(new_n219), .ZN(new_n786));
  OR3_X1    g0586(.A1(KEYINPUT98), .A2(G13), .A3(G33), .ZN(new_n787));
  OAI21_X1  g0587(.A(KEYINPUT98), .B1(G13), .B2(G33), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n265), .B1(G20), .B2(new_n350), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n777), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n218), .A2(new_n608), .A3(new_n278), .A4(G190), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n351), .B1(new_n797), .B2(new_n203), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n218), .A2(new_n608), .A3(new_n286), .A4(new_n278), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n218), .B1(new_n801), .B2(G190), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n800), .A2(new_n207), .B1(new_n802), .B2(new_n228), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n218), .A2(new_n286), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n608), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n798), .B(new_n803), .C1(G58), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n218), .A2(G190), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n805), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G77), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n801), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G159), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT32), .Z(new_n815));
  NOR2_X1   g0615(.A1(new_n278), .A2(G179), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n809), .A2(new_n816), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G87), .A2(new_n818), .B1(new_n820), .B2(G107), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n808), .A2(new_n811), .A3(new_n815), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT99), .Z(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n802), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n351), .B1(new_n799), .B2(G326), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n819), .ZN(new_n828));
  XNOR2_X1  g0628(.A(KEYINPUT33), .B(G317), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n825), .B(new_n828), .C1(new_n796), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n810), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  INV_X1    g0632(.A(G329), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n831), .A2(new_n832), .B1(new_n812), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n817), .B(KEYINPUT100), .Z(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(G303), .ZN(new_n837));
  INV_X1    g0637(.A(G322), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n830), .B(new_n837), .C1(new_n838), .C2(new_n806), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n823), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n795), .B1(new_n840), .B2(new_n792), .ZN(new_n841));
  INV_X1    g0641(.A(new_n791), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n794), .B(new_n841), .C1(new_n779), .C2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n780), .A2(new_n843), .ZN(G396));
  NAND2_X1  g0644(.A1(new_n685), .A2(new_n704), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n446), .A2(new_n703), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n444), .A2(new_n703), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n545), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n446), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n851), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n685), .A2(new_n704), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n852), .A2(new_n768), .A3(G330), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n795), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n855), .A2(new_n858), .A3(new_n795), .ZN(new_n859));
  INV_X1    g0659(.A(new_n769), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n852), .A2(new_n854), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n857), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n431), .B1(new_n819), .B2(new_n291), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n800), .A2(new_n643), .B1(new_n802), .B2(new_n228), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n863), .B(new_n864), .C1(G294), .C2(new_n807), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n813), .A2(G311), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G283), .A2(new_n796), .B1(new_n810), .B2(G116), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT101), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n836), .A2(G107), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n865), .A2(new_n866), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n799), .A2(G137), .B1(new_n810), .B2(G159), .ZN(new_n871));
  INV_X1    g0671(.A(G143), .ZN(new_n872));
  INV_X1    g0672(.A(G150), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n871), .B1(new_n872), .B2(new_n806), .C1(new_n873), .C2(new_n797), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT34), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n802), .A2(new_n202), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n819), .A2(new_n203), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(new_n836), .C2(G50), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n875), .A2(new_n781), .A3(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(G132), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n812), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n870), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n795), .B1(new_n882), .B2(new_n792), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n789), .A2(new_n792), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n251), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n883), .B(new_n885), .C1(new_n853), .C2(new_n790), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n862), .A2(new_n886), .ZN(G384));
  AOI21_X1  g0687(.A(new_n518), .B1(new_n516), .B2(new_n520), .ZN(new_n888));
  INV_X1    g0688(.A(new_n518), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n531), .B2(new_n480), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT18), .B1(new_n534), .B2(new_n538), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n531), .A2(new_n540), .A3(new_n537), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n888), .A2(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n529), .A2(KEYINPUT16), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n483), .B1(new_n895), .B2(new_n530), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n701), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n484), .B1(new_n515), .B2(new_n894), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n470), .A2(G179), .A3(new_n477), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n701), .C1(new_n350), .C2(new_n479), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n531), .A2(new_n480), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n902), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n516), .B1(new_n896), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(KEYINPUT103), .A3(KEYINPUT37), .ZN(new_n908));
  INV_X1    g0708(.A(new_n701), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n534), .B1(new_n538), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n516), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n905), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n898), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n898), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n398), .B(new_n703), .C1(new_n391), .C2(new_n397), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n398), .A2(new_n703), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n399), .A2(new_n400), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n851), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT40), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n910), .A2(new_n516), .A3(new_n912), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n912), .B1(new_n910), .B2(new_n516), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n534), .A2(new_n909), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n533), .B2(new_n542), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n916), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n918), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n925), .A2(KEYINPUT40), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n926), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n547), .A2(new_n920), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(G330), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n547), .B1(new_n743), .B2(new_n744), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n692), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n938), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n399), .A2(new_n703), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n917), .B2(new_n918), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n932), .A2(new_n918), .A3(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n542), .A2(new_n909), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n921), .A2(new_n923), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n854), .B2(new_n847), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n947), .B1(new_n950), .B2(new_n919), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n941), .B(new_n952), .Z(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n217), .B2(new_n774), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n223), .B1(new_n552), .B2(KEYINPUT35), .ZN(new_n955));
  INV_X1    g0755(.A(new_n215), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n955), .B(new_n956), .C1(KEYINPUT35), .C2(new_n552), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  OAI21_X1  g0758(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n213), .A2(new_n959), .B1(G50), .B2(new_n203), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n773), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT105), .ZN(G367));
  AND2_X1   g0763(.A1(new_n555), .A2(new_n557), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n735), .B(new_n739), .C1(new_n964), .C2(new_n704), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n586), .A2(new_n589), .A3(new_n703), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(KEYINPUT42), .B1(new_n967), .B2(new_n718), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  INV_X1    g0770(.A(new_n718), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n590), .B1(new_n965), .B2(new_n674), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n704), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT109), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n704), .A2(new_n618), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n621), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n616), .A2(new_n978), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n979), .A2(KEYINPUT106), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT106), .B1(new_n979), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n712), .A2(new_n716), .A3(new_n969), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n986));
  NAND3_X1  g0786(.A1(new_n981), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT108), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n985), .A2(new_n988), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n977), .A2(new_n984), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n977), .A2(new_n984), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n724), .B(KEYINPUT41), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n967), .B2(new_n719), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n720), .A2(new_n969), .A3(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n967), .A2(new_n719), .A3(KEYINPUT44), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n720), .B2(new_n969), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n716), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n715), .B1(new_n736), .B2(new_n703), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n718), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n712), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n712), .A2(new_n1010), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1008), .A2(new_n770), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n996), .B1(new_n1015), .B2(new_n770), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n991), .B(new_n994), .C1(new_n1016), .C2(new_n776), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n781), .B1(G97), .B2(new_n820), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n812), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT111), .Z(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n835), .A2(new_n1022), .A3(new_n223), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1022), .B1(new_n817), .B2(new_n223), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n302), .B2(new_n802), .C1(new_n800), .C2(new_n832), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n797), .A2(new_n824), .B1(new_n831), .B2(new_n827), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1021), .B(new_n1027), .C1(new_n643), .C2(new_n806), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G58), .A2(new_n818), .B1(new_n820), .B2(G77), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n873), .B2(new_n806), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G143), .A2(new_n799), .B1(new_n796), .B2(G159), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n203), .B2(new_n802), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n351), .B1(new_n831), .B2(new_n207), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(G137), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(new_n812), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT47), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n795), .B1(new_n1038), .B2(new_n792), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n782), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n793), .B1(new_n219), .B2(new_n439), .C1(new_n243), .C2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n981), .A2(new_n791), .A3(new_n982), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1017), .A2(new_n1043), .ZN(G387));
  NOR2_X1   g0844(.A1(new_n716), .A2(new_n842), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n351), .A2(new_n219), .A3(new_n725), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n441), .A2(G50), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  INV_X1    g0848(.A(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(G45), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n725), .B1(G68), .B2(G77), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n1049), .C2(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n782), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n240), .A2(new_n358), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1046), .B1(G107), .B2(new_n219), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n793), .B1(new_n1055), .B2(KEYINPUT113), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(KEYINPUT113), .B2(new_n1055), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n800), .A2(new_n838), .B1(new_n831), .B2(new_n643), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n806), .A2(new_n1019), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n797), .A2(new_n832), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n1062));
  INV_X1    g0862(.A(new_n802), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n1061), .A2(new_n1062), .B1(G283), .B2(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n824), .B2(new_n817), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT49), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n781), .B1(G326), .B2(new_n813), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n223), .C2(new_n819), .ZN(new_n1068));
  INV_X1    g0868(.A(G159), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n800), .A2(new_n1069), .B1(new_n819), .B2(new_n228), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n818), .A2(G77), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n873), .B2(new_n812), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT114), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(new_n481), .B2(new_n797), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1070), .B(new_n1074), .C1(new_n1073), .C2(new_n1072), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n781), .C1(new_n203), .C2(new_n831), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1063), .A2(new_n599), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n207), .B2(new_n806), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT115), .Z(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT117), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n1045), .B(new_n1057), .C1(new_n1081), .C2(new_n792), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1082), .A2(new_n777), .B1(new_n776), .B2(new_n1013), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1013), .A2(new_n770), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1013), .A2(new_n770), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n724), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(KEYINPUT120), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1000), .A2(new_n717), .A3(new_n1004), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n717), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(new_n724), .A3(new_n1015), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n802), .A2(new_n251), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n807), .A2(G159), .B1(new_n799), .B2(G150), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1093), .B(new_n1095), .C1(G50), .C2(new_n796), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G68), .A2(new_n818), .B1(new_n820), .B2(G87), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n781), .B(new_n1097), .C1(new_n872), .C2(new_n812), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT118), .Z(new_n1099));
  OAI211_X1 g0899(.A(new_n1096), .B(new_n1099), .C1(new_n441), .C2(new_n831), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT119), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n800), .A2(new_n1019), .B1(new_n832), .B2(new_n806), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n797), .A2(new_n643), .B1(new_n819), .B2(new_n302), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n817), .A2(new_n827), .B1(new_n812), .B2(new_n838), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n431), .B1(new_n802), .B2(new_n223), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1103), .B(new_n1107), .C1(new_n824), .C2(new_n831), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n795), .B1(new_n1109), .B2(new_n792), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n793), .B1(new_n228), .B2(new_n219), .C1(new_n247), .C2(new_n1040), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n967), .A2(new_n791), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n776), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1088), .B1(new_n1092), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1092), .A2(new_n1115), .A3(new_n1088), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(G390));
  NOR2_X1   g0919(.A1(new_n851), .A2(new_n694), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n920), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n949), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n898), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT38), .B1(new_n898), .B2(new_n914), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT39), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n932), .A2(new_n918), .A3(new_n943), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n950), .C2(new_n942), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n942), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n703), .B1(new_n741), .B2(new_n684), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n846), .B1(new_n1129), .B2(new_n850), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1128), .B(new_n933), .C1(new_n1130), .C2(new_n949), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1122), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n854), .A2(new_n847), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n948), .B1(new_n768), .B2(new_n1120), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n1122), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n768), .A2(new_n948), .A3(new_n1120), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1121), .A2(new_n949), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1130), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n402), .A2(new_n464), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n546), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1141), .A2(G330), .A3(new_n1142), .A4(new_n920), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n939), .A2(new_n692), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1140), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1137), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1127), .A2(new_n1147), .A3(new_n1131), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1133), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1144), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1127), .A2(new_n1147), .A3(new_n1131), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1132), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n724), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n776), .B1(new_n1151), .B2(new_n1132), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1125), .A2(new_n789), .A3(new_n1126), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n481), .A2(new_n884), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n351), .B1(new_n797), .B2(new_n1035), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n799), .A2(G128), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n1069), .B2(new_n802), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G50), .C2(new_n820), .ZN(new_n1160));
  XOR2_X1   g0960(.A(KEYINPUT54), .B(G143), .Z(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n831), .A2(new_n1162), .B1(new_n812), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT53), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n817), .B2(new_n873), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n818), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1160), .B(new_n1168), .C1(new_n880), .C2(new_n806), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n831), .A2(new_n228), .B1(new_n806), .B2(new_n223), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n836), .B2(G87), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n800), .A2(new_n827), .B1(new_n797), .B2(new_n302), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1172), .A2(new_n351), .A3(new_n877), .A4(new_n1093), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n824), .C2(new_n812), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n795), .B1(new_n1175), .B2(new_n792), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1155), .A2(new_n1156), .A3(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1154), .A2(KEYINPUT121), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT121), .B1(new_n1154), .B2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1153), .B1(new_n1178), .B2(new_n1179), .ZN(G378));
  OAI21_X1  g0980(.A(new_n429), .B1(new_n460), .B2(new_n463), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n450), .A2(new_n452), .A3(new_n701), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT55), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT55), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n1183), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT56), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1186), .A2(KEYINPUT56), .A3(new_n1189), .ZN(new_n1193));
  AND2_X1   g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n789), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n884), .A2(new_n207), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G58), .A2(new_n820), .B1(new_n813), .B2(G283), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1071), .C1(new_n302), .C2(new_n806), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G68), .B2(new_n1063), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n781), .A2(new_n723), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n800), .A2(new_n223), .B1(new_n797), .B2(new_n228), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n599), .B2(new_n810), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT58), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G125), .A2(new_n799), .B1(new_n796), .B2(G132), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n807), .A2(G128), .B1(new_n810), .B2(G137), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1063), .A2(G150), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n818), .A2(new_n1161), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n813), .A2(G124), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n820), .C2(G159), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1204), .B(new_n1214), .C1(new_n1200), .C2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n795), .B1(new_n1216), .B2(new_n792), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1195), .A2(new_n1196), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n925), .A2(new_n933), .A3(KEYINPUT40), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n920), .A2(new_n924), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n918), .B2(new_n917), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G330), .B(new_n1221), .C1(new_n1223), .C2(KEYINPUT40), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1224), .A2(new_n946), .A3(new_n951), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n946), .B2(new_n951), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1220), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n952), .A2(new_n935), .A3(G330), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(new_n946), .A3(new_n951), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1194), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1219), .B1(new_n1231), .B2(new_n776), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1227), .A2(new_n1230), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n724), .B1(new_n1233), .B2(KEYINPUT57), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1152), .A2(new_n1145), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1228), .A2(new_n1194), .A3(new_n1229), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1194), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1235), .B(KEYINPUT57), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1232), .B1(new_n1234), .B2(new_n1239), .ZN(G375));
  OAI22_X1  g1040(.A1(new_n831), .A2(new_n302), .B1(new_n812), .B2(new_n643), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n836), .B2(G97), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n807), .A2(G283), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n351), .B1(new_n820), .B2(G77), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT122), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1077), .B1(new_n797), .B2(new_n223), .C1(new_n824), .C2(new_n800), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1243), .A3(new_n1245), .A4(new_n1247), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(G58), .A2(new_n820), .B1(new_n813), .B2(G128), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n1249), .B1(new_n880), .B2(new_n800), .C1(new_n797), .C2(new_n1162), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G159), .B2(new_n836), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n831), .A2(new_n873), .B1(new_n802), .B2(new_n207), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(KEYINPUT123), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n781), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n806), .A2(new_n1035), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1248), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n795), .B1(new_n1256), .B2(new_n792), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n948), .B2(new_n790), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n203), .B2(new_n884), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1140), .B2(new_n776), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1136), .A2(new_n1144), .A3(new_n1139), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n995), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1262), .B2(new_n1150), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(KEYINPUT124), .ZN(G381));
  INV_X1    g1064(.A(new_n1154), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1177), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1153), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G375), .A2(G396), .A3(G393), .A4(new_n1268), .ZN(new_n1269));
  NOR4_X1   g1069(.A1(G390), .A2(G387), .A3(G381), .A4(G384), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G407));
  OAI21_X1  g1071(.A(new_n776), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1218), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT57), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n730), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1273), .B1(new_n1276), .B2(new_n1238), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1268), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n702), .A3(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(G407), .A2(G213), .A3(new_n1279), .ZN(G409));
  NAND3_X1  g1080(.A1(G387), .A2(new_n1118), .A3(new_n1117), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1118), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1043), .B(new_n1017), .C1(new_n1282), .C2(new_n1116), .ZN(new_n1283));
  INV_X1    g1083(.A(G396), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G393), .B(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1231), .A2(new_n995), .A3(new_n1235), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1268), .B1(new_n1232), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1277), .B2(G378), .ZN(new_n1291));
  INV_X1    g1091(.A(G213), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(G343), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT60), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1261), .A2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1136), .A2(new_n1144), .A3(KEYINPUT60), .A4(new_n1139), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1146), .A3(new_n724), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1260), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT125), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G384), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n862), .A2(KEYINPUT125), .A3(new_n886), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1301), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n1260), .A3(new_n1297), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(new_n1291), .A2(KEYINPUT62), .A3(new_n1293), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT62), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G378), .B(new_n1232), .C1(new_n1234), .C2(new_n1239), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1289), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1278), .B1(new_n1310), .B2(new_n1273), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1293), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1308), .B1(new_n1312), .B2(new_n1305), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1307), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1293), .ZN(new_n1316));
  INV_X1    g1116(.A(G2897), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1305), .B(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1315), .B1(new_n1312), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1288), .B1(new_n1314), .B2(new_n1322), .ZN(new_n1323));
  AOI211_X1 g1123(.A(new_n1293), .B(new_n1306), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1305), .B(new_n1318), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1325), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1324), .B1(new_n1326), .B2(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1316), .A4(new_n1305), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1288), .ZN(new_n1330));
  NOR3_X1   g1130(.A1(new_n1327), .A2(KEYINPUT61), .A3(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(KEYINPUT126), .B1(new_n1323), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1312), .A2(new_n1305), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1312), .A2(new_n1320), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1333), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1336), .A2(new_n1315), .A3(new_n1288), .A4(new_n1329), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1307), .A2(new_n1321), .A3(new_n1313), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1337), .B(new_n1338), .C1(new_n1288), .C2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1332), .A2(new_n1340), .ZN(G405));
  NOR2_X1   g1141(.A1(new_n1277), .A2(new_n1268), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1309), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(KEYINPUT127), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT127), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1346), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1345), .A2(new_n1306), .A3(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1344), .A2(KEYINPUT127), .A3(new_n1305), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1288), .ZN(G402));
endmodule


