//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1281,
    new_n1282, new_n1283;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g0008(.A(KEYINPUT65), .B(G238), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n208), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n208), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g0023(.A(G50), .B1(G58), .B2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n206), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AND4_X1   g0028(.A1(new_n218), .A2(new_n222), .A3(new_n223), .A4(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  AND2_X1   g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  OAI211_X1 g0048(.A(G264), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT83), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT83), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(G264), .A4(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n247), .A2(new_n248), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G303), .ZN(new_n259));
  INV_X1    g0059(.A(G1698), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(G257), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n250), .A2(new_n257), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n226), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n205), .A2(G45), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT5), .A2(G41), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT5), .A2(G41), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT68), .B1(new_n263), .B2(new_n226), .ZN(new_n271));
  AND2_X1   g0071(.A1(G1), .A2(G13), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n270), .A2(G274), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G45), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G1), .ZN(new_n278));
  INV_X1    g0078(.A(new_n269), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n267), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n280), .A2(new_n271), .A3(G270), .A4(new_n275), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n265), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT21), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G116), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n205), .A2(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n285), .A2(new_n289), .A3(new_n226), .A4(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n288), .B1(new_n291), .B2(new_n287), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n290), .A2(new_n226), .B1(G20), .B2(new_n287), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  INV_X1    g0094(.A(G97), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n294), .B(new_n206), .C1(G33), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT20), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(KEYINPUT20), .A3(new_n296), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n283), .A2(new_n284), .A3(G169), .A4(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n276), .A2(new_n281), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n264), .B2(new_n262), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n293), .A2(KEYINPUT20), .A3(new_n296), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n297), .ZN(new_n306));
  OAI21_X1  g0106(.A(G169), .B1(new_n306), .B2(new_n292), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT21), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n304), .A2(G179), .A3(new_n301), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n265), .A2(G190), .A3(new_n282), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n311), .B(new_n300), .C1(new_n312), .C2(new_n304), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT84), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n309), .A2(KEYINPUT84), .A3(new_n310), .A4(new_n313), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n290), .A2(new_n226), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n206), .A2(G33), .ZN(new_n321));
  XNOR2_X1  g0121(.A(new_n321), .B(KEYINPUT69), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G50), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n210), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G20), .A2(G33), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(G20), .B1(G150), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n320), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT70), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n286), .A2(new_n319), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n326), .B1(new_n205), .B2(G20), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(new_n326), .B2(new_n286), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT9), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n271), .A2(new_n275), .A3(new_n341), .A4(G274), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n271), .A2(new_n275), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(G226), .A3(new_n340), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n258), .A2(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G222), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n260), .B1(new_n253), .B2(new_n254), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(G223), .B1(new_n258), .B2(G77), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n264), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n342), .B(new_n344), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G200), .B2(new_n351), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n339), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT10), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(KEYINPUT72), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n355), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT72), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n339), .A2(new_n354), .A3(new_n361), .A4(KEYINPUT10), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n351), .A2(G179), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n351), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n338), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n360), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n255), .A2(G232), .A3(G1698), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n255), .A2(G226), .A3(new_n260), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n264), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n271), .A2(new_n275), .A3(G238), .A4(new_n340), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n342), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT13), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n372), .B2(new_n375), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  INV_X1    g0181(.A(new_n370), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n345), .B2(G226), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n350), .B1(new_n383), .B2(new_n368), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT13), .B1(new_n384), .B2(new_n374), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n377), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n387), .A3(G169), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT73), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n377), .A2(G179), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n379), .A2(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n321), .B(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G77), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n206), .A2(new_n252), .ZN(new_n399));
  OR3_X1    g0199(.A1(new_n399), .A2(KEYINPUT74), .A3(new_n326), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n326), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT74), .B1(new_n210), .B2(G20), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n319), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT11), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT11), .B(new_n319), .C1(new_n398), .C2(new_n403), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT12), .B1(new_n285), .B2(G68), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n285), .A2(KEYINPUT12), .A3(G68), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n210), .B1(new_n205), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n408), .A2(new_n409), .B1(new_n335), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n394), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n412), .B1(new_n386), .B2(G200), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n390), .A2(G190), .A3(new_n392), .A4(new_n377), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n323), .B1(new_n205), .B2(G20), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n335), .B1(new_n286), .B2(new_n323), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT7), .B1(new_n258), .B2(new_n206), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n253), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n254), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n327), .A2(new_n210), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G58), .A2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n329), .A2(G159), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT16), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n320), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n424), .A2(KEYINPUT16), .A3(new_n430), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n420), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n271), .A2(new_n275), .A3(G232), .A4(new_n340), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G87), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT75), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(KEYINPUT75), .A2(G33), .A3(G87), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  MUX2_X1   g0241(.A(G223), .B(G226), .S(G1698), .Z(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n255), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n342), .B(new_n436), .C1(new_n443), .C2(new_n350), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n364), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(G179), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n435), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n253), .A2(new_n206), .A3(new_n254), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT7), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n210), .B1(new_n451), .B2(new_n422), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n432), .B1(new_n452), .B2(new_n429), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(new_n434), .A3(new_n319), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n419), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n448), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n343), .A2(G244), .A3(new_n340), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n460), .A2(new_n342), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n255), .A2(G232), .A3(new_n260), .ZN(new_n462));
  INV_X1    g0262(.A(G107), .ZN(new_n463));
  INV_X1    g0263(.A(new_n347), .ZN(new_n464));
  OAI221_X1 g0264(.A(new_n462), .B1(new_n463), .B2(new_n255), .C1(new_n464), .C2(new_n209), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n264), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G200), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n335), .B(G77), .C1(G1), .C2(new_n206), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n286), .A2(new_n397), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT15), .B(G87), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n321), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(G20), .B2(G77), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n323), .B(KEYINPUT71), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n475), .B2(new_n399), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n476), .B2(new_n319), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n468), .B(new_n477), .C1(new_n352), .C2(new_n467), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n467), .A2(new_n364), .ZN(new_n479));
  INV_X1    g0279(.A(new_n477), .ZN(new_n480));
  INV_X1    g0280(.A(G179), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n461), .A2(new_n466), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n442), .A2(new_n255), .ZN(new_n485));
  INV_X1    g0285(.A(new_n441), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n264), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n488), .A2(new_n352), .A3(new_n342), .A4(new_n436), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n444), .A2(new_n312), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g0291(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n435), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n454), .A3(new_n419), .ZN(new_n495));
  OR2_X1    g0295(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n459), .A2(new_n484), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n367), .A2(new_n417), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n294), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n502), .B1(new_n347), .B2(G250), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n260), .C1(new_n247), .C2(new_n248), .ZN(new_n504));
  XOR2_X1   g0304(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n260), .A2(KEYINPUT4), .A3(G244), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT80), .B1(new_n258), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n507), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT80), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n255), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n503), .A2(new_n506), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n264), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n280), .A2(new_n271), .A3(G257), .A4(new_n275), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n276), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(G179), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n512), .B2(new_n264), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n364), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT6), .ZN(new_n520));
  AND2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n202), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n463), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT77), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n399), .B2(new_n397), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n329), .A2(KEYINPUT77), .A3(G77), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n524), .A2(G20), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n463), .B1(new_n451), .B2(new_n422), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT78), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI211_X1 g0331(.A(KEYINPUT78), .B(new_n463), .C1(new_n451), .C2(new_n422), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n319), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n286), .A2(new_n295), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n291), .B2(new_n295), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n519), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n519), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  INV_X1    g0341(.A(new_n537), .ZN(new_n542));
  OR2_X1    g0342(.A1(new_n518), .A2(new_n312), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n518), .A2(G190), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n539), .A2(new_n541), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n206), .B1(new_n370), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G87), .B2(new_n203), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n206), .B(G68), .C1(new_n247), .C2(new_n248), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n321), .B2(new_n295), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n319), .ZN(new_n553));
  XOR2_X1   g0353(.A(KEYINPUT15), .B(G87), .Z(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n285), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT82), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT82), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  INV_X1    g0360(.A(new_n291), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n558), .A2(new_n560), .B1(G87), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G244), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n563));
  OAI211_X1 g0363(.A(G238), .B(new_n260), .C1(new_n247), .C2(new_n248), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n564), .C1(new_n252), .C2(new_n287), .ZN(new_n565));
  AOI21_X1  g0365(.A(G250), .B1(new_n205), .B2(G45), .ZN(new_n566));
  INV_X1    g0366(.A(G274), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n278), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n565), .A2(new_n264), .B1(new_n343), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(new_n312), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(G190), .B2(new_n569), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n559), .B1(new_n553), .B2(new_n556), .ZN(new_n572));
  AOI211_X1 g0372(.A(KEYINPUT82), .B(new_n555), .C1(new_n552), .C2(new_n319), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n572), .A2(new_n573), .B1(new_n291), .B2(new_n472), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n569), .A2(G169), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n565), .A2(new_n264), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n343), .A2(new_n568), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(new_n481), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n562), .A2(new_n571), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n280), .A2(new_n271), .A3(new_n275), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(G1698), .C1(new_n247), .C2(new_n248), .ZN(new_n582));
  OAI211_X1 g0382(.A(G250), .B(new_n260), .C1(new_n247), .C2(new_n248), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G294), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n581), .A2(G264), .B1(new_n585), .B2(new_n264), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n586), .A2(new_n276), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n481), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n276), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n364), .ZN(new_n590));
  XOR2_X1   g0390(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n463), .A3(G20), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n594), .C1(new_n287), .C2(new_n321), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT87), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n255), .A2(new_n206), .A3(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n598), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n255), .A2(new_n206), .A3(G87), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n591), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT87), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n595), .B(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n591), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(new_n599), .A4(new_n601), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n320), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n463), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT25), .B1(new_n286), .B2(new_n463), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n610), .A2(new_n611), .B1(new_n463), .B2(new_n291), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n588), .B(new_n590), .C1(new_n608), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n603), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n319), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n586), .A2(new_n352), .A3(new_n276), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n587), .B2(G200), .ZN(new_n617));
  INV_X1    g0417(.A(new_n612), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n580), .A2(new_n613), .A3(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n318), .A2(new_n501), .A3(new_n546), .A4(new_n620), .ZN(G372));
  NAND2_X1  g0421(.A1(new_n360), .A2(new_n362), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n414), .A2(new_n415), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n413), .B1(new_n623), .B2(new_n483), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n499), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n622), .B1(new_n625), .B2(new_n459), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT91), .ZN(new_n627));
  INV_X1    g0427(.A(new_n366), .ZN(new_n628));
  OR3_X1    g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n501), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n539), .A2(new_n541), .A3(new_n580), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n574), .A2(new_n579), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n561), .A2(G87), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n572), .B2(new_n573), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT88), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(KEYINPUT88), .B(new_n636), .C1(new_n572), .C2(new_n573), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n635), .B1(new_n641), .B2(new_n571), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n518), .A2(new_n364), .ZN(new_n644));
  AOI211_X1 g0444(.A(new_n481), .B(new_n515), .C1(new_n264), .C2(new_n512), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n517), .B(KEYINPUT90), .C1(new_n364), .C2(new_n518), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(new_n537), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n642), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n635), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n634), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n613), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n309), .A2(new_n310), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n539), .A2(new_n541), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n612), .B1(new_n614), .B2(new_n319), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n545), .A2(new_n542), .B1(new_n657), .B2(new_n617), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n658), .A3(new_n642), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n655), .B1(new_n659), .B2(KEYINPUT89), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT89), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n656), .A2(new_n658), .A3(new_n642), .A4(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n652), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n631), .B1(new_n632), .B2(new_n663), .ZN(G369));
  NAND3_X1  g0464(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n301), .A2(new_n670), .ZN(new_n671));
  MUX2_X1   g0471(.A(new_n654), .B(new_n318), .S(new_n671), .Z(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n653), .A2(new_n670), .ZN(new_n675));
  INV_X1    g0475(.A(new_n670), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n613), .B(new_n619), .C1(new_n657), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT92), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n654), .A2(new_n676), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n613), .B2(new_n670), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT93), .Z(new_n685));
  NAND2_X1  g0485(.A1(new_n681), .A2(new_n685), .ZN(G399));
  INV_X1    g0486(.A(new_n219), .ZN(new_n687));
  OR3_X1    g0487(.A1(new_n687), .A2(KEYINPUT94), .A3(G41), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT94), .B1(new_n687), .B2(G41), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n691), .A2(new_n205), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n225), .B2(new_n691), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT28), .Z(new_n696));
  NAND2_X1  g0496(.A1(new_n642), .A2(new_n648), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(KEYINPUT26), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n539), .A2(new_n649), .A3(new_n580), .A4(new_n541), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(KEYINPUT98), .A3(new_n651), .A4(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT98), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n651), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n649), .B1(new_n642), .B2(new_n648), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n659), .A2(new_n655), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n700), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n663), .A2(new_n670), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(KEYINPUT29), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT97), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT31), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n265), .A2(new_n586), .A3(new_n569), .A4(new_n282), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n645), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(KEYINPUT30), .B1(new_n517), .B2(new_n712), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n304), .A2(G179), .A3(new_n569), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n587), .A2(new_n518), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n670), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n715), .A2(new_n716), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n717), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n722), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(new_n710), .B(new_n711), .C1(new_n721), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n723), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n676), .A2(new_n711), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT95), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT95), .ZN(new_n729));
  INV_X1    g0529(.A(new_n727), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n719), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n318), .A2(new_n546), .A3(new_n620), .A4(new_n676), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n725), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n719), .A2(new_n720), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n670), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n710), .B1(new_n737), .B2(new_n711), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n709), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n696), .B1(new_n741), .B2(G1), .ZN(G364));
  AND2_X1   g0542(.A1(new_n206), .A2(G13), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n205), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n674), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G330), .B2(new_n672), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n219), .A2(new_n255), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT99), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G355), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G116), .B2(new_n219), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n242), .A2(new_n277), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n687), .A2(new_n255), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n277), .B2(new_n225), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT100), .ZN(new_n758));
  OAI21_X1  g0558(.A(G20), .B1(new_n758), .B2(G169), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n364), .A2(KEYINPUT100), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n272), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT101), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT101), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n746), .B1(new_n757), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n206), .A2(new_n481), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(KEYINPUT102), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(G317), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G311), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(G179), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n781), .ZN(new_n785));
  INV_X1    g0585(.A(G329), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n771), .A2(G190), .A3(new_n312), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n255), .B(new_n787), .C1(G322), .C2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n772), .A2(new_n352), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G326), .B1(new_n793), .B2(G303), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n352), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n206), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n784), .A2(new_n352), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n797), .A2(G294), .B1(new_n799), .B2(G283), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n780), .A2(new_n790), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT104), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n295), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n255), .B1(new_n782), .B2(new_n397), .C1(new_n327), .C2(new_n788), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(G87), .C2(new_n793), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n777), .A2(G68), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n791), .A2(G50), .B1(new_n799), .B2(G107), .ZN(new_n808));
  INV_X1    g0608(.A(new_n785), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G159), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT32), .Z(new_n811));
  NAND4_X1  g0611(.A1(new_n806), .A2(new_n807), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n801), .A2(new_n802), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n803), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n770), .B1(new_n814), .B2(new_n764), .ZN(new_n815));
  INV_X1    g0615(.A(new_n767), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n672), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT105), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n748), .A2(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n480), .A2(new_n670), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n484), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT108), .B1(new_n483), .B2(new_n676), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n477), .B1(new_n467), .B2(new_n364), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT108), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n823), .A2(new_n824), .A3(new_n482), .A4(new_n670), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n676), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n708), .A2(new_n827), .B1(new_n663), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n746), .B1(new_n829), .B2(new_n740), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n740), .B2(new_n829), .ZN(new_n831));
  INV_X1    g0631(.A(new_n746), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n764), .A2(new_n765), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n397), .ZN(new_n834));
  INV_X1    g0634(.A(new_n764), .ZN(new_n835));
  INV_X1    g0635(.A(new_n782), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n789), .A2(G143), .B1(new_n836), .B2(G159), .ZN(new_n837));
  INV_X1    g0637(.A(G137), .ZN(new_n838));
  INV_X1    g0638(.A(new_n791), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n777), .B2(G150), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n255), .B1(new_n785), .B2(new_n844), .C1(new_n326), .C2(new_n792), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n796), .A2(new_n327), .B1(new_n798), .B2(new_n210), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n842), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G303), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n839), .A2(new_n848), .B1(new_n782), .B2(new_n287), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n777), .B2(G283), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT106), .ZN(new_n851));
  INV_X1    g0651(.A(G294), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n258), .B1(new_n785), .B2(new_n783), .C1(new_n788), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n792), .A2(new_n463), .ZN(new_n854));
  INV_X1    g0654(.A(G87), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n798), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g0656(.A1(new_n853), .A2(new_n804), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n847), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n835), .B1(new_n858), .B2(KEYINPUT107), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n834), .B1(new_n766), .B2(new_n827), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n831), .A2(new_n862), .ZN(G384));
  OR2_X1    g0663(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(G116), .A3(new_n227), .A4(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OAI211_X1 g0667(.A(new_n225), .B(G77), .C1(new_n327), .C2(new_n210), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n326), .A2(G68), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n205), .B(G13), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n484), .A2(new_n820), .B1(new_n822), .B2(new_n825), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n412), .A2(new_n670), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n413), .A2(new_n416), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n412), .B(new_n670), .C1(new_n623), .C2(new_n394), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n668), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n455), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n498), .B2(new_n458), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n448), .A2(new_n455), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n879), .A3(new_n495), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n882), .A2(new_n879), .A3(new_n885), .A4(new_n495), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT38), .B1(new_n881), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n877), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n711), .B1(new_n721), .B2(new_n724), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n736), .A4(new_n670), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n733), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n872), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n881), .A2(new_n887), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n881), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n733), .A2(new_n891), .A3(new_n892), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .A4(new_n877), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT110), .ZN(new_n903));
  OR3_X1    g0703(.A1(new_n903), .A2(new_n632), .A3(new_n893), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n903), .B1(new_n632), .B2(new_n893), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(G330), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n875), .A2(new_n876), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n542), .A2(new_n544), .A3(new_n543), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n519), .A2(new_n540), .A3(new_n537), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n540), .B1(new_n519), .B2(new_n537), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n909), .B(new_n619), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n558), .A2(new_n560), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT88), .B1(new_n913), .B2(new_n636), .ZN(new_n914));
  INV_X1    g0714(.A(new_n640), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n571), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n651), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT89), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n655), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n662), .A3(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n634), .A2(new_n650), .A3(new_n651), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n828), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n483), .A2(new_n670), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT109), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT109), .ZN(new_n925));
  INV_X1    g0725(.A(new_n923), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n925), .B(new_n926), .C1(new_n663), .C2(new_n828), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n908), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n899), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n458), .A2(new_n668), .ZN(new_n930));
  INV_X1    g0730(.A(new_n899), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT39), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n899), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n413), .A2(new_n670), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n930), .A3(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n707), .B(new_n501), .C1(new_n708), .C2(KEYINPUT29), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n631), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n937), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n906), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n205), .B2(new_n743), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n906), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n871), .B1(new_n942), .B2(new_n943), .ZN(G367));
  OAI21_X1  g0744(.A(new_n546), .B1(new_n542), .B2(new_n676), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n648), .A2(new_n670), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n948), .A2(new_n683), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT42), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n656), .B1(new_n948), .B2(new_n613), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n676), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n639), .A2(new_n640), .A3(new_n670), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n642), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n651), .B2(new_n953), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n950), .A2(new_n952), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n956), .B(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n680), .A2(new_n947), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n690), .B(KEYINPUT41), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n685), .A2(new_n947), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT45), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n685), .A2(new_n947), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n680), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n675), .A2(new_n677), .A3(new_n682), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n683), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT111), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n673), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n673), .B(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n971), .B1(new_n972), .B2(new_n969), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n963), .A2(new_n681), .A3(new_n965), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n967), .A2(new_n741), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n961), .B1(new_n975), .B2(new_n741), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n960), .B1(new_n976), .B2(new_n745), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT112), .B1(new_n792), .B2(new_n287), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT46), .Z(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n852), .B2(new_n776), .ZN(new_n980));
  AOI22_X1  g0780(.A1(G107), .A2(new_n797), .B1(new_n791), .B2(G311), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n255), .B1(new_n836), .B2(G283), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n789), .A2(G303), .B1(new_n809), .B2(G317), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n799), .A2(G97), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n797), .A2(G68), .B1(new_n793), .B2(G58), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n791), .A2(G143), .B1(new_n799), .B2(G77), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n258), .B1(new_n789), .B2(G150), .ZN(new_n988));
  AOI22_X1  g0788(.A1(G50), .A2(new_n836), .B1(new_n809), .B2(G137), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G159), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n776), .A2(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n980), .A2(new_n985), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n835), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n754), .A2(new_n237), .B1(new_n687), .B2(new_n554), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n832), .B1(new_n997), .B2(new_n768), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(new_n955), .C2(new_n816), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n977), .A2(new_n999), .ZN(G387));
  NAND3_X1  g0800(.A1(new_n675), .A2(new_n677), .A3(new_n767), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n750), .A2(new_n693), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n219), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n755), .B1(new_n234), .B2(G45), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n475), .A2(G50), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1006));
  OR2_X1    g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n693), .C1(G68), .C2(G77), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1003), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n746), .B1(new_n1011), .B2(new_n769), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n789), .A2(G317), .B1(new_n836), .B2(G303), .ZN(new_n1013));
  INV_X1    g0813(.A(G322), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1013), .B1(new_n1014), .B2(new_n839), .C1(new_n776), .C2(new_n783), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT48), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  INV_X1    g0818(.A(G283), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n796), .A2(new_n1019), .B1(new_n792), .B2(new_n852), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT115), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT49), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n798), .A2(new_n287), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n255), .B(new_n1026), .C1(G326), .C2(new_n809), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n776), .A2(new_n323), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n788), .A2(new_n326), .B1(new_n782), .B2(new_n210), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n258), .B(new_n1030), .C1(G150), .C2(new_n809), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n792), .A2(new_n397), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G97), .B2(new_n799), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n554), .A2(new_n797), .B1(new_n791), .B2(G159), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1028), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1012), .B1(new_n1036), .B2(new_n764), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n973), .A2(new_n745), .B1(new_n1001), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n741), .A2(new_n973), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n691), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n741), .A2(new_n973), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(new_n974), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n681), .B1(new_n963), .B2(new_n965), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1043), .A2(new_n744), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n948), .A2(new_n767), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n755), .A2(new_n245), .B1(new_n295), .B2(new_n219), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n746), .B1(new_n1047), .B2(new_n769), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n258), .B(new_n856), .C1(G143), .C2(new_n809), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n796), .A2(new_n397), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G68), .B2(new_n793), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n326), .B2(new_n776), .C1(new_n475), .C2(new_n782), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G150), .A2(new_n791), .B1(new_n789), .B2(G159), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n258), .B1(new_n785), .B2(new_n1014), .C1(new_n852), .C2(new_n782), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n796), .A2(new_n287), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n463), .A2(new_n798), .B1(new_n792), .B2(new_n1019), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n776), .B2(new_n848), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G317), .A2(new_n791), .B1(new_n789), .B2(G311), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT52), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n1053), .A2(new_n1055), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1048), .B1(new_n1063), .B2(new_n764), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1045), .B1(new_n1046), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n975), .A3(new_n691), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(G390));
  NAND3_X1  g0868(.A1(new_n900), .A2(G330), .A3(new_n827), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n908), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n706), .A2(new_n676), .A3(new_n827), .ZN(new_n1071));
  AND3_X1   g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n926), .ZN(new_n1072));
  OAI211_X1 g0872(.A(G330), .B(new_n827), .C1(new_n734), .C2(new_n738), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(new_n908), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n908), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n900), .A2(G330), .A3(new_n827), .A4(new_n907), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n924), .A2(new_n927), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n501), .A2(G330), .A3(new_n900), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n631), .A2(new_n938), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT116), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n932), .A2(new_n934), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n928), .B2(new_n935), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n931), .A2(new_n935), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n1071), .A2(new_n926), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n1089), .B2(new_n908), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1087), .A2(new_n1090), .A3(new_n1074), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1077), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1085), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1077), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT116), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1072), .A2(new_n1074), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1097), .B1(new_n1098), .B2(new_n1083), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1087), .A2(new_n1090), .A3(new_n1074), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1096), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1093), .A2(new_n1101), .A3(new_n691), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n255), .B1(new_n788), .B2(new_n844), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n791), .A2(G128), .B1(new_n799), .B2(G50), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n991), .B2(new_n796), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G125), .C2(new_n809), .ZN(new_n1106));
  INV_X1    g0906(.A(G150), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n792), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT117), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n777), .A2(G137), .B1(new_n836), .B2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1106), .B(new_n1110), .C1(new_n1111), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1114), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n776), .A2(new_n463), .B1(new_n295), .B2(new_n782), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT119), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n258), .B1(new_n788), .B2(new_n287), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G294), .B2(new_n809), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n210), .A2(new_n798), .B1(new_n792), .B2(new_n855), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1050), .B(new_n1124), .C1(G283), .C2(new_n791), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1115), .A2(new_n1117), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n764), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n833), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n746), .C1(new_n324), .C2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1086), .B2(new_n765), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n745), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1102), .A2(new_n1133), .ZN(G378));
  NAND3_X1  g0934(.A1(new_n1096), .A2(new_n1100), .A3(new_n1081), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1084), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n338), .A2(new_n878), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT122), .Z(new_n1139));
  NAND2_X1  g0939(.A1(new_n367), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n360), .A3(new_n362), .A4(new_n366), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1143), .B(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n894), .A2(G330), .A3(new_n901), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n1147), .A3(KEYINPUT123), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT123), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n894), .A2(new_n1150), .A3(new_n901), .A4(G330), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1143), .B(new_n1144), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1149), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n936), .A2(new_n930), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(new_n928), .B2(new_n899), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1147), .A2(KEYINPUT123), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n937), .A2(new_n1159), .A3(new_n1148), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1137), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n690), .B1(new_n1136), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1135), .A2(new_n1084), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(KEYINPUT57), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1152), .A2(new_n765), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n839), .A2(new_n287), .B1(new_n798), .B2(new_n327), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1032), .B(new_n1167), .C1(G68), .C2(new_n797), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n255), .A2(G41), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n788), .A2(new_n463), .B1(new_n782), .B2(new_n472), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(G283), .C2(new_n809), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1168), .B(new_n1171), .C1(new_n295), .C2(new_n776), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT58), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1169), .B(new_n326), .C1(G33), .C2(G41), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n789), .A2(G128), .B1(new_n836), .B2(G137), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n792), .B2(new_n1112), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G150), .A2(new_n797), .B1(new_n791), .B2(G125), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT120), .Z(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G132), .C2(new_n777), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT121), .Z(new_n1183));
  OR2_X1    g0983(.A1(new_n1183), .A2(KEYINPUT59), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n991), .B2(new_n798), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n1183), .B2(KEYINPUT59), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1174), .B(new_n1177), .C1(new_n1184), .C2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1188), .A2(new_n835), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n832), .B(new_n1189), .C1(new_n326), .C2(new_n833), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1165), .A2(new_n745), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1164), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1098), .A2(new_n1083), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n961), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n908), .A2(new_n765), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n746), .B1(new_n1129), .B2(G68), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n777), .A2(new_n1113), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n788), .A2(new_n838), .B1(new_n782), .B2(new_n1107), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n258), .B(new_n1200), .C1(G128), .C2(new_n809), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n791), .A2(G132), .B1(new_n799), .B2(G58), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n797), .A2(G50), .B1(new_n793), .B2(G159), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n839), .A2(new_n852), .B1(new_n782), .B2(new_n463), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n777), .B2(G116), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT124), .Z(new_n1207));
  OAI21_X1  g1007(.A(new_n258), .B1(new_n788), .B2(new_n1019), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G303), .B2(new_n809), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n797), .A2(new_n554), .B1(new_n799), .B2(G77), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(new_n295), .C2(new_n792), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1207), .B2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1198), .B1(new_n1212), .B2(new_n764), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1081), .A2(new_n745), .B1(new_n1197), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1196), .A2(new_n1214), .ZN(G381));
  OR4_X1    g1015(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1102), .A2(new_n1133), .A3(new_n1218), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1191), .A3(new_n1164), .ZN(new_n1221));
  OR4_X1    g1021(.A1(G387), .A2(new_n1216), .A3(G381), .A4(new_n1221), .ZN(G407));
  OAI211_X1 g1022(.A(G407), .B(G213), .C1(G343), .C2(new_n1221), .ZN(G409));
  INV_X1    g1023(.A(G390), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G387), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n977), .A2(G390), .A3(new_n999), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g1027(.A(G393), .B(G396), .Z(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(new_n1228), .A3(new_n1226), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT61), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n669), .A2(G213), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(G2897), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1098), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n691), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1193), .A2(KEYINPUT60), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1238), .B1(new_n1194), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1214), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n862), .B(new_n831), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1239), .A2(new_n1194), .ZN(new_n1243));
  OAI211_X1 g1043(.A(G384), .B(new_n1214), .C1(new_n1243), .C2(new_n1238), .ZN(new_n1244));
  AOI211_X1 g1044(.A(KEYINPUT127), .B(new_n1236), .C1(new_n1242), .C2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT127), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G2897), .B(new_n1235), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1245), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1136), .A2(new_n1195), .A3(new_n1165), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1191), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1217), .A2(new_n1252), .A3(new_n1219), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1091), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1161), .B1(new_n1254), .B2(new_n1083), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n691), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT57), .B1(new_n1136), .B2(new_n1165), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G378), .B(new_n1191), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT126), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT126), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1164), .A2(new_n1260), .A3(G378), .A4(new_n1191), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1253), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1250), .B1(new_n1262), .B2(new_n1235), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1262), .A2(new_n1235), .A3(new_n1246), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1233), .B(new_n1263), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1253), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1246), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1234), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1232), .B1(new_n1266), .B2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1263), .A2(new_n1233), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1271), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1264), .A2(KEYINPUT63), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1279), .ZN(G405));
  NAND2_X1  g1080(.A1(new_n1220), .A2(G375), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1267), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1270), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1232), .ZN(G402));
endmodule


