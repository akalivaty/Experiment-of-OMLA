//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n547, new_n549, new_n550, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n592, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127, new_n1128;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n452), .A2(new_n457), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n464), .A3(G137), .ZN(new_n465));
  NAND2_X1  g040(.A1(G101), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G125), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n474), .B2(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n480), .A3(new_n473), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(KEYINPUT69), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n492), .A2(new_n462), .A3(new_n464), .A4(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n462), .A2(new_n464), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(new_n492), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT4), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n471), .B2(G126), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n495), .A2(G2105), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n505), .A2(new_n509), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n517), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XNOR2_X1  g097(.A(new_n506), .B(KEYINPUT6), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n510), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n511), .A2(new_n513), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n525), .A2(new_n528), .A3(new_n529), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  AOI22_X1  g108(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n519), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n527), .A2(G90), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n524), .A2(G52), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  AND2_X1   g114(.A1(new_n527), .A2(G81), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n519), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT71), .B(G43), .Z(new_n543));
  NOR2_X1   g118(.A1(new_n509), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g119(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND3_X1  g126(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G65), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n526), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n527), .A2(G91), .B1(new_n556), .B2(G651), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G299));
  NAND2_X1  g133(.A1(new_n524), .A2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n527), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  AOI22_X1  g137(.A1(G48), .A2(new_n524), .B1(new_n527), .B2(G86), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G61), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n526), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G651), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(KEYINPUT72), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT72), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n566), .B2(G651), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n563), .B1(new_n568), .B2(new_n570), .ZN(G305));
  NAND2_X1  g146(.A1(new_n527), .A2(G85), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n524), .A2(G47), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n519), .C2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G290));
  NAND2_X1  g153(.A1(G301), .A2(G868), .ZN(new_n579));
  INV_X1    g154(.A(G92), .ZN(new_n580));
  OR3_X1    g155(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G79), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n526), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n524), .A2(G54), .B1(new_n584), .B2(G651), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT10), .B1(new_n515), .B2(new_n580), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n579), .B1(new_n588), .B2(G868), .ZN(G284));
  XOR2_X1   g164(.A(G284), .B(KEYINPUT74), .Z(G321));
  NAND2_X1  g165(.A1(G286), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(G299), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G297));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(G868), .ZN(G280));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n588), .B1(new_n595), .B2(G860), .ZN(G148));
  NOR2_X1   g171(.A1(new_n545), .A2(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n587), .A2(G559), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n597), .B1(new_n599), .B2(G868), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT75), .ZN(G323));
  XNOR2_X1  g176(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g177(.A1(new_n482), .A2(G123), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n485), .A2(G135), .ZN(new_n604));
  OAI21_X1  g179(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n473), .A2(G111), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n603), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT77), .B(G2096), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT76), .B(G2100), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT78), .B(G2438), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(G2427), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT80), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n618), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n624), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G14), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(G401));
  XNOR2_X1  g208(.A(G2067), .B(G2678), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT81), .Z(new_n635));
  XOR2_X1   g210(.A(G2072), .B(G2078), .Z(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(KEYINPUT17), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n637), .B(new_n639), .C1(new_n635), .C2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n636), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n642), .A2(new_n634), .A3(new_n638), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT18), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n635), .A2(new_n640), .A3(new_n638), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XOR2_X1   g223(.A(G1971), .B(G1976), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(KEYINPUT20), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n655), .A2(new_n656), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n651), .A2(new_n654), .A3(new_n657), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n656), .C2(new_n655), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT83), .B(G1981), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G229));
  NOR2_X1   g243(.A1(G16), .A2(G24), .ZN(new_n669));
  XNOR2_X1  g244(.A(G290), .B(KEYINPUT84), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n669), .B1(new_n670), .B2(G16), .ZN(new_n671));
  INV_X1    g246(.A(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G22), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G166), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1971), .ZN(new_n677));
  NOR2_X1   g252(.A1(G16), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(G16), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT33), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(G6), .B(G305), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n673), .B(KEYINPUT85), .C1(KEYINPUT34), .C2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n482), .A2(G119), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n485), .A2(G131), .ZN(new_n691));
  OAI21_X1  g266(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n473), .A2(G107), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR3_X1   g272(.A1(new_n688), .A2(new_n689), .A3(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT36), .Z(new_n699));
  NAND2_X1  g274(.A1(KEYINPUT24), .A2(G34), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(KEYINPUT24), .A2(G34), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n701), .A2(new_n702), .A3(G29), .ZN(new_n703));
  INV_X1    g278(.A(G160), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G29), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G2084), .ZN(new_n707));
  NAND2_X1  g282(.A1(G171), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G5), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  NOR2_X1   g285(.A1(G4), .A2(G16), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n588), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT86), .B(G1348), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI221_X1 g290(.A(new_n707), .B1(new_n709), .B2(new_n710), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n710), .B2(new_n709), .ZN(new_n717));
  NOR2_X1   g292(.A1(G27), .A2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G164), .B2(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(G2078), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n482), .A2(G129), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n485), .A2(G141), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND4_X1  g300(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n727), .A2(new_n728), .A3(G29), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(G29), .B2(G32), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n731), .B2(new_n607), .ZN(new_n736));
  OR2_X1    g311(.A1(G29), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  AOI22_X1  g314(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  INV_X1    g315(.A(G139), .ZN(new_n741));
  OAI221_X1 g316(.A(new_n739), .B1(new_n473), .B2(new_n740), .C1(new_n484), .C2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n737), .B1(new_n742), .B2(new_n731), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT90), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G2084), .B2(new_n706), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n720), .A2(new_n736), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n731), .A2(G26), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT88), .Z(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G140), .B2(new_n485), .ZN(new_n754));
  INV_X1    g329(.A(G128), .ZN(new_n755));
  OAI21_X1  g330(.A(KEYINPUT87), .B1(new_n481), .B2(new_n755), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n755), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n749), .B(new_n750), .C1(new_n758), .C2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n749), .B2(new_n750), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT89), .B(G2067), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n731), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n731), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT29), .B(G2090), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n767), .A2(G28), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(G28), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n768), .A2(new_n769), .A3(G29), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n719), .A2(G2078), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n770), .B(new_n771), .C1(new_n744), .C2(new_n743), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n674), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n674), .ZN(new_n774));
  INV_X1    g349(.A(G1966), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT31), .B(G11), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n674), .A2(G19), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n545), .B2(new_n674), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n713), .A2(new_n715), .B1(G1341), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n780), .ZN(new_n781));
  NOR3_X1   g356(.A1(new_n762), .A2(new_n766), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n779), .A2(G1341), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n674), .A2(KEYINPUT23), .A3(G20), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G20), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n592), .C2(new_n674), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT92), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1956), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n748), .A2(new_n782), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT93), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n699), .A2(new_n792), .ZN(G150));
  INV_X1    g368(.A(G150), .ZN(G311));
  AOI22_X1  g369(.A1(G55), .A2(new_n524), .B1(new_n527), .B2(G93), .ZN(new_n795));
  NAND2_X1  g370(.A1(G80), .A2(G543), .ZN(new_n796));
  INV_X1    g371(.A(G67), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n526), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT94), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n795), .B1(new_n799), .B2(new_n519), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT95), .ZN(new_n801));
  INV_X1    g376(.A(G860), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT37), .ZN(new_n804));
  INV_X1    g379(.A(new_n545), .ZN(new_n805));
  MUX2_X1   g380(.A(new_n800), .B(new_n801), .S(new_n805), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n588), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT38), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT39), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT96), .Z(new_n811));
  OAI21_X1  g386(.A(new_n802), .B1(new_n809), .B2(KEYINPUT39), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(G145));
  XNOR2_X1  g388(.A(new_n742), .B(new_n611), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n503), .B(KEYINPUT97), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n694), .B(new_n726), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n485), .A2(G142), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n473), .A2(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G130), .B2(new_n482), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(new_n758), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n607), .B(new_n489), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n704), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(G37), .B1(new_n825), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n826), .B1(new_n825), .B2(new_n829), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g409(.A(new_n806), .B(new_n599), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n588), .B(G299), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT41), .Z(new_n837));
  AND2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT42), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(G290), .B(G288), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(G305), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n847), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n843), .A2(new_n844), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT100), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n841), .B1(new_n838), .B2(new_n840), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n842), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n851), .B1(new_n842), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(G868), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(G868), .B2(new_n801), .ZN(G295));
  OAI21_X1  g431(.A(new_n855), .B1(G868), .B2(new_n801), .ZN(G331));
  XNOR2_X1  g432(.A(G168), .B(G301), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n806), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n806), .A2(new_n858), .ZN(new_n860));
  OR3_X1    g435(.A1(new_n859), .A2(new_n860), .A3(new_n839), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n837), .B1(new_n859), .B2(new_n860), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n848), .A2(new_n850), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n861), .A2(new_n862), .A3(new_n850), .A4(new_n848), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT43), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n865), .A2(new_n870), .A3(new_n867), .A4(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n871), .A2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT44), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n869), .A2(KEYINPUT102), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n868), .A2(new_n880), .A3(KEYINPUT43), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n874), .B1(new_n878), .B2(new_n882), .ZN(G397));
  INV_X1    g458(.A(G8), .ZN(new_n884));
  INV_X1    g459(.A(G1384), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n496), .A2(new_n497), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n462), .A2(new_n464), .A3(G126), .ZN(new_n887));
  INV_X1    g462(.A(new_n501), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n886), .A2(new_n473), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n890));
  OAI211_X1 g465(.A(KEYINPUT45), .B(new_n885), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT109), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n503), .A2(new_n896), .A3(KEYINPUT45), .A4(new_n885), .ZN(new_n897));
  INV_X1    g472(.A(G40), .ZN(new_n898));
  AOI211_X1 g473(.A(new_n898), .B(new_n467), .C1(new_n474), .C2(new_n477), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n892), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n775), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(KEYINPUT50), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n887), .A2(new_n888), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n492), .B1(new_n471), .B2(G138), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(G2105), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n493), .A2(new_n494), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n473), .ZN(new_n907));
  AOI21_X1  g482(.A(G1384), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT50), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT110), .B(G2084), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(new_n910), .A3(new_n899), .A4(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n884), .B1(new_n901), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G286), .A2(G8), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT118), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT51), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT118), .ZN(new_n917));
  NAND3_X1  g492(.A1(G286), .A2(new_n917), .A3(G8), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT120), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT120), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n902), .A2(new_n910), .A3(new_n899), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n923), .A2(new_n911), .B1(new_n900), .B2(new_n775), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n921), .B(new_n922), .C1(new_n924), .C2(new_n884), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n915), .A2(new_n918), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n926), .A2(KEYINPUT119), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(KEYINPUT119), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n913), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n920), .B(new_n925), .C1(new_n929), .C2(new_n916), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n901), .A2(new_n912), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n926), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT121), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n895), .A2(new_n899), .A3(new_n891), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(G2078), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT122), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n902), .A2(new_n910), .A3(new_n899), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n710), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n938), .A2(new_n939), .ZN(new_n944));
  INV_X1    g519(.A(new_n891), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n945), .A2(new_n898), .A3(new_n467), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n476), .A2(G2105), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n936), .A2(G2078), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n946), .A2(new_n947), .A3(new_n895), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(G301), .B(KEYINPUT54), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n900), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n948), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n943), .A2(new_n944), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n953), .B1(new_n956), .B2(new_n952), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT104), .B(G2090), .Z(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n902), .A2(new_n910), .A3(new_n899), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1971), .ZN(new_n963));
  OAI211_X1 g538(.A(G40), .B(G160), .C1(new_n908), .C2(KEYINPUT45), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n945), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n937), .A2(KEYINPUT103), .A3(new_n963), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n972));
  OAI21_X1  g547(.A(G8), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n958), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n937), .A2(KEYINPUT103), .A3(new_n963), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT103), .B1(new_n937), .B2(new_n963), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n961), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n971), .A2(new_n972), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(KEYINPUT105), .A3(G8), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT123), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n679), .A2(G1976), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n899), .A2(new_n908), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT106), .B1(new_n985), .B2(G8), .ZN(new_n986));
  INV_X1    g561(.A(new_n467), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT67), .B1(new_n476), .B2(G2105), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n468), .B(new_n473), .C1(new_n475), .C2(new_n469), .ZN(new_n989));
  OAI211_X1 g564(.A(G40), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(KEYINPUT106), .B(G8), .C1(new_n990), .C2(new_n893), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n982), .B(new_n984), .C1(new_n986), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n563), .B(new_n994), .C1(new_n568), .C2(new_n570), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT107), .B(G86), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n567), .B1(new_n515), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n524), .A2(G48), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n995), .B2(new_n999), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n986), .A2(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n990), .A2(new_n893), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n884), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1006), .A2(new_n991), .B1(G1976), .B2(new_n679), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n993), .B(new_n1003), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n884), .B1(new_n965), .B2(new_n961), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(new_n978), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n980), .A2(new_n981), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n981), .B1(new_n980), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n957), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT124), .B1(new_n935), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT61), .ZN(new_n1017));
  INV_X1    g592(.A(new_n937), .ZN(new_n1018));
  XNOR2_X1  g593(.A(KEYINPUT56), .B(G2072), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT111), .B(G1956), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n941), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT112), .Z(new_n1025));
  NAND2_X1  g600(.A1(new_n553), .A2(KEYINPUT113), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT114), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G299), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(KEYINPUT114), .A3(new_n592), .ZN(new_n1031));
  OR2_X1    g606(.A1(KEYINPUT114), .A2(KEYINPUT57), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT115), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1030), .A2(new_n1035), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1022), .A2(new_n1025), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1022), .A2(new_n1025), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1017), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g615(.A1(new_n923), .A2(new_n714), .B1(G2067), .B2(new_n985), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(new_n588), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(KEYINPUT60), .ZN(new_n1043));
  INV_X1    g618(.A(G1996), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1018), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT58), .B(G1341), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n985), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n805), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1041), .A2(KEYINPUT60), .A3(new_n587), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1043), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT61), .A3(new_n1037), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1040), .A2(new_n1052), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1037), .A2(new_n588), .A3(new_n1041), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n913), .A2(new_n928), .ZN(new_n1060));
  INV_X1    g635(.A(new_n927), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n916), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n920), .A2(new_n925), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n932), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n930), .A2(KEYINPUT121), .A3(new_n932), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n980), .A2(new_n1012), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT123), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n980), .A2(new_n1012), .A3(new_n981), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1068), .A2(new_n1072), .A3(new_n1073), .A4(new_n957), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1016), .A2(new_n1059), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n679), .A2(new_n983), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT108), .ZN(new_n1077));
  OR3_X1    g652(.A1(new_n1077), .A2(new_n1002), .A3(new_n1001), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1078), .A2(new_n995), .B1(new_n991), .B2(new_n1006), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n913), .A2(G168), .ZN(new_n1080));
  OR3_X1    g655(.A1(new_n1011), .A2(new_n1080), .A3(KEYINPUT63), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1009), .B1(new_n1081), .B2(new_n980), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n977), .A2(new_n978), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OR3_X1    g659(.A1(new_n1084), .A2(new_n1009), .A3(new_n1080), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1079), .B(new_n1082), .C1(KEYINPUT63), .C2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT62), .B1(new_n933), .B2(new_n934), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1066), .A2(new_n1088), .A3(new_n1067), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n956), .A2(G171), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT125), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1087), .A2(new_n1089), .A3(new_n1091), .A4(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1075), .A2(new_n1086), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(new_n758), .B(G2067), .Z(new_n1097));
  XNOR2_X1  g672(.A(new_n726), .B(new_n1044), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n696), .B2(new_n694), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n696), .B2(new_n694), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n576), .A2(new_n672), .A3(new_n577), .ZN(new_n1102));
  NAND2_X1  g677(.A1(G290), .A2(G1986), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n895), .A2(new_n990), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1096), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1044), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n1108), .B(KEYINPUT46), .Z(new_n1109));
  NAND2_X1  g684(.A1(new_n1097), .A2(new_n727), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n1105), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT47), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1105), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n694), .A2(new_n696), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1099), .A2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n758), .A2(G2067), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1101), .A2(new_n1113), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT126), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1102), .A2(new_n1113), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT48), .Z(new_n1121));
  AOI211_X1 g696(.A(new_n1112), .B(new_n1117), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1107), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g698(.A1(G227), .A2(new_n459), .ZN(new_n1125));
  NOR2_X1   g699(.A1(new_n1125), .A2(KEYINPUT127), .ZN(new_n1126));
  NOR3_X1   g700(.A1(G401), .A2(G229), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g701(.A1(new_n1125), .A2(KEYINPUT127), .ZN(new_n1128));
  NAND4_X1  g702(.A1(new_n872), .A2(new_n833), .A3(new_n1127), .A4(new_n1128), .ZN(G225));
  INV_X1    g703(.A(G225), .ZN(G308));
endmodule


