//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n465), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI211_X1 g045(.A(new_n466), .B(new_n467), .C1(G2105), .C2(new_n470), .ZN(G160));
  INV_X1    g046(.A(new_n461), .ZN(new_n472));
  INV_X1    g047(.A(new_n460), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n459), .B1(new_n473), .B2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n460), .B2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n483), .B(KEYINPUT4), .C1(new_n461), .C2(new_n460), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n486), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n489), .A2(new_n487), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(new_n486), .A4(new_n490), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  NAND2_X1  g072(.A1(KEYINPUT69), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(KEYINPUT69), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(new_n504), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n509), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n505), .A2(new_n515), .ZN(G166));
  AND2_X1   g091(.A1(new_n502), .A2(new_n512), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  INV_X1    g093(.A(new_n501), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT5), .B1(KEYINPUT69), .B2(G543), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n500), .A2(new_n522), .A3(new_n501), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n521), .A2(new_n523), .A3(G63), .A4(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n510), .A2(G51), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n518), .A2(new_n524), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n523), .A3(G64), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n533), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n510), .A2(G43), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n521), .A2(new_n523), .A3(G56), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n504), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI211_X1 g123(.A(KEYINPUT71), .B(new_n504), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n510), .A2(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT72), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n510), .A2(new_n558), .A3(G53), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(KEYINPUT72), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n517), .A2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n519), .A2(new_n520), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n568), .ZN(G299));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n510), .A2(G49), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(KEYINPUT73), .A3(G49), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n573), .A2(new_n574), .B1(new_n517), .B2(G87), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n521), .A2(new_n523), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n576), .B2(G74), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n577), .A3(KEYINPUT74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n565), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n510), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n502), .A2(G86), .A3(new_n512), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n517), .A2(KEYINPUT75), .A3(G86), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n576), .A2(G60), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n504), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n510), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  NAND3_X1  g175(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n513), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n565), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G284));
  XNOR2_X1  g188(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  AND4_X1   g190(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n568), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  AND2_X1   g193(.A1(new_n605), .A2(new_n609), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NOR2_X1   g196(.A1(new_n550), .A2(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g201(.A(KEYINPUT3), .B(G2104), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n464), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n474), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n476), .A2(G123), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n636), .A2(KEYINPUT78), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(KEYINPUT78), .B2(new_n636), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT80), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT81), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(KEYINPUT81), .ZN(new_n654));
  OAI22_X1  g229(.A1(new_n653), .A2(new_n654), .B1(new_n650), .B2(new_n648), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n655), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n646), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n662), .A2(new_n645), .A3(new_n658), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n661), .B2(new_n663), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT18), .Z(new_n675));
  INV_X1    g250(.A(new_n672), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n673), .B1(new_n676), .B2(new_n670), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n670), .B(new_n678), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n677), .B1(new_n679), .B2(new_n676), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n676), .A3(new_n673), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n631), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT84), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT85), .ZN(new_n687));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n690), .A2(new_n691), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n697), .B(new_n696), .S(new_n689), .Z(new_n698));
  OR3_X1    g273(.A1(new_n695), .A2(new_n698), .A3(G1981), .ZN(new_n699));
  OAI21_X1  g274(.A(G1981), .B1(new_n695), .B2(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n700), .A3(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(G1986), .B1(new_n699), .B2(new_n700), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n687), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(new_n687), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n701), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n704), .A2(new_n707), .A3(new_n709), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(G229));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n640), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(KEYINPUT96), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT30), .B(G28), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT31), .A2(G11), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n718), .A2(new_n714), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G21), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G168), .B2(new_n723), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n716), .B(new_n722), .C1(G1966), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(G5), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G171), .B2(new_n723), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n726), .B1(G1966), .B2(new_n725), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT98), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n714), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2084), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n714), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT26), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G129), .B2(new_n476), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n739), .B1(new_n744), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n748));
  NAND2_X1  g323(.A1(G103), .A2(G2104), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n474), .A2(G139), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n627), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n459), .B2(new_n753), .ZN(new_n754));
  MUX2_X1   g329(.A(G33), .B(new_n754), .S(G29), .Z(new_n755));
  AOI21_X1  g330(.A(new_n747), .B1(G2072), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n745), .A2(new_n746), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n756), .B(new_n757), .C1(G2072), .C2(new_n755), .ZN(new_n758));
  INV_X1    g333(.A(G2090), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n714), .A2(G35), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n714), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  AOI211_X1 g337(.A(new_n738), .B(new_n758), .C1(new_n759), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n723), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n550), .B2(new_n723), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G1341), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n714), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT28), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n474), .A2(G140), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n476), .A2(G128), .ZN(new_n770));
  OR2_X1    g345(.A1(G104), .A2(G2105), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n771), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n768), .B1(new_n774), .B2(new_n714), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT95), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n729), .A2(new_n730), .B1(G1341), .B2(new_n765), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n763), .A2(new_n766), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n762), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n619), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G4), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT93), .B(G1348), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n780), .A2(G2090), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n723), .A2(G20), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT100), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n616), .B2(new_n723), .ZN(new_n789));
  INV_X1    g364(.A(G1956), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n785), .B(new_n791), .C1(new_n782), .C2(new_n784), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n714), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT99), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2078), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n732), .A2(new_n779), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n474), .A2(G131), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT86), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G107), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n476), .B2(G119), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT87), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G29), .ZN(new_n808));
  INV_X1    g383(.A(G25), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(G29), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n813), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n808), .A2(new_n811), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT88), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n815), .B1(new_n808), .B2(new_n811), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n810), .B(new_n813), .C1(new_n807), .C2(G29), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n723), .A2(G24), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n599), .B2(new_n723), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G1986), .Z(new_n824));
  AND3_X1   g399(.A1(new_n817), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n826));
  INV_X1    g401(.A(G6), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n827), .A2(G16), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G305), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT32), .B(G1981), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n723), .A2(G23), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n578), .B2(G16), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT33), .B(G1976), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT90), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n723), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n723), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(G1971), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(G1971), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n840), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n834), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n831), .A2(new_n832), .A3(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n837), .A2(new_n839), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n835), .A2(new_n845), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT91), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n845), .A2(new_n848), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n852), .A2(KEYINPUT91), .A3(new_n835), .A4(new_n847), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n825), .B(new_n826), .C1(new_n854), .C2(KEYINPUT34), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT34), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n817), .A2(new_n821), .A3(new_n824), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT92), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT36), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n798), .B1(new_n862), .B2(new_n864), .ZN(G311));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n863), .B1(new_n859), .B2(new_n860), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n797), .B1(new_n866), .B2(new_n867), .ZN(G150));
  NOR2_X1   g443(.A1(new_n610), .A2(new_n620), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n521), .A2(new_n523), .A3(G67), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G651), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n510), .A2(G55), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n513), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT101), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n504), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n881), .A2(new_n882), .A3(new_n878), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n880), .A2(new_n883), .B1(new_n548), .B2(new_n549), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n544), .A2(new_n545), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(G651), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n542), .B1(new_n886), .B2(KEYINPUT71), .ZN(new_n887));
  INV_X1    g462(.A(new_n549), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n875), .A4(new_n879), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n871), .B(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(KEYINPUT39), .ZN(new_n893));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(G860), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n875), .A2(KEYINPUT101), .A3(new_n879), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n882), .B1(new_n881), .B2(new_n878), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n899), .ZN(G145));
  XNOR2_X1  g475(.A(G160), .B(new_n640), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n480), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n754), .B(new_n744), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n474), .A2(G142), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n476), .A2(G130), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n459), .A2(G118), .ZN(new_n907));
  OAI21_X1  g482(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n904), .B(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(new_n773), .B(new_n491), .Z(new_n911));
  OR2_X1    g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n805), .B(new_n629), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n903), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  INV_X1    g494(.A(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n902), .A4(new_n915), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT105), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n918), .A2(new_n922), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g504(.A(new_n611), .B1(new_n880), .B2(new_n883), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n623), .B(KEYINPUT106), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n888), .A2(new_n887), .B1(new_n896), .B2(new_n897), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n548), .A2(new_n549), .A3(new_n881), .A4(new_n878), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n931), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT107), .B1(new_n619), .B2(G299), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n616), .A2(new_n937), .A3(new_n610), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n619), .A2(G299), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n940), .A2(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(KEYINPUT41), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n599), .B(G303), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n578), .B(G305), .Z(new_n947));
  XNOR2_X1  g522(.A(new_n946), .B(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT42), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n945), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n930), .B1(new_n950), .B2(new_n611), .ZN(G295));
  OAI21_X1  g526(.A(new_n930), .B1(new_n950), .B2(new_n611), .ZN(G331));
  INV_X1    g527(.A(new_n948), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n533), .A2(KEYINPUT108), .A3(new_n537), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n504), .B1(new_n530), .B2(new_n531), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n536), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(G168), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(G301), .A2(new_n955), .A3(G286), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n932), .B2(new_n933), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n940), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n884), .A2(new_n889), .A3(new_n959), .A4(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  INV_X1    g540(.A(new_n960), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n934), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n962), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n961), .A2(new_n963), .ZN(new_n970));
  OAI22_X1  g545(.A1(new_n968), .A2(new_n969), .B1(new_n944), .B2(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(KEYINPUT110), .B(new_n962), .C1(new_n964), .C2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n953), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n961), .A2(new_n963), .A3(new_n940), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n965), .B1(new_n934), .B2(new_n966), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n963), .A2(KEYINPUT109), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n961), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n940), .B(KEYINPUT41), .Z(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G37), .B1(new_n980), .B2(new_n948), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n973), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n981), .B(KEYINPUT43), .C1(new_n948), .C2(new_n980), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n982), .B2(KEYINPUT43), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n980), .B2(new_n948), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n967), .A2(new_n964), .B1(new_n890), .B2(new_n960), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n974), .B1(new_n991), .B2(new_n944), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n923), .B1(new_n992), .B2(new_n953), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT43), .B1(new_n992), .B2(new_n953), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n981), .A2(new_n995), .A3(KEYINPUT111), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n988), .A2(new_n997), .A3(KEYINPUT112), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT112), .B1(new_n988), .B2(new_n997), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n987), .B1(new_n998), .B2(new_n999), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n491), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G40), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n470), .B2(G2105), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n462), .A2(new_n465), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT67), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n465), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n467), .A2(new_n466), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT113), .A3(new_n1006), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1004), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n773), .B(G2067), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT116), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n742), .B2(new_n743), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT115), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n744), .B2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n805), .B(new_n815), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1016), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n1016), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n807), .A2(new_n815), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT125), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1025), .A2(new_n1032), .B1(G2067), .B2(new_n773), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1027), .A2(new_n1030), .B1(new_n1033), .B2(new_n1016), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1024), .B(KEYINPUT46), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1016), .B1(new_n744), .B2(new_n1017), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT126), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1038), .A2(KEYINPUT47), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT47), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT113), .B1(new_n1014), .B2(new_n1006), .ZN(new_n1045));
  AND4_X1   g620(.A1(KEYINPUT113), .A2(new_n1006), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g622(.A(new_n490), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT4), .B1(new_n627), .B2(new_n483), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n1050), .B2(new_n493), .ZN(new_n1051));
  OAI22_X1  g626(.A1(new_n1045), .A2(new_n1046), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g627(.A(KEYINPUT50), .B(G1384), .C1(new_n492), .C2(new_n495), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n790), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n1055));
  NAND3_X1  g630(.A1(G299), .A2(new_n1055), .A3(KEYINPUT57), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n568), .A2(new_n562), .A3(new_n563), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1055), .A2(KEYINPUT57), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1055), .A2(KEYINPUT57), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1057), .A2(new_n560), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n494), .B1(new_n1050), .B2(new_n493), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n486), .A2(new_n490), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n489), .A2(new_n487), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(KEYINPUT68), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1001), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1003), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1013), .A2(new_n1015), .B1(new_n1051), .B2(KEYINPUT45), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1054), .A2(new_n1061), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1051), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(G2067), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1045), .A2(new_n1046), .B1(KEYINPUT50), .B2(new_n1002), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1047), .B1(new_n496), .B2(new_n1001), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n783), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n610), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1061), .B1(new_n1054), .B2(new_n1070), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1071), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1054), .A2(new_n1061), .A3(new_n1070), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1078), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1061), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1047), .B1(new_n491), .B2(new_n1001), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n496), .A2(new_n1047), .A3(new_n1001), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1956), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1083), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT61), .A3(new_n1071), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  INV_X1    g666(.A(new_n783), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1066), .A2(KEYINPUT50), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n491), .A2(new_n1047), .A3(new_n1001), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1072), .A2(G2067), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1091), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1073), .A2(new_n1076), .A3(KEYINPUT60), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(new_n1099), .A3(new_n619), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1082), .A2(new_n1090), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1051), .A2(KEYINPUT45), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT45), .B1(new_n496), .B2(new_n1001), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1103), .A2(new_n1104), .A3(G1996), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT58), .B(G1341), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1051), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n550), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT59), .B(new_n550), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(new_n619), .C2(new_n1099), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1079), .B1(new_n1101), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g690(.A(G1971), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1093), .A2(new_n759), .A3(new_n1095), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G303), .A2(G8), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT55), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1117), .A2(new_n1118), .A3(new_n1115), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1120), .A2(G8), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G8), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1107), .B2(new_n1051), .ZN(new_n1127));
  INV_X1    g702(.A(G1976), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n580), .A2(new_n1128), .A3(new_n581), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n575), .A2(new_n577), .A3(G1976), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1072), .A2(G8), .A3(new_n1131), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT52), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n586), .A2(G651), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n510), .A2(G48), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n588), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(G1981), .ZN(new_n1138));
  INV_X1    g713(.A(G1981), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n587), .A2(new_n1139), .A3(new_n590), .A4(new_n591), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1140), .A3(KEYINPUT49), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1127), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1132), .A2(new_n1134), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1971), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1086), .A2(new_n759), .A3(new_n1087), .ZN(new_n1149));
  OAI21_X1  g724(.A(G8), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1122), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1125), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1074), .A2(new_n1075), .A3(G2084), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1013), .A2(new_n1015), .B1(new_n1003), .B2(new_n1002), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1155));
  AOI21_X1  g730(.A(G1966), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(G8), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(G286), .A2(G8), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1158), .B2(KEYINPUT122), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1155), .A2(new_n1107), .A3(new_n1004), .ZN(new_n1163));
  INV_X1    g738(.A(G1966), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G2084), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1093), .A2(new_n1166), .A3(new_n1095), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(G8), .B(new_n1160), .C1(new_n1168), .C2(G286), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1162), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(G8), .A3(G286), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT53), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n1173), .B2(G2078), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n730), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1172), .A2(new_n1005), .A3(G2078), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1014), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n459), .B1(new_n470), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1178), .B2(new_n470), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1102), .A2(new_n1177), .A3(new_n1004), .A4(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1174), .A2(new_n1175), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G301), .B(KEYINPUT54), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1163), .A2(new_n1172), .A3(G2078), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n1183), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1170), .A2(new_n1171), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1114), .A2(new_n1152), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  AOI211_X1 g765(.A(new_n1126), .B(G286), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1151), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1146), .B1(new_n1192), .B2(new_n1125), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1124), .A2(G8), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1122), .B1(new_n1194), .B2(new_n1119), .ZN(new_n1195));
  OAI211_X1 g770(.A(G8), .B(G168), .C1(new_n1153), .C2(new_n1156), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1146), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1190), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT120), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n582), .A2(new_n1128), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1138), .A2(new_n1140), .A3(KEYINPUT49), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT49), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1203), .B2(new_n1127), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1140), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1145), .A2(new_n1128), .A3(new_n582), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1207), .A2(KEYINPUT120), .A3(new_n1140), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1127), .B(KEYINPUT119), .Z(new_n1209));
  AND3_X1   g784(.A1(new_n1206), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1193), .A2(new_n1198), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1189), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1212), .B1(new_n1189), .B2(new_n1211), .ZN(new_n1214));
  AND2_X1   g789(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1215));
  AOI21_X1  g790(.A(G301), .B1(new_n1215), .B2(new_n1186), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1152), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n1218));
  AND3_X1   g793(.A1(new_n1170), .A2(new_n1218), .A3(new_n1171), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1218), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NOR3_X1   g796(.A1(new_n1213), .A2(new_n1214), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(new_n1028), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT114), .ZN(new_n1224));
  NAND2_X1  g799(.A1(G290), .A2(G1986), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1226), .B(new_n1016), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1027), .A2(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1228), .B(KEYINPUT117), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1044), .B1(new_n1222), .B2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g805(.A1(new_n711), .A2(new_n712), .ZN(new_n1232));
  INV_X1    g806(.A(G319), .ZN(new_n1233));
  NOR2_X1   g807(.A1(G227), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g808(.A1(new_n1232), .A2(new_n668), .A3(KEYINPUT127), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g809(.A(KEYINPUT127), .ZN(new_n1236));
  OAI21_X1  g810(.A(new_n1234), .B1(new_n666), .B2(new_n667), .ZN(new_n1237));
  OAI21_X1  g811(.A(new_n1236), .B1(G229), .B2(new_n1237), .ZN(new_n1238));
  AOI22_X1  g812(.A1(new_n1235), .A2(new_n1238), .B1(new_n925), .B2(new_n927), .ZN(new_n1239));
  AND2_X1   g813(.A1(new_n984), .A2(new_n986), .ZN(new_n1240));
  AND2_X1   g814(.A1(new_n1239), .A2(new_n1240), .ZN(G308));
  NAND2_X1  g815(.A1(new_n1239), .A2(new_n1240), .ZN(G225));
endmodule


