//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n194), .A2(KEYINPUT74), .A3(G146), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(G146), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT74), .B1(new_n194), .B2(G146), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(G119), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  OR2_X1    g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G128), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n201), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT73), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n206), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n193), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n197), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n203), .A2(new_n204), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(G110), .B2(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT75), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT75), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n218), .B(new_n221), .C1(G110), .C2(new_n211), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n227));
  XOR2_X1   g041(.A(new_n225), .B(new_n227), .Z(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n206), .A2(new_n213), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n223), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n232), .A3(new_n188), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n229), .A2(new_n232), .A3(KEYINPUT25), .A4(new_n188), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n190), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n232), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n189), .A2(G902), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n242));
  INV_X1    g056(.A(G221), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT9), .B(G234), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n243), .B1(new_n245), .B2(new_n188), .ZN(new_n246));
  INV_X1    g060(.A(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g063(.A(G107), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G104), .ZN(new_n251));
  INV_X1    g065(.A(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(G107), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n248), .A2(new_n251), .A3(new_n252), .A4(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n247), .A2(G107), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n250), .A2(G104), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(G143), .B(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G128), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n215), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n258), .B1(G128), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n254), .B(new_n257), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n257), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n259), .B1(G143), .B2(new_n215), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n200), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n271), .A3(new_n260), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G137), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT11), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT64), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(G137), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n282), .A2(new_n283), .B1(KEYINPUT64), .B2(new_n278), .ZN(new_n284));
  OAI21_X1  g098(.A(G131), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n279), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n281), .A2(G134), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n279), .B1(new_n275), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G131), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n271), .B2(new_n260), .ZN(new_n296));
  INV_X1    g110(.A(new_n266), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n265), .A2(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n292), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n248), .A2(new_n251), .A3(new_n253), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G101), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n254), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n262), .A2(new_n268), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n262), .B2(new_n268), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n258), .B2(new_n304), .ZN(new_n311));
  INV_X1    g125(.A(new_n304), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n269), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(KEYINPUT66), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n300), .A2(new_n315), .A3(G101), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n302), .A2(new_n310), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n298), .A2(new_n299), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT12), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n273), .A2(new_n319), .A3(new_n292), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n294), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(G110), .B(G140), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n226), .A2(G227), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n265), .A2(new_n295), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n296), .A2(new_n297), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n317), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n292), .ZN(new_n329));
  INV_X1    g143(.A(new_n324), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(new_n318), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n188), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G469), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT76), .B(G469), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n330), .B1(new_n329), .B2(new_n318), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n336), .A2(new_n337), .B1(new_n321), .B2(new_n324), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n328), .A2(new_n292), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n299), .B1(new_n298), .B2(new_n317), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n324), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n188), .B(new_n335), .C1(new_n338), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n246), .B1(new_n334), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G214), .B1(G237), .B2(G902), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n208), .A2(G116), .ZN(new_n347));
  INV_X1    g161(.A(G116), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT2), .B(G113), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n302), .A2(new_n352), .A3(new_n316), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G122), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n350), .A2(new_n351), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n208), .A3(G116), .ZN(new_n357));
  OAI211_X1 g171(.A(G113), .B(new_n357), .C1(new_n350), .C2(new_n356), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n297), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n354), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n271), .A2(new_n260), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n191), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n311), .A2(new_n313), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G224), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G953), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT7), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n354), .B(KEYINPUT8), .ZN(new_n371));
  AND4_X1   g185(.A1(new_n355), .A2(new_n358), .A3(new_n254), .A4(new_n257), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n355), .A2(new_n358), .B1(new_n254), .B2(new_n257), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n362), .B(new_n364), .C1(new_n368), .C2(new_n367), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n360), .A2(new_n370), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n188), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(new_n365), .B(new_n367), .Z(new_n380));
  NAND2_X1  g194(.A1(new_n353), .A2(new_n359), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n382));
  INV_X1    g196(.A(new_n354), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n383), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n376), .A2(KEYINPUT78), .A3(new_n188), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G210), .B1(G237), .B2(G902), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT79), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n391), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n379), .A2(new_n387), .A3(new_n393), .A4(new_n388), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n346), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n344), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G475), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n198), .A2(new_n197), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(new_n195), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n196), .A2(KEYINPUT81), .A3(new_n197), .A4(new_n198), .ZN(new_n402));
  NOR2_X1   g216(.A1(G237), .A2(G953), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(G143), .A3(G214), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G143), .B1(new_n403), .B2(G214), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(G131), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n290), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n401), .A2(new_n402), .A3(new_n409), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G113), .B(G122), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n247), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n290), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n407), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n193), .B(new_n215), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT80), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n423), .A3(new_n418), .ZN(new_n424));
  OAI21_X1  g238(.A(KEYINPUT80), .B1(new_n407), .B2(new_n419), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n414), .A2(new_n427), .ZN(new_n430));
  INV_X1    g244(.A(new_n416), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI211_X1 g246(.A(KEYINPUT83), .B(new_n416), .C1(new_n414), .C2(new_n427), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n398), .B1(new_n434), .B2(new_n188), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G122), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G116), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n250), .B1(new_n438), .B2(KEYINPUT14), .ZN(new_n439));
  XNOR2_X1  g253(.A(G116), .B(G122), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n200), .A2(G143), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n202), .A2(G143), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n274), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n274), .B1(new_n442), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n441), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n443), .A2(KEYINPUT13), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT85), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n200), .A2(G143), .B1(KEYINPUT13), .B2(new_n443), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n274), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n348), .A2(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n438), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT84), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G107), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n250), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n445), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n448), .B1(new_n452), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n244), .A2(new_n187), .A3(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n448), .B(new_n463), .C1(new_n452), .C2(new_n461), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT86), .B1(new_n467), .B2(new_n188), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n469), .B(G902), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(G478), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n468), .A2(new_n470), .B1(KEYINPUT15), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(G234), .A2(G237), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(G952), .A3(new_n226), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(G898), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(G902), .A3(G953), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n471), .A2(KEYINPUT15), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n467), .A2(new_n188), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n472), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n193), .B(KEYINPUT19), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n197), .B1(new_n484), .B2(G146), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n410), .B2(new_n412), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n431), .B1(new_n486), .B2(new_n426), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n428), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT82), .B1(new_n428), .B2(new_n487), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(KEYINPUT20), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n488), .A2(KEYINPUT82), .A3(new_n493), .A4(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n436), .A2(new_n482), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n242), .B1(new_n397), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n436), .A2(new_n482), .A3(new_n495), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n396), .A2(new_n498), .A3(KEYINPUT87), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n403), .A2(G210), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT26), .B(G101), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n308), .A2(new_n303), .A3(new_n309), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT66), .B1(new_n311), .B2(new_n313), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n507), .B1(new_n510), .B2(new_n292), .ZN(new_n511));
  AND4_X1   g325(.A1(new_n507), .A2(new_n292), .A3(new_n310), .A4(new_n314), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n275), .B2(new_n288), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n361), .A2(new_n291), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(new_n352), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n506), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT69), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT30), .A4(new_n515), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n292), .A2(new_n310), .A3(new_n314), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT67), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n292), .A2(new_n507), .A3(new_n310), .A4(new_n314), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n515), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n292), .A2(new_n363), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n352), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n519), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT69), .B(new_n532), .C1(new_n521), .C2(new_n526), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n518), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT31), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n513), .A2(new_n517), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n529), .A2(new_n352), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT28), .B1(new_n517), .B2(new_n522), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n506), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n518), .B(new_n545), .C1(new_n534), .C2(new_n535), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT71), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT32), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n539), .B(new_n506), .C1(new_n534), .C2(new_n535), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n505), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT29), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n542), .B(KEYINPUT72), .Z(new_n557));
  INV_X1    g371(.A(new_n513), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n352), .B1(new_n558), .B2(new_n516), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n539), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n560), .B2(new_n538), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n505), .A2(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n188), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G472), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n241), .B(new_n500), .C1(new_n552), .C2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(G101), .ZN(G3));
  NOR2_X1   g381(.A1(new_n550), .A2(new_n551), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n547), .A2(new_n188), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G472), .ZN(new_n570));
  INV_X1    g384(.A(new_n241), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n334), .A2(new_n343), .ZN(new_n572));
  INV_X1    g386(.A(new_n246), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n395), .A2(new_n478), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n492), .A2(new_n494), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(new_n435), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n467), .B(KEYINPUT33), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n471), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT88), .B(G478), .C1(new_n467), .C2(new_n188), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT88), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n585), .B1(new_n480), .B2(new_n471), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n583), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(KEYINPUT89), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n578), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n577), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  NAND2_X1  g409(.A1(new_n472), .A2(new_n481), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n435), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n490), .B1(KEYINPUT90), .B2(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g413(.A1(KEYINPUT90), .A2(KEYINPUT20), .ZN(new_n600));
  MUX2_X1   g414(.A(new_n490), .B(new_n599), .S(new_n600), .Z(new_n601));
  XNOR2_X1  g415(.A(new_n478), .B(KEYINPUT91), .ZN(new_n602));
  AND4_X1   g416(.A1(new_n395), .A2(new_n598), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n577), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT35), .B(G107), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  NAND2_X1  g422(.A1(new_n235), .A2(new_n236), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n189), .ZN(new_n610));
  OR4_X1    g424(.A1(KEYINPUT36), .A2(new_n231), .A3(new_n223), .A4(new_n230), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n231), .A2(new_n223), .B1(KEYINPUT36), .B2(new_n230), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n611), .A2(new_n240), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT94), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n237), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n500), .A2(new_n568), .A3(new_n570), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT37), .B(G110), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT95), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n619), .B(new_n621), .ZN(G12));
  NAND2_X1  g436(.A1(new_n547), .A2(new_n549), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT71), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT32), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n565), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n618), .A2(new_n397), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n474), .B1(new_n477), .B2(G900), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n598), .A2(new_n601), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  XOR2_X1   g449(.A(new_n631), .B(KEYINPUT39), .Z(new_n636));
  NOR2_X1   g450(.A1(new_n574), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT96), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n534), .A2(new_n535), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n506), .B1(new_n640), .B2(new_n539), .ZN(new_n641));
  INV_X1    g455(.A(new_n560), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n188), .B1(new_n642), .B2(new_n505), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n627), .A2(new_n553), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n638), .A2(KEYINPUT40), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n392), .A2(new_n394), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT38), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n436), .A2(new_n495), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n596), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n610), .A2(new_n614), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n648), .A2(new_n650), .A3(new_n346), .A4(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n639), .A2(new_n645), .A3(new_n646), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT97), .B(G143), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G45));
  OAI211_X1 g469(.A(new_n587), .B(new_n631), .C1(new_n579), .C2(new_n435), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n630), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n552), .B2(new_n565), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  AND3_X1   g473(.A1(new_n294), .A2(new_n318), .A3(new_n320), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n341), .A2(KEYINPUT77), .B1(new_n660), .B2(new_n330), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n336), .A2(new_n337), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G469), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n343), .B(new_n573), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n629), .A2(new_n592), .A3(new_n241), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT41), .B(G113), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G15));
  NAND4_X1  g483(.A1(new_n629), .A2(new_n241), .A3(new_n603), .A4(new_n666), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G116), .ZN(G18));
  INV_X1    g485(.A(new_n343), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n341), .A2(KEYINPUT77), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n660), .A2(new_n330), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n662), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n664), .B1(new_n675), .B2(new_n188), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n677), .A2(new_n678), .A3(new_n573), .A4(new_n395), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n647), .A2(new_n345), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT98), .B1(new_n665), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(new_n496), .A3(new_n618), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n552), .B2(new_n565), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NOR2_X1   g499(.A1(new_n650), .A2(new_n680), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n666), .A3(new_n602), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n561), .A2(new_n506), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n537), .A2(new_n546), .A3(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n569), .A2(G472), .B1(new_n549), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n241), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n690), .A2(new_n693), .A3(new_n241), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n687), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n437), .ZN(G24));
  AOI21_X1  g510(.A(new_n656), .B1(new_n679), .B2(new_n681), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n651), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G125), .ZN(G27));
  NAND2_X1  g513(.A1(G469), .A2(G902), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT100), .Z(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n343), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n325), .B(KEYINPUT101), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(KEYINPUT102), .A3(G469), .A4(new_n331), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n325), .A2(KEYINPUT101), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n321), .B2(new_n324), .ZN(new_n708));
  OAI211_X1 g522(.A(G469), .B(new_n331), .C1(new_n706), .C2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n703), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n392), .A2(new_n573), .A3(new_n345), .A4(new_n394), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n656), .A2(KEYINPUT42), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n629), .A2(new_n241), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(KEYINPUT32), .B1(new_n547), .B2(new_n549), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n241), .B1(new_n565), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n656), .A2(new_n712), .A3(new_n713), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT42), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n290), .ZN(G33));
  INV_X1    g537(.A(new_n632), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n629), .A2(new_n241), .A3(new_n724), .A4(new_n714), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT103), .B(G134), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G36));
  NOR2_X1   g541(.A1(new_n647), .A2(new_n346), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n568), .A2(new_n570), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n651), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n733), .A3(new_n651), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n580), .A2(new_n587), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT43), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n729), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(KEYINPUT105), .C1(new_n740), .C2(new_n739), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n704), .A2(KEYINPUT45), .A3(new_n331), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n664), .B1(new_n332), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n701), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n343), .B1(new_n746), .B2(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n573), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n749), .A2(new_n636), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n739), .A2(new_n740), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n737), .B1(new_n732), .B2(new_n734), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n728), .B1(new_n754), .B2(KEYINPUT44), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n742), .A2(new_n751), .A3(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT106), .B(G137), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G39));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n749), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n749), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n629), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n656), .A2(new_n241), .A3(new_n729), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  INV_X1    g581(.A(G952), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n737), .A2(new_n474), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n729), .A2(new_n665), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(new_n718), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n768), .B(G953), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n474), .B(new_n737), .C1(new_n692), .C2(new_n694), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n682), .ZN(new_n777));
  INV_X1    g591(.A(new_n770), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n645), .A2(new_n571), .A3(new_n474), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n590), .A2(new_n591), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT48), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n772), .A2(KEYINPUT118), .A3(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n775), .A2(new_n777), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n677), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n573), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n786), .B1(new_n763), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n787), .B2(new_n763), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n728), .A3(new_n776), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n648), .A2(new_n346), .A3(new_n666), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n776), .A2(KEYINPUT50), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n692), .A2(new_n694), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n769), .A3(new_n791), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n792), .A2(new_n796), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n799), .A2(new_n801), .B1(KEYINPUT117), .B2(new_n800), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n779), .A2(new_n580), .A3(new_n588), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n769), .A2(new_n651), .A3(new_n690), .A4(new_n770), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n776), .B(new_n728), .C1(new_n763), .C2(new_n786), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT117), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n805), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n792), .A2(new_n796), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT51), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n784), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n689), .A2(new_n549), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n570), .A2(new_n697), .A3(new_n651), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n629), .B2(new_n633), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n610), .A2(new_n573), .A3(new_n614), .A4(new_n631), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT111), .B1(new_n817), .B2(new_n712), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n573), .A2(new_n631), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n237), .A2(new_n613), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n705), .A2(new_n711), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n703), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n686), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n553), .A2(new_n644), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n552), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n658), .A4(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n634), .A2(new_n658), .A3(new_n826), .A4(new_n698), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n813), .B(new_n827), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n667), .A2(new_n670), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT108), .B1(new_n580), .B2(new_n588), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT108), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n649), .A2(new_n837), .A3(new_n587), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n395), .A2(new_n602), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n568), .A3(new_n570), .A4(new_n575), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n566), .A2(new_n684), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n835), .A2(new_n843), .A3(new_n695), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n598), .A2(new_n495), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n840), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n619), .B1(new_n576), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n619), .B(KEYINPUT109), .C1(new_n576), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n570), .A2(new_n719), .A3(new_n651), .A4(new_n814), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n690), .A2(KEYINPUT110), .A3(new_n651), .A4(new_n719), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n601), .A2(new_n728), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n597), .A2(new_n631), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n858), .A2(new_n574), .A3(new_n435), .A4(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n629), .A2(new_n618), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n725), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n722), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n844), .A2(new_n852), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n833), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n827), .A2(new_n813), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n831), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n834), .A2(new_n864), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n828), .A2(new_n830), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n827), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n844), .A3(new_n852), .A4(new_n863), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT53), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n868), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n872), .A2(KEYINPUT114), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n834), .A2(new_n864), .A3(new_n867), .A4(KEYINPUT53), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n812), .A2(new_n875), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n768), .A2(new_n226), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n241), .A2(new_n573), .A3(new_n345), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n736), .B(new_n887), .C1(KEYINPUT49), .C2(new_n785), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT107), .Z(new_n889));
  OAI21_X1  g703(.A(new_n648), .B1(new_n785), .B2(KEYINPUT49), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n889), .A2(new_n645), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n886), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT119), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n886), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n895), .ZN(G75));
  NOR2_X1   g710(.A1(new_n226), .A2(G952), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n188), .B1(new_n880), .B2(new_n882), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(new_n391), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n386), .A2(new_n384), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n380), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT55), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n898), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n900), .B2(new_n904), .ZN(G51));
  AND3_X1   g720(.A1(new_n872), .A2(KEYINPUT114), .A3(new_n868), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT114), .B1(new_n872), .B2(new_n868), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n882), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n883), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n701), .B(KEYINPUT57), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n675), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n899), .A2(new_n743), .A3(new_n745), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n897), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  INV_X1    g731(.A(new_n488), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n897), .ZN(G60));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT59), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n911), .A2(new_n581), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n875), .A2(new_n883), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n581), .B1(new_n925), .B2(new_n923), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n926), .A3(new_n897), .ZN(G63));
  AND2_X1   g741(.A1(new_n611), .A2(new_n612), .ZN(new_n928));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n909), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n930), .B1(new_n880), .B2(new_n882), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n897), .B1(new_n937), .B2(new_n928), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n239), .B1(new_n909), .B2(new_n931), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n932), .A2(new_n898), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n942), .A2(KEYINPUT121), .A3(new_n939), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n936), .A3(new_n940), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT121), .B1(new_n942), .B2(new_n939), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n945), .A2(new_n946), .A3(new_n934), .A4(new_n933), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n944), .A2(new_n947), .ZN(G66));
  AND2_X1   g762(.A1(new_n844), .A2(new_n852), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n475), .B2(new_n366), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n901), .B1(G898), .B2(new_n226), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  AOI21_X1  g770(.A(new_n226), .B1(G227), .B2(G900), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n729), .B(new_n638), .C1(new_n845), .C2(new_n839), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(new_n629), .A3(new_n241), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT124), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n816), .A2(new_n658), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n653), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n961), .A2(new_n964), .A3(new_n766), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(G953), .B1(new_n757), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n527), .A2(new_n531), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(new_n483), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n958), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n751), .A2(new_n686), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n766), .B(new_n725), .C1(new_n718), .C2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(new_n722), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n757), .A2(new_n976), .A3(new_n962), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n757), .B2(new_n962), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n226), .B(new_n975), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n957), .A2(KEYINPUT126), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G72));
  INV_X1    g797(.A(new_n641), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  NAND4_X1  g800(.A1(new_n874), .A2(new_n554), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(KEYINPUT127), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n757), .A2(new_n967), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n949), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n987), .B(new_n898), .C1(new_n991), .C2(new_n984), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(new_n993));
  INV_X1    g807(.A(new_n949), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n554), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(G57));
endmodule


