//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT31), .B(G50gat), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G228gat), .ZN(new_n207));
  INV_X1    g006(.A(G233gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n213));
  INV_X1    g012(.A(G211gat), .ZN(new_n214));
  OR2_X1    g013(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n213), .B1(new_n217), .B2(KEYINPUT22), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT72), .A2(G218gat), .ZN(new_n220));
  OAI21_X1  g019(.A(G211gat), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT22), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT73), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(G197gat), .B(G204gat), .Z(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n212), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n212), .ZN(new_n228));
  AOI211_X1 g027(.A(new_n225), .B(new_n228), .C1(new_n218), .C2(new_n223), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n211), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n217), .A2(new_n213), .A3(KEYINPUT22), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT73), .B1(new_n221), .B2(new_n222), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n228), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n224), .A2(new_n226), .A3(new_n212), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT74), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  INV_X1    g036(.A(G141gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G148gat), .ZN(new_n239));
  INV_X1    g038(.A(G148gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G141gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G155gat), .B(G162gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G162gat), .ZN(new_n247));
  INV_X1    g046(.A(G155gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT78), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G155gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT2), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT79), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT79), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT78), .B(G155gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n255), .B(KEYINPUT2), .C1(new_n256), .C2(new_n247), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n246), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT76), .B(KEYINPUT2), .Z(new_n259));
  AND3_X1   g058(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT75), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT75), .B1(new_n239), .B2(new_n241), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n244), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n230), .A2(new_n236), .B1(new_n237), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n258), .A2(new_n264), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n237), .B1(new_n227), .B2(new_n229), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n210), .B1(new_n267), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT86), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n237), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n227), .A2(new_n229), .A3(new_n211), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT74), .B1(new_n234), .B2(new_n235), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT29), .B1(new_n234), .B2(new_n235), .ZN(new_n278));
  INV_X1    g077(.A(new_n265), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT86), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n210), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n273), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n258), .A2(new_n264), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n258), .B2(new_n264), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n278), .B2(KEYINPUT3), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n277), .A2(new_n289), .A3(new_n209), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n206), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  AOI211_X1 g091(.A(new_n205), .B(new_n290), .C1(new_n273), .C2(new_n283), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n204), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G227gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(new_n208), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT64), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G169gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n300), .A2(new_n305), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n304), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n297), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n320), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n315), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n310), .B1(new_n324), .B2(new_n306), .ZN(new_n325));
  OR3_X1    g124(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT23), .A3(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT25), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT27), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G183gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n335), .B2(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(G190gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n334), .A2(new_n336), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT28), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n310), .B1(KEYINPUT26), .B2(new_n306), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n346), .A3(new_n327), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n345), .A2(new_n347), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n330), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G127gat), .ZN(new_n352));
  INV_X1    g151(.A(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT1), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G113gat), .A2(G120gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n358), .B1(G113gat), .B2(G120gat), .ZN(new_n359));
  AND2_X1   g158(.A1(G113gat), .A2(G120gat), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n359), .A2(new_n360), .A3(G127gat), .ZN(new_n361));
  OAI21_X1  g160(.A(G134gat), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G127gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n355), .A2(new_n363), .A3(new_n356), .ZN(new_n364));
  INV_X1    g163(.A(G134gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n359), .A2(new_n360), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n352), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n318), .A2(new_n329), .B1(new_n344), .B2(new_n348), .ZN(new_n370));
  INV_X1    g169(.A(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n296), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT34), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n372), .A3(new_n296), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  XOR2_X1   g175(.A(G15gat), .B(G43gat), .Z(new_n377));
  XNOR2_X1  g176(.A(G71gat), .B(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n375), .B(KEYINPUT32), .C1(new_n376), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n376), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n374), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n381), .ZN(new_n386));
  INV_X1    g185(.A(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT70), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n374), .A2(new_n389), .A3(new_n384), .A4(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n282), .B1(new_n281), .B2(new_n210), .ZN(new_n392));
  AOI211_X1 g191(.A(KEYINPUT86), .B(new_n209), .C1(new_n277), .C2(new_n280), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n291), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n205), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n284), .A2(new_n206), .A3(new_n291), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n203), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n294), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n268), .A2(KEYINPUT80), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n258), .A2(new_n264), .A3(new_n285), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT3), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n266), .A2(new_n371), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n368), .A2(new_n258), .A3(new_n264), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n409), .B2(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(KEYINPUT82), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n368), .A2(new_n258), .A3(new_n264), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n405), .B(new_n410), .C1(KEYINPUT4), .C2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n286), .A2(new_n287), .A3(new_n368), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT5), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n368), .A2(new_n258), .A3(new_n264), .A4(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT83), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n413), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n421), .A2(new_n422), .B1(new_n403), .B2(new_n404), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT84), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT83), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n420), .A2(new_n426), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AND4_X1   g228(.A1(KEYINPUT84), .A2(new_n429), .A3(new_n405), .A4(new_n424), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n418), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(KEYINPUT6), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n431), .A2(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n418), .B(new_n435), .C1(new_n425), .C2(new_n430), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n431), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n436), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n350), .B2(new_n237), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n370), .A2(new_n446), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n236), .B(new_n230), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n446), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n350), .A2(new_n447), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n451), .B(new_n452), .C1(new_n275), .C2(new_n276), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n458), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT30), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(new_n463), .A3(new_n458), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n294), .A2(new_n391), .A3(new_n397), .A4(KEYINPUT88), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n400), .A2(new_n445), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT35), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n439), .A2(new_n443), .A3(new_n444), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n294), .A2(new_n397), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n385), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n387), .A2(new_n386), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n388), .A2(new_n390), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n472), .A2(new_n479), .A3(KEYINPUT35), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n468), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n391), .A2(KEYINPUT36), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n474), .A2(new_n476), .B1(new_n388), .B2(new_n390), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(new_n484), .B2(KEYINPUT36), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n454), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT37), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n459), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n458), .B1(new_n454), .B2(new_n486), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n450), .A2(new_n453), .A3(KEYINPUT87), .A4(KEYINPUT37), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n490), .A2(new_n461), .A3(new_n496), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n444), .A2(new_n439), .A3(new_n443), .A4(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  OR3_X1    g298(.A1(new_n416), .A2(new_n414), .A3(new_n407), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT39), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n429), .A2(new_n405), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n407), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n407), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n435), .B1(new_n504), .B2(KEYINPUT39), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n504), .A2(KEYINPUT39), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT39), .A3(new_n500), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(KEYINPUT40), .A3(new_n435), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n440), .A2(new_n464), .A3(new_n462), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n397), .B(new_n294), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n472), .ZN(new_n513));
  OAI221_X1 g312(.A(new_n485), .B1(new_n498), .B2(new_n512), .C1(new_n471), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n482), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G29gat), .ZN(new_n519));
  INV_X1    g318(.A(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n520), .B2(new_n517), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(KEYINPUT15), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT89), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n525), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT15), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n526), .A2(new_n522), .A3(KEYINPUT15), .A4(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G22gat), .Z(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(G1gat), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT90), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n535), .A2(new_n538), .A3(new_n543), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n547), .A3(new_n530), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n549), .A3(new_n544), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n532), .A2(new_n546), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT92), .B1(new_n542), .B2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n529), .A2(new_n530), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n542), .A2(KEYINPUT92), .A3(new_n544), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n551), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n557), .B(KEYINPUT13), .Z(new_n561));
  INV_X1    g360(.A(new_n556), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n551), .A2(new_n556), .A3(KEYINPUT18), .A4(new_n557), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n560), .A2(new_n564), .A3(new_n571), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(KEYINPUT93), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G57gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n586), .A2(G64gat), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT94), .B(G57gat), .Z(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(G64gat), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n580), .B1(KEYINPUT9), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n585), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT21), .ZN(new_n593));
  INV_X1    g392(.A(new_n555), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(new_n552), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT95), .B(KEYINPUT21), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n591), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT96), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n605), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n603), .B(new_n605), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n599), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n609), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n615), .A2(new_n616), .A3(new_n597), .A4(new_n598), .ZN(new_n617));
  XNOR2_X1  g416(.A(G134gat), .B(G162gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(G232gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n618), .B(new_n621), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G99gat), .B(G106gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  NAND2_X1  g424(.A1(G85gat), .A2(G92gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT7), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(KEYINPUT8), .A2(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n554), .B1(new_n635), .B2(KEYINPUT17), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n531), .A2(new_n547), .A3(new_n633), .A4(new_n634), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n636), .B(new_n637), .C1(new_n620), .C2(new_n619), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n623), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n641), .A2(new_n642), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  NAND3_X1  g447(.A1(new_n638), .A2(new_n643), .A3(new_n623), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n648), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n644), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n614), .A2(new_n617), .A3(new_n650), .A4(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(G230gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n208), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n625), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n592), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n635), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n633), .A2(new_n659), .A3(new_n592), .A4(new_n634), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT10), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n657), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n656), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n674), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n666), .A3(new_n671), .A4(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n654), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n515), .A2(new_n579), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n445), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n534), .ZN(G1324gat));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n465), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n539), .B2(new_n684), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n681), .B2(new_n485), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n479), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n681), .B2(new_n693), .ZN(G1326gat));
  NOR2_X1   g493(.A1(new_n681), .A2(new_n513), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AND2_X1   g496(.A1(new_n614), .A2(new_n617), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n648), .B1(new_n645), .B2(new_n649), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n652), .A2(new_n651), .A3(new_n644), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n698), .A2(new_n701), .A3(new_n679), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n515), .A2(new_n579), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n516), .A3(new_n469), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n482), .A2(new_n514), .A3(KEYINPUT107), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n467), .A2(KEYINPUT35), .B1(new_n471), .B2(new_n480), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n485), .B1(new_n498), .B2(new_n512), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n513), .B1(new_n445), .B2(new_n465), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n699), .B2(new_n700), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n653), .A2(new_n650), .A3(KEYINPUT108), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n707), .A2(new_n713), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n709), .A2(new_n712), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n721), .B2(new_n701), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n678), .B(KEYINPUT105), .ZN(new_n724));
  INV_X1    g523(.A(new_n698), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n575), .A3(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n726), .B(KEYINPUT106), .Z(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n445), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n706), .A2(new_n729), .ZN(G1328gat));
  NOR3_X1   g529(.A1(new_n703), .A2(G36gat), .A3(new_n465), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  OAI21_X1  g531(.A(G36gat), .B1(new_n728), .B2(new_n465), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1329gat));
  INV_X1    g533(.A(G43gat), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n485), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n723), .A2(new_n727), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n703), .B2(new_n479), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT47), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n739), .B(new_n742), .C1(new_n728), .C2(new_n736), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n513), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n723), .A2(new_n727), .A3(new_n746), .ZN(new_n747));
  OR2_X1    g546(.A1(KEYINPUT109), .A2(KEYINPUT48), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n515), .A2(new_n472), .A3(new_n579), .A4(new_n702), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n749), .A2(new_n745), .B1(KEYINPUT109), .B2(KEYINPUT48), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n748), .B1(new_n747), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1331gat));
  NOR3_X1   g552(.A1(new_n724), .A2(new_n575), .A3(new_n654), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n707), .A2(new_n713), .A3(new_n469), .A4(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(KEYINPUT110), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n756), .A2(new_n588), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n588), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1332gat));
  NAND3_X1  g559(.A1(new_n707), .A2(new_n713), .A3(new_n754), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n707), .A2(new_n713), .A3(new_n763), .A4(new_n754), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n762), .A2(new_n470), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT49), .B(G64gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1333gat));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n485), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n762), .A2(new_n764), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n761), .B2(new_n479), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n772), .A2(KEYINPUT50), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT50), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1334gat));
  NAND3_X1  g575(.A1(new_n762), .A2(new_n472), .A3(new_n764), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n698), .A2(new_n575), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n679), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n720), .B2(new_n722), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n445), .ZN(new_n783));
  INV_X1    g582(.A(new_n701), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n515), .A2(KEYINPUT51), .A3(new_n784), .A4(new_n779), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n784), .B(new_n779), .C1(new_n709), .C2(new_n712), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n469), .A2(new_n629), .A3(new_n679), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n783), .B1(new_n790), .B2(new_n791), .ZN(G1336gat));
  INV_X1    g591(.A(new_n724), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n630), .A3(new_n470), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT112), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g595(.A(new_n465), .B(new_n780), .C1(new_n720), .C2(new_n722), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n797), .B2(new_n630), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n795), .B(KEYINPUT113), .Z(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n788), .B2(new_n785), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n470), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n782), .B2(new_n485), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n479), .A2(G99gat), .A3(new_n678), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n790), .B2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(G106gat), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n781), .B2(new_n472), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n513), .A2(G106gat), .A3(new_n724), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n789), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT53), .B1(new_n809), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n513), .B(new_n780), .C1(new_n720), .C2(new_n722), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n814), .B(new_n811), .C1(new_n815), .C2(new_n808), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n661), .A2(new_n662), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT10), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n656), .A3(new_n664), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n666), .A3(KEYINPUT54), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n657), .C1(new_n663), .C2(new_n665), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n672), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n677), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n822), .A2(new_n672), .A3(new_n824), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n562), .A2(new_n563), .A3(new_n561), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n557), .B1(new_n551), .B2(new_n556), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n570), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n574), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n827), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n718), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n827), .A2(new_n575), .A3(new_n830), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n679), .A2(new_n834), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n717), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n725), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n698), .A2(new_n701), .A3(new_n678), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n575), .ZN(new_n843));
  INV_X1    g642(.A(new_n575), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n680), .A2(KEYINPUT114), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n445), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n465), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n400), .A2(new_n466), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n353), .A3(new_n575), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n472), .A2(new_n479), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n853), .A3(new_n579), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(G113gat), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n854), .B2(G113gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n852), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  AOI21_X1  g658(.A(G120gat), .B1(new_n851), .B2(new_n679), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n849), .A2(new_n853), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n861), .A2(new_n354), .A3(new_n724), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(new_n862), .ZN(G1341gat));
  NAND3_X1  g662(.A1(new_n851), .A2(new_n363), .A3(new_n698), .ZN(new_n864));
  OAI21_X1  g663(.A(G127gat), .B1(new_n861), .B2(new_n725), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1342gat));
  NOR2_X1   g665(.A1(new_n470), .A2(new_n701), .ZN(new_n867));
  XNOR2_X1  g666(.A(KEYINPUT69), .B(G134gat), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n847), .A2(new_n850), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT56), .Z(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n861), .B2(new_n701), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1343gat));
  NAND3_X1  g671(.A1(new_n485), .A2(new_n469), .A3(new_n465), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n513), .B1(new_n840), .B2(new_n846), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n845), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n717), .A2(new_n827), .A3(new_n830), .A4(new_n834), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT55), .B1(new_n828), .B2(KEYINPUT116), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n822), .A2(new_n880), .A3(new_n672), .A4(new_n824), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n826), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n579), .A2(new_n882), .B1(new_n679), .B2(new_n834), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n878), .B1(new_n883), .B2(new_n784), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n877), .B1(new_n884), .B2(new_n725), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT57), .B1(new_n885), .B2(new_n513), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n876), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n579), .ZN(new_n888));
  OAI21_X1  g687(.A(G141gat), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n485), .A2(new_n472), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n847), .A2(new_n465), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n238), .A3(new_n579), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n887), .B2(new_n844), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n893), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n894), .B1(new_n896), .B2(new_n890), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n240), .A2(KEYINPUT59), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n887), .B2(new_n678), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n821), .A2(new_n666), .A3(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n824), .A2(new_n672), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT116), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n829), .A3(new_n881), .ZN(new_n903));
  INV_X1    g702(.A(new_n578), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT93), .B1(new_n573), .B2(new_n574), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n903), .B(new_n827), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n784), .B1(new_n906), .B2(new_n838), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n835), .A2(new_n701), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n725), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n842), .A2(new_n579), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n513), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT120), .B1(new_n912), .B2(KEYINPUT57), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n835), .A2(new_n701), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n915), .B1(new_n883), .B2(new_n784), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n916), .B2(new_n725), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n914), .B(new_n875), .C1(new_n917), .C2(new_n513), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n830), .A2(new_n677), .A3(new_n825), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n838), .B1(new_n920), .B2(new_n844), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n718), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n698), .B1(new_n922), .B2(new_n878), .ZN(new_n923));
  OAI211_X1 g722(.A(KEYINPUT57), .B(new_n472), .C1(new_n923), .C2(new_n877), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT119), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n840), .A2(new_n846), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n472), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n919), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n873), .A2(new_n678), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n240), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n899), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n892), .A2(new_n240), .A3(new_n679), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT117), .Z(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1345gat));
  NAND3_X1  g736(.A1(new_n892), .A2(new_n256), .A3(new_n698), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n887), .A2(new_n725), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n256), .ZN(G1346gat));
  OAI21_X1  g739(.A(G162gat), .B1(new_n887), .B2(new_n718), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n847), .A2(new_n247), .A3(new_n867), .A4(new_n891), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT121), .Z(G1347gat));
  AOI21_X1  g743(.A(new_n469), .B1(new_n840), .B2(new_n846), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n945), .A2(new_n470), .A3(new_n850), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n946), .A2(new_n301), .A3(new_n303), .A4(new_n575), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n469), .A2(new_n465), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n927), .A2(new_n853), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(G169gat), .B1(new_n949), .B2(new_n888), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1348gat));
  NAND3_X1  g750(.A1(new_n946), .A2(new_n305), .A3(new_n679), .ZN(new_n952));
  OAI21_X1  g751(.A(G176gat), .B1(new_n949), .B2(new_n724), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1349gat));
  INV_X1    g753(.A(new_n949), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n333), .B1(new_n955), .B2(new_n698), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n698), .A2(new_n342), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g757(.A(new_n958), .B(KEYINPUT60), .Z(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n949), .B2(new_n701), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT61), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n339), .A3(new_n717), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1351gat));
  NAND3_X1  g762(.A1(new_n891), .A2(KEYINPUT122), .A3(new_n470), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT122), .B1(new_n891), .B2(new_n470), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT123), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n966), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n968), .A2(new_n969), .A3(new_n945), .A4(new_n964), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n575), .ZN(new_n972));
  AOI22_X1  g771(.A1(new_n913), .A2(new_n918), .B1(new_n926), .B2(new_n928), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n948), .A2(new_n485), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n579), .A2(G197gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(G1352gat));
  NOR4_X1   g776(.A1(new_n965), .A2(G204gat), .A3(new_n678), .A4(new_n966), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT62), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n973), .A2(new_n724), .A3(new_n974), .ZN(new_n980));
  OAI21_X1  g779(.A(G204gat), .B1(new_n980), .B2(KEYINPUT124), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n793), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1353gat));
  NAND2_X1  g782(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n973), .A2(new_n725), .A3(new_n974), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n984), .B(new_n987), .C1(new_n988), .C2(new_n214), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n930), .A2(new_n485), .A3(new_n698), .A4(new_n948), .ZN(new_n990));
  NAND4_X1  g789(.A1(new_n990), .A2(new_n985), .A3(new_n986), .A4(G211gat), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n967), .A2(new_n214), .A3(new_n698), .A4(new_n970), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(G1354gat));
  NAND2_X1  g793(.A1(new_n215), .A2(new_n216), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n784), .A2(new_n995), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n973), .A2(new_n974), .A3(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n967), .A2(new_n717), .A3(new_n970), .ZN(new_n1000));
  INV_X1    g799(.A(G218gat), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(new_n1002), .ZN(new_n1004));
  OAI21_X1  g803(.A(KEYINPUT127), .B1(new_n1004), .B2(new_n997), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1355gat));
endmodule


