//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G137), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(G128), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n194), .B(new_n196), .C1(new_n197), .C2(KEYINPUT23), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G119), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n199), .A2(new_n196), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  OAI22_X1  g015(.A1(new_n198), .A2(G110), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n205), .A2(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n210), .A3(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n206), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT71), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n199), .A2(new_n196), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT24), .B(G110), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n198), .A2(G110), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n211), .ZN(new_n224));
  AOI21_X1  g038(.A(G146), .B1(new_n207), .B2(new_n210), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n214), .B(new_n215), .C1(new_n223), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n221), .B(new_n222), .C1(new_n225), .C2(new_n224), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n215), .B1(new_n229), .B2(new_n214), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n192), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n214), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n191), .ZN(new_n233));
  AOI21_X1  g047(.A(G902), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n187), .B1(new_n234), .B2(KEYINPUT73), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT73), .ZN(new_n236));
  INV_X1    g050(.A(new_n233), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(KEYINPUT72), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n227), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n239), .B2(new_n192), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n236), .B(KEYINPUT25), .C1(new_n240), .C2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G217), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(G234), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n235), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(G902), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT74), .Z(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n247), .B2(new_n240), .ZN(new_n248));
  NOR2_X1   g062(.A1(G472), .A2(G902), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  XOR2_X1   g064(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(G137), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT11), .A3(G134), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n257), .A3(new_n260), .A4(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XOR2_X1   g078(.A(KEYINPUT0), .B(G128), .Z(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n212), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(G143), .B(G146), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT0), .B(G128), .C1(new_n272), .C2(KEYINPUT64), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT2), .B(G113), .Z(new_n279));
  XNOR2_X1  g093(.A(G116), .B(G119), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n264), .A2(KEYINPUT67), .A3(new_n274), .A4(new_n275), .ZN(new_n283));
  AOI21_X1  g097(.A(G128), .B1(new_n267), .B2(new_n269), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n268), .A2(KEYINPUT1), .A3(G146), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT65), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n285), .B(new_n288), .C1(new_n272), .C2(G128), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT1), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n267), .A2(new_n269), .A3(new_n290), .A4(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n255), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n253), .A2(G137), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(new_n261), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n278), .A2(new_n282), .A3(new_n283), .A4(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n274), .A2(new_n262), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n297), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n281), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n251), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n275), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT66), .B1(new_n259), .B2(new_n261), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n271), .A2(new_n273), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n297), .A2(new_n282), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT28), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(G237), .A2(G953), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G210), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(KEYINPUT27), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G101), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT68), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n300), .A2(KEYINPUT30), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n278), .A2(new_n283), .A3(new_n297), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(KEYINPUT30), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n298), .B(new_n315), .C1(new_n319), .C2(new_n282), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n310), .A2(new_n316), .B1(new_n320), .B2(KEYINPUT31), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n276), .A2(new_n277), .B1(new_n292), .B2(new_n296), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n283), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n281), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n298), .A4(new_n315), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n250), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n298), .B1(new_n319), .B2(new_n282), .ZN(new_n329));
  INV_X1    g143(.A(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n302), .A2(new_n309), .A3(new_n316), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n318), .A2(new_n281), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(new_n298), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT70), .B(new_n335), .C1(new_n306), .C2(new_n307), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n330), .A2(new_n333), .ZN(new_n343));
  AOI21_X1  g157(.A(G902), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n328), .A2(KEYINPUT32), .B1(new_n345), .B2(G472), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n320), .A2(KEYINPUT31), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n316), .B1(new_n302), .B2(new_n309), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n327), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n249), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n248), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  AND4_X1   g168(.A1(G143), .A2(new_n354), .A3(new_n189), .A4(G214), .ZN(new_n355));
  AOI21_X1  g169(.A(G143), .B1(new_n311), .B2(G214), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n203), .A2(G125), .ZN(new_n359));
  OAI21_X1  g173(.A(G146), .B1(new_n208), .B2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n357), .A2(new_n358), .B1(new_n213), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT84), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n189), .A3(G214), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n268), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n311), .A2(G143), .A3(G214), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n358), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n362), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g182(.A(KEYINPUT84), .B(new_n358), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n361), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n361), .B(KEYINPUT85), .C1(new_n368), .C2(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(G104), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G131), .B1(new_n355), .B2(new_n356), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT17), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n364), .A2(new_n260), .A3(new_n365), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n207), .A2(new_n210), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n212), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT17), .B(G131), .C1(new_n355), .C2(new_n356), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n211), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n374), .A2(new_n377), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT88), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT19), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT19), .B1(new_n204), .B2(new_n206), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n390), .B(new_n212), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n211), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT19), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n395), .B1(new_n208), .B2(new_n359), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT19), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n390), .B1(new_n398), .B2(new_n212), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n389), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n212), .B1(new_n391), .B2(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT87), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n402), .A2(KEYINPUT88), .A3(new_n211), .A4(new_n393), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT86), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n378), .A2(new_n404), .A3(new_n380), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n378), .B2(new_n380), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n374), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n388), .B1(new_n409), .B2(new_n377), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT89), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n410), .A2(new_n411), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n377), .B1(new_n374), .B2(new_n408), .ZN(new_n416));
  AOI211_X1 g230(.A(new_n376), .B(new_n386), .C1(new_n372), .C2(new_n373), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n412), .B(new_n414), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT90), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT20), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n377), .B1(new_n374), .B2(new_n387), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n243), .B1(new_n423), .B2(new_n417), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT91), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(KEYINPUT91), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  OAI21_X1  g245(.A(G221), .B1(new_n431), .B2(G902), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n432), .B(KEYINPUT75), .Z(new_n433));
  INV_X1    g247(.A(G469), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(new_n243), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n189), .A2(G227), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n436), .B(new_n437), .Z(new_n438));
  NOR2_X1   g252(.A1(new_n284), .A2(new_n286), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT76), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n291), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n272), .A2(KEYINPUT76), .A3(new_n290), .A4(G128), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G104), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT3), .B1(new_n444), .B2(G107), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT3), .ZN(new_n446));
  INV_X1    g260(.A(G107), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G104), .ZN(new_n448));
  INV_X1    g262(.A(G101), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(G107), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n444), .A2(G107), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n447), .A2(G104), .ZN(new_n453));
  OAI21_X1  g267(.A(G101), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n443), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n445), .A2(new_n448), .A3(new_n450), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G101), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT4), .A3(new_n451), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n462), .A3(G101), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n274), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n264), .A2(new_n275), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n451), .A2(new_n454), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n457), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n292), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n458), .A2(new_n464), .A3(new_n465), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n456), .A2(new_n457), .B1(new_n292), .B2(new_n467), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n465), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n438), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n438), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n287), .A2(new_n466), .A3(new_n289), .A4(new_n291), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n456), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n303), .A2(new_n304), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT12), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n262), .A2(KEYINPUT12), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n456), .B2(new_n475), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n469), .B(new_n474), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n435), .B1(new_n482), .B2(new_n434), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n477), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n480), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT77), .B1(new_n486), .B2(new_n470), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n488), .B(new_n469), .C1(new_n478), .C2(new_n480), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n438), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n469), .A2(new_n474), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT78), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n458), .A2(new_n464), .A3(new_n468), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n477), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n469), .A2(KEYINPUT78), .A3(new_n474), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(G469), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n433), .B1(new_n483), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n305), .A2(G125), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT80), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n287), .A2(new_n289), .A3(new_n205), .A4(new_n291), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n305), .A2(new_n506), .A3(G125), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT81), .B(G224), .Z(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(G953), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n504), .A2(new_n505), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n503), .A2(new_n505), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n510), .B2(new_n509), .ZN(new_n514));
  XNOR2_X1  g328(.A(G110), .B(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT8), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n279), .A2(new_n280), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n451), .A3(new_n454), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n280), .A2(new_n519), .A3(KEYINPUT5), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n280), .B2(KEYINPUT5), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n195), .A3(G116), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT79), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n523), .A2(new_n195), .A3(KEYINPUT79), .A4(G116), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n526), .A2(G113), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n518), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n280), .A2(KEYINPUT5), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n530), .A2(G113), .A3(new_n526), .A4(new_n527), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n455), .B1(new_n517), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n516), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n281), .A2(new_n461), .A3(new_n463), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n455), .A2(new_n531), .A3(new_n517), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n515), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n512), .A2(new_n514), .A3(new_n533), .A4(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n537), .A2(new_n243), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  INV_X1    g353(.A(new_n515), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n536), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n509), .B(KEYINPUT82), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n504), .A2(new_n505), .A3(new_n507), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n545));
  INV_X1    g359(.A(new_n543), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n539), .A2(new_n548), .A3(new_n540), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n542), .A2(new_n544), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n502), .B1(new_n538), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n538), .A2(new_n550), .A3(new_n502), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n501), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n499), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G116), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n447), .B1(new_n557), .B2(KEYINPUT14), .ZN(new_n558));
  XNOR2_X1  g372(.A(G116), .B(G122), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n268), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n193), .A2(G143), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n253), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n253), .B1(new_n562), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n561), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(KEYINPUT93), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n560), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n562), .A2(new_n563), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n572), .A2(new_n253), .B1(G107), .B2(new_n559), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n559), .A2(G107), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n193), .A2(G143), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(KEYINPUT13), .B2(new_n563), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT92), .B1(new_n562), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n268), .A2(G128), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n580), .B(new_n562), .C1(new_n581), .C2(new_n577), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G134), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n573), .B(new_n574), .C1(new_n579), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n570), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n431), .A2(new_n242), .A3(G953), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n570), .A2(new_n588), .A3(new_n584), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT95), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT95), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n570), .A2(new_n588), .A3(new_n584), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n243), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(KEYINPUT15), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n595), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(G952), .A3(new_n189), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT21), .B(G898), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(G902), .A3(G953), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n430), .A2(new_n555), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n353), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n349), .B2(new_n243), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n350), .ZN(new_n613));
  INV_X1    g427(.A(new_n433), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n490), .A2(G469), .A3(new_n497), .ZN(new_n615));
  INV_X1    g429(.A(new_n481), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n474), .B1(new_n495), .B2(new_n469), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n434), .B(new_n243), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n435), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n614), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n613), .A2(new_n248), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n592), .A2(new_n623), .A3(new_n594), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n592), .A2(KEYINPUT96), .A3(new_n623), .A4(new_n594), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n590), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n596), .A2(G902), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n595), .A2(new_n596), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n628), .A2(KEYINPUT97), .A3(new_n629), .A4(new_n630), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n430), .A2(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n538), .A2(new_n550), .A3(new_n502), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n500), .B(new_n605), .C1(new_n638), .C2(new_n551), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n622), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G104), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n421), .A2(new_n418), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n425), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n639), .A2(new_n646), .A3(new_n599), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n622), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(new_n244), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n236), .B1(new_n240), .B2(G902), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n187), .ZN(new_n653));
  INV_X1    g467(.A(new_n247), .ZN(new_n654));
  INV_X1    g468(.A(new_n239), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n653), .A2(new_n241), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n613), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n607), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AOI21_X1  g476(.A(new_n658), .B1(new_n346), .B2(new_n352), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n604), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n601), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n645), .A2(new_n425), .A3(new_n598), .A4(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n500), .B1(new_n638), .B2(new_n551), .ZN(new_n667));
  OR3_X1    g481(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT99), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT99), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n621), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  AOI21_X1  g486(.A(KEYINPUT32), .B1(new_n349), .B2(new_n249), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n610), .A2(new_n243), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n336), .A2(new_n298), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n610), .B1(new_n675), .B2(new_n316), .ZN(new_n676));
  AOI211_X1 g490(.A(KEYINPUT100), .B(new_n674), .C1(new_n676), .C2(new_n320), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n320), .ZN(new_n679));
  INV_X1    g493(.A(new_n674), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n673), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n349), .A2(KEYINPUT32), .A3(new_n249), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n681), .A2(new_n677), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n352), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n638), .A2(new_n551), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n690), .B(KEYINPUT38), .Z(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n422), .A2(KEYINPUT91), .A3(new_n425), .ZN(new_n693));
  AOI21_X1  g507(.A(KEYINPUT91), .B1(new_n422), .B2(new_n425), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n658), .A2(new_n500), .A3(new_n598), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n689), .A2(new_n697), .A3(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n665), .B(KEYINPUT39), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n499), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT40), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT102), .B1(new_n689), .B2(new_n697), .ZN(new_n704));
  OR3_X1    g518(.A1(new_n703), .A2(KEYINPUT103), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT103), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n268), .ZN(G45));
  OAI211_X1 g522(.A(new_n636), .B(new_n665), .C1(new_n693), .C2(new_n694), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n555), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n663), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n345), .A2(G472), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n352), .A2(new_n713), .A3(new_n684), .ZN(new_n714));
  INV_X1    g528(.A(new_n248), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n243), .B1(new_n616), .B2(new_n617), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n614), .A3(new_n618), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT104), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n720), .A3(new_n614), .A4(new_n618), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n714), .A2(new_n715), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n430), .A2(new_n636), .A3(new_n640), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT41), .B(G113), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  INV_X1    g541(.A(new_n647), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT105), .B1(new_n723), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n353), .A2(new_n730), .A3(new_n647), .A4(new_n722), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR3_X1   g547(.A1(new_n693), .A2(new_n694), .A3(new_n606), .ZN(new_n734));
  INV_X1    g548(.A(new_n718), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n554), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n718), .B2(new_n667), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n658), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n714), .A2(new_n734), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  OAI21_X1  g556(.A(new_n316), .B1(new_n337), .B2(new_n341), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n347), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT107), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n347), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n327), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n611), .B1(new_n748), .B2(new_n249), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n599), .B1(new_n428), .B2(new_n429), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n719), .A2(new_n640), .A3(new_n721), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n749), .A2(new_n715), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  AOI211_X1 g567(.A(new_n658), .B(new_n611), .C1(new_n748), .C2(new_n249), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n709), .A2(KEYINPUT108), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n430), .A2(new_n756), .A3(new_n636), .A4(new_n665), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .A4(new_n739), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G125), .ZN(G27));
  NAND3_X1  g573(.A1(new_n552), .A2(new_n500), .A3(new_n553), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n690), .A2(new_n762), .A3(new_n500), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT42), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n621), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n755), .A2(new_n757), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n352), .A2(KEYINPUT110), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(new_n346), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n673), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n248), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n761), .A2(new_n499), .A3(new_n763), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n353), .A2(new_n755), .A3(new_n757), .A4(new_n773), .ZN(new_n774));
  AOI22_X1  g588(.A1(new_n767), .A2(new_n772), .B1(new_n774), .B2(new_n765), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n260), .ZN(G33));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n666), .B(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n714), .A2(new_n778), .A3(new_n773), .A4(new_n715), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  AND2_X1   g594(.A1(new_n490), .A2(new_n497), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n782));
  OAI21_X1  g596(.A(G469), .B1(new_n781), .B2(KEYINPUT45), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n435), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(KEYINPUT46), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n618), .B1(new_n785), .B2(KEYINPUT46), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n614), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n699), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n764), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n613), .A2(new_n740), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT43), .B1(new_n695), .B2(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n695), .A2(new_n636), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n792), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n790), .B(new_n791), .C1(new_n797), .C2(KEYINPUT44), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n256), .ZN(G39));
  INV_X1    g615(.A(KEYINPUT47), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n788), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT47), .B(new_n614), .C1(new_n786), .C2(new_n787), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR4_X1   g619(.A1(new_n709), .A2(new_n714), .A3(new_n715), .A4(new_n764), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  NOR3_X1   g622(.A1(new_n248), .A2(new_n501), .A3(new_n433), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n717), .A2(new_n618), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT49), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n692), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n689), .A2(new_n812), .A3(new_n794), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n749), .A2(new_n715), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n601), .B(new_n814), .C1(new_n795), .C2(new_n796), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n739), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n791), .A2(new_n735), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n689), .A2(new_n248), .A3(new_n601), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n637), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(G952), .A3(new_n189), .A4(new_n819), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n601), .B(new_n817), .C1(new_n795), .C2(new_n796), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n772), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT48), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(KEYINPUT121), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(KEYINPUT121), .B(KEYINPUT48), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n820), .B(new_n824), .C1(new_n822), .C2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n501), .B1(new_n827), .B2(KEYINPUT50), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n691), .A2(new_n718), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n815), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n827), .A2(KEYINPUT50), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n430), .A2(new_n636), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n821), .A2(new_n754), .B1(new_n818), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n810), .A2(new_n433), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n803), .A2(new_n804), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n815), .A2(new_n791), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n838), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n830), .A2(new_n831), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n835), .A2(new_n842), .A3(KEYINPUT51), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n837), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n835), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n826), .B(new_n844), .C1(new_n846), .C2(KEYINPUT51), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n657), .A2(new_n654), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n665), .B(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n245), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT117), .B1(new_n621), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n658), .A2(new_n499), .A3(new_n853), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n554), .B(new_n598), .C1(new_n693), .C2(new_n694), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n683), .B1(new_n682), .B2(new_n684), .ZN(new_n858));
  AND4_X1   g672(.A1(new_n683), .A2(new_n352), .A3(new_n684), .A4(new_n686), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n663), .B1(new_n710), .B2(new_n670), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n861), .A3(new_n758), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n752), .B(new_n741), .C1(new_n724), .C2(new_n723), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n731), .B2(new_n729), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n767), .A2(new_n772), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n774), .A2(new_n765), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n860), .A2(new_n861), .A3(new_n758), .A4(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n863), .A2(new_n865), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n755), .A2(new_n757), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT115), .A3(new_n754), .A4(new_n773), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n754), .A2(new_n773), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n876), .B2(new_n872), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n430), .A2(new_n599), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT114), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n640), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n695), .A2(new_n598), .A3(new_n640), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT114), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n883), .A3(new_n622), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n724), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n430), .A2(KEYINPUT113), .A3(new_n636), .A4(new_n640), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n622), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n607), .B1(new_n659), .B2(new_n353), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI211_X1 g704(.A(new_n598), .B(new_n646), .C1(new_n601), .C2(new_n664), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n714), .A2(new_n773), .A3(new_n891), .A4(new_n740), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n779), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n878), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n848), .B1(new_n871), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n863), .A2(new_n870), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n884), .A2(new_n893), .A3(new_n888), .A4(new_n889), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n877), .B2(new_n874), .ZN(new_n898));
  INV_X1    g712(.A(new_n864), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n732), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n775), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT53), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n900), .B2(new_n775), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n865), .A2(KEYINPUT118), .A3(new_n868), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n898), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n895), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n847), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT122), .Z(new_n915));
  OAI21_X1  g729(.A(new_n813), .B1(new_n913), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n189), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n243), .B1(new_n909), .B2(new_n895), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n542), .A2(new_n549), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n547), .A2(new_n544), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n550), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n918), .B1(new_n920), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n920), .B2(new_n926), .ZN(G51));
  NAND2_X1  g742(.A1(new_n909), .A2(new_n895), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT54), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(KEYINPUT123), .A3(new_n911), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n929), .A2(new_n932), .A3(KEYINPUT54), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n435), .B(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n473), .A2(new_n481), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n919), .A2(new_n784), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n917), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  AND3_X1   g755(.A1(new_n919), .A2(new_n410), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n410), .B1(new_n919), .B2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n917), .ZN(G60));
  AND2_X1   g758(.A1(new_n628), .A2(new_n629), .ZN(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT59), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n945), .A2(new_n931), .A3(new_n933), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n904), .B2(new_n911), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n918), .B1(new_n950), .B2(new_n945), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n909), .B2(new_n895), .ZN(new_n955));
  INV_X1    g769(.A(new_n240), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n657), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n918), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n957), .A2(KEYINPUT61), .A3(new_n918), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(G66));
  OAI21_X1  g777(.A(G953), .B1(new_n508), .B2(new_n602), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n865), .A2(new_n890), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(G953), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n921), .B1(G898), .B2(new_n189), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G69));
  XOR2_X1   g782(.A(new_n319), .B(new_n398), .Z(new_n969));
  OR2_X1    g783(.A1(new_n637), .A2(new_n879), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n970), .A2(new_n353), .A3(new_n699), .A4(new_n773), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n807), .B(new_n971), .C1(new_n798), .C2(new_n799), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n861), .A2(new_n758), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n705), .A2(new_n706), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(KEYINPUT62), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n976));
  AOI211_X1 g790(.A(G953), .B(new_n969), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n969), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n807), .B1(new_n798), .B2(new_n799), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n790), .A2(new_n554), .A3(new_n750), .A4(new_n772), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n973), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n868), .A2(new_n779), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n189), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(G900), .A2(G953), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n977), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(G227), .A2(G900), .ZN(new_n991));
  AND4_X1   g805(.A1(G953), .A2(new_n990), .A3(new_n991), .A4(new_n969), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n989), .A2(new_n992), .ZN(G72));
  XNOR2_X1  g807(.A(new_n329), .B(KEYINPUT127), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n975), .A2(new_n976), .A3(new_n965), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n674), .B(KEYINPUT63), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  AOI211_X1 g812(.A(new_n330), .B(new_n995), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n982), .A2(new_n965), .A3(new_n984), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n315), .B(new_n994), .C1(new_n1000), .C2(new_n998), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n331), .A2(new_n320), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n903), .A2(new_n997), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n918), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n999), .A2(new_n1001), .A3(new_n1004), .ZN(G57));
endmodule


