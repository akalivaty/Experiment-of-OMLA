//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND4_X1  g038(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n465), .B1(new_n459), .B2(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n458), .A2(new_n464), .B1(new_n468), .B2(G101), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n464), .A2(new_n458), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT65), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n471), .A2(new_n475), .ZN(G160));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n460), .A2(new_n462), .ZN(new_n479));
  OR2_X1    g054(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G2105), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n463), .A3(new_n481), .ZN(new_n485));
  OAI221_X1 g060(.A(new_n478), .B1(new_n482), .B2(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NOR2_X1   g062(.A1(new_n463), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n460), .A2(new_n462), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(KEYINPUT69), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n460), .A2(new_n462), .A3(new_n492), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n463), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n498), .B(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G651), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n503), .A2(new_n505), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G50), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n507), .B(KEYINPUT70), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n503), .A2(new_n505), .A3(new_n513), .A4(new_n515), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n510), .A2(new_n502), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n517), .ZN(G166));
  XNOR2_X1  g093(.A(KEYINPUT71), .B(G51), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n506), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(new_n509), .A3(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(KEYINPUT72), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(KEYINPUT7), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT7), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  NOR3_X1   g105(.A1(new_n524), .A2(new_n529), .A3(new_n530), .ZN(G168));
  NAND3_X1  g106(.A1(new_n513), .A2(new_n515), .A3(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n503), .A2(new_n505), .A3(G52), .A4(G543), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n521), .A2(new_n509), .A3(G90), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(G171));
  NAND3_X1  g114(.A1(new_n521), .A2(new_n509), .A3(G81), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n521), .A2(G43), .A3(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n513), .A2(new_n515), .A3(G56), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n502), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n548), .A2(new_n553), .ZN(G188));
  NAND4_X1  g129(.A1(new_n503), .A2(new_n505), .A3(G53), .A4(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT9), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n521), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n556), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n513), .A2(new_n515), .ZN(new_n563));
  INV_X1    g138(.A(G65), .ZN(new_n564));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(new_n512), .ZN(new_n566));
  AND4_X1   g141(.A1(new_n503), .A2(new_n505), .A3(new_n513), .A4(new_n515), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n566), .A2(G651), .B1(new_n567), .B2(G91), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n560), .A2(new_n562), .A3(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n535), .A2(new_n570), .A3(new_n536), .A4(new_n537), .ZN(new_n571));
  INV_X1    g146(.A(G90), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n536), .B1(new_n516), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n502), .B1(new_n532), .B2(new_n533), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT76), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G301));
  NOR2_X1   g151(.A1(new_n529), .A2(new_n530), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n577), .A2(new_n520), .A3(new_n522), .A4(new_n523), .ZN(G286));
  OR2_X1    g153(.A1(new_n508), .A2(new_n517), .ZN(G303));
  NAND2_X1  g154(.A1(new_n567), .A2(G87), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n506), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n567), .A2(G86), .B1(new_n506), .B2(G48), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n502), .B2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n567), .A2(G85), .B1(new_n506), .B2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n502), .B2(new_n588), .ZN(G290));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n516), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n521), .A2(new_n509), .A3(KEYINPUT10), .A4(G92), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n513), .A2(new_n515), .A3(G66), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n506), .B2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G301), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G284));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(new_n600), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n600), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n600), .B2(G168), .ZN(G280));
  NAND3_X1  g182(.A1(new_n521), .A2(G54), .A3(G543), .ZN(new_n608));
  INV_X1    g183(.A(new_n596), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(new_n509), .B2(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n608), .B1(new_n610), .B2(new_n502), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n592), .B2(new_n593), .ZN(new_n612));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G860), .ZN(G148));
  AND2_X1   g189(.A1(new_n543), .A2(new_n544), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n541), .B(new_n540), .C1(new_n615), .C2(new_n502), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n600), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n599), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n600), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n491), .A2(new_n468), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT13), .Z(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n623), .A2(KEYINPUT77), .A3(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n627), .B1(new_n482), .B2(new_n628), .C1(new_n629), .C2(new_n485), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  OAI21_X1  g206(.A(new_n623), .B1(KEYINPUT77), .B2(new_n624), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n624), .A2(KEYINPUT77), .ZN(new_n633));
  NAND4_X1  g208(.A1(new_n625), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(G2451), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT15), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2435), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n638), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT80), .A4(G14), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI21_X1  g239(.A(KEYINPUT17), .B1(new_n656), .B2(new_n657), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n658), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n663), .B(new_n664), .C1(new_n666), .C2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n685), .A2(KEYINPUT20), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(KEYINPUT20), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n679), .A2(new_n680), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n681), .A2(new_n684), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n686), .A2(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n683), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT84), .Z(new_n692));
  INV_X1    g267(.A(KEYINPUT85), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n693), .B1(new_n690), .B2(new_n692), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n695), .A2(G1991), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G1991), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n690), .A2(new_n692), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT85), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n698), .B1(new_n700), .B2(new_n694), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n677), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(G1991), .B1(new_n695), .B2(new_n696), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n698), .A3(new_n694), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(G1996), .A3(new_n706), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n704), .B1(new_n702), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n676), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n702), .A2(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(new_n703), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n702), .A2(new_n704), .A3(new_n707), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n712), .A2(new_n675), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1971), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(G6), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n521), .A2(G543), .ZN(new_n723));
  INV_X1    g298(.A(G48), .ZN(new_n724));
  INV_X1    g299(.A(G86), .ZN(new_n725));
  OAI22_X1  g300(.A1(new_n723), .A2(new_n724), .B1(new_n516), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n509), .A2(G61), .ZN(new_n727));
  NAND2_X1  g302(.A1(G73), .A2(G543), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n502), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n722), .B1(new_n730), .B2(new_n718), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT32), .B(G1981), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT87), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G23), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT88), .Z(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G288), .B2(new_n718), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT33), .B(G1976), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n721), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT34), .ZN(new_n742));
  INV_X1    g317(.A(new_n482), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n743), .A2(KEYINPUT86), .A3(G119), .ZN(new_n744));
  INV_X1    g319(.A(new_n485), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G131), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT86), .ZN(new_n747));
  INV_X1    g322(.A(G119), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n482), .B2(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(G95), .A2(G2105), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n750), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n744), .A2(new_n746), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  MUX2_X1   g327(.A(G25), .B(new_n752), .S(G29), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT35), .B(G1991), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n753), .B(new_n754), .Z(new_n755));
  MUX2_X1   g330(.A(G24), .B(G290), .S(G16), .Z(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(G1986), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n742), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n716), .B(new_n717), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G29), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2090), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  AND2_X1   g341(.A1(new_n761), .A2(G26), .ZN(new_n767));
  OR2_X1    g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT91), .Z(new_n770));
  INV_X1    g345(.A(G128), .ZN(new_n771));
  INV_X1    g346(.A(G140), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n770), .B1(new_n482), .B2(new_n771), .C1(new_n772), .C2(new_n485), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(G29), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n767), .B(new_n774), .S(KEYINPUT28), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT26), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  AOI22_X1  g355(.A1(G105), .A2(new_n468), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G129), .ZN(new_n782));
  INV_X1    g357(.A(G141), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n781), .B1(new_n482), .B2(new_n782), .C1(new_n783), .C2(new_n485), .ZN(new_n784));
  MUX2_X1   g359(.A(G32), .B(new_n784), .S(G29), .Z(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n630), .A2(new_n761), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G171), .B2(G16), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  INV_X1    g366(.A(G28), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT30), .ZN(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n792), .B2(KEYINPUT30), .ZN(new_n794));
  OR2_X1    g369(.A1(KEYINPUT31), .A2(G11), .ZN(new_n795));
  NAND2_X1  g370(.A1(KEYINPUT31), .A2(G11), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n790), .A2(G1961), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n788), .A2(new_n791), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n718), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n612), .B2(new_n718), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1348), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n787), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n776), .B(new_n803), .C1(G2090), .C2(new_n764), .ZN(new_n804));
  NAND2_X1  g379(.A1(G168), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G16), .B2(G21), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G29), .A2(G33), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT92), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n491), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n814));
  INV_X1    g389(.A(G139), .ZN(new_n815));
  OAI221_X1 g390(.A(new_n813), .B1(new_n814), .B2(new_n463), .C1(new_n485), .C2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(new_n761), .ZN(new_n817));
  INV_X1    g392(.A(G2072), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(G164), .A2(G29), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G27), .B2(G29), .ZN(new_n821));
  INV_X1    g396(.A(G2078), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n808), .B(new_n823), .C1(new_n822), .C2(new_n821), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n718), .A2(G20), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n825), .B(new_n826), .C1(G299), .C2(G16), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  INV_X1    g403(.A(G1956), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G34), .ZN(new_n831));
  AOI21_X1  g406(.A(G29), .B1(new_n831), .B2(KEYINPUT24), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n832), .A2(KEYINPUT94), .B1(KEYINPUT24), .B2(new_n831), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(KEYINPUT94), .B2(new_n832), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G160), .B2(G29), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G2084), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT95), .ZN(new_n839));
  NOR2_X1   g414(.A1(G16), .A2(G19), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n546), .B2(G16), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1341), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n836), .A2(new_n837), .B1(new_n817), .B2(new_n818), .ZN(new_n843));
  AOI211_X1 g418(.A(new_n842), .B(new_n843), .C1(new_n807), .C2(new_n806), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n824), .A2(new_n830), .A3(new_n839), .A4(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n766), .A2(new_n804), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n758), .A2(new_n759), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n847), .A2(KEYINPUT89), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT36), .B1(new_n758), .B2(new_n716), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n760), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(G150));
  INV_X1    g425(.A(G150), .ZN(G311));
  XNOR2_X1  g426(.A(KEYINPUT98), .B(G860), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n513), .A2(new_n515), .A3(G67), .ZN(new_n853));
  NAND2_X1  g428(.A1(G80), .A2(G543), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G651), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n503), .A2(new_n505), .A3(G55), .A4(G543), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n521), .A2(new_n509), .A3(G93), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n856), .A2(KEYINPUT97), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n857), .B1(new_n516), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n502), .B1(new_n853), .B2(new_n854), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n864), .A3(new_n546), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n616), .A2(new_n866), .A3(new_n860), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n612), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n852), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n873), .B1(new_n872), .B2(new_n871), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(new_n852), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT37), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(G145));
  XNOR2_X1  g452(.A(new_n752), .B(new_n816), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n743), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n745), .A2(G142), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n463), .A2(KEYINPUT99), .A3(G118), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT99), .B1(new_n463), .B2(G118), .ZN(new_n882));
  OR2_X1    g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(G2104), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n879), .B(new_n880), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G164), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n878), .A2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n486), .B(new_n630), .Z(new_n890));
  XNOR2_X1  g465(.A(new_n773), .B(G160), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n892), .B(new_n893), .C1(new_n887), .C2(new_n888), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n622), .B(KEYINPUT100), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n784), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n895), .A2(new_n899), .A3(new_n896), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g480(.A1(new_n866), .A2(new_n600), .ZN(new_n906));
  NAND2_X1  g481(.A1(G303), .A2(new_n730), .ZN(new_n907));
  NAND2_X1  g482(.A1(G166), .A2(G305), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G290), .B(G288), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n910), .A3(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(KEYINPUT102), .A2(KEYINPUT42), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G299), .A2(new_n612), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n561), .B1(new_n556), .B2(new_n558), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n521), .A2(new_n509), .A3(G91), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n565), .A2(new_n512), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n509), .B2(G65), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n502), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n599), .A3(new_n562), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n919), .A2(new_n926), .A3(KEYINPUT101), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n925), .A2(new_n599), .A3(new_n929), .A4(new_n562), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n919), .A2(new_n926), .A3(KEYINPUT41), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n868), .B(new_n618), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n919), .A2(new_n926), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n935), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n918), .B(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n906), .B1(new_n938), .B2(new_n600), .ZN(G295));
  XNOR2_X1  g514(.A(G295), .B(KEYINPUT103), .ZN(G331));
  AOI21_X1  g515(.A(G286), .B1(new_n575), .B2(new_n571), .ZN(new_n941));
  INV_X1    g516(.A(new_n524), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n538), .B1(new_n942), .B2(new_n577), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n867), .B(new_n865), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(G301), .A2(G168), .ZN(new_n945));
  NAND2_X1  g520(.A1(G171), .A2(G286), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n868), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n927), .A2(KEYINPUT41), .A3(new_n930), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(KEYINPUT41), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n946), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n865), .A2(new_n867), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n952), .A2(new_n956), .B1(new_n948), .B2(new_n949), .ZN(new_n957));
  INV_X1    g532(.A(new_n936), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n914), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n913), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT43), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n955), .B1(new_n948), .B2(new_n951), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n965), .B1(new_n966), .B2(new_n933), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n931), .A2(new_n932), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n944), .B2(new_n947), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n968), .B(KEYINPUT105), .C1(new_n969), .C2(new_n955), .ZN(new_n970));
  INV_X1    g545(.A(new_n948), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n936), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n914), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n969), .B2(new_n955), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n976), .A2(new_n965), .B1(new_n936), .B2(new_n971), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(KEYINPUT107), .A3(new_n914), .A4(new_n970), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n964), .A2(new_n975), .A3(new_n902), .A4(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n967), .A2(new_n970), .A3(new_n972), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n963), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n975), .A2(new_n983), .A3(new_n978), .A4(new_n902), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  AOI21_X1  g560(.A(G37), .B1(new_n973), .B2(new_n974), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(KEYINPUT108), .A3(new_n964), .A4(new_n978), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n959), .B2(new_n963), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n986), .A2(new_n978), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(G397));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n494), .A2(new_n495), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n494), .A2(new_n495), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n998), .A2(new_n999), .B1(new_n488), .B2(new_n489), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT4), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n498), .B(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n997), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n475), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(G40), .A3(new_n469), .A4(new_n470), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n773), .B(G2067), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n784), .B(new_n677), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n752), .A2(new_n754), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n752), .A2(new_n754), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(G290), .B(G1986), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1009), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1008), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n497), .B2(new_n499), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT45), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1024), .B2(G2078), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1008), .B1(new_n1022), .B2(new_n1004), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1003), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1026), .A2(new_n1028), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1022), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n471), .A2(new_n1033), .A3(new_n475), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1025), .A2(new_n1029), .A3(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1038), .A2(new_n602), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1034), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT50), .B(G1384), .C1(new_n497), .C2(new_n499), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n1041), .A2(G2084), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1966), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(G168), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT51), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1044), .B2(new_n1043), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1034), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1022), .A2(KEYINPUT45), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n807), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1008), .B1(new_n1003), .B2(KEYINPUT50), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n837), .A3(new_n1032), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1046), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1052), .B1(new_n1058), .B2(new_n1049), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1051), .B1(new_n1059), .B2(KEYINPUT51), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1040), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(new_n1052), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT62), .B1(new_n1066), .B2(new_n1051), .ZN(new_n1067));
  INV_X1    g642(.A(G288), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G1976), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT112), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1034), .A2(new_n1022), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(G8), .ZN(new_n1073));
  AOI211_X1 g648(.A(KEYINPUT111), .B(new_n1046), .C1(new_n1034), .C2(new_n1022), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(G8), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT111), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1071), .A3(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n1070), .ZN(new_n1082));
  OR3_X1    g657(.A1(new_n1068), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G303), .A2(G8), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1971), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT110), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1088), .A2(new_n1089), .B1(G2090), .B2(new_n1035), .ZN(new_n1090));
  INV_X1    g665(.A(G1971), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1034), .B1(new_n1022), .B2(new_n1004), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1003), .A2(new_n1027), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(KEYINPUT110), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1087), .B(G8), .C1(new_n1090), .C2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1085), .B(KEYINPUT55), .ZN(new_n1097));
  INV_X1    g672(.A(G2090), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1088), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1100), .B2(new_n1046), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT114), .B(G1981), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(G305), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1102), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n730), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(G305), .A2(KEYINPUT116), .A3(G1981), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  INV_X1    g684(.A(G1981), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n730), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1112), .A3(KEYINPUT49), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1107), .A2(new_n1112), .A3(new_n1115), .A4(KEYINPUT49), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT49), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1084), .A2(new_n1096), .A3(new_n1101), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1062), .A2(new_n1063), .A3(new_n1067), .A4(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1084), .A2(new_n1121), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1094), .A2(KEYINPUT110), .B1(new_n1099), .B2(new_n1098), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1046), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1128), .A2(new_n1087), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1058), .A2(G168), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1125), .A2(new_n1129), .A3(new_n1096), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT57), .B(new_n924), .C1(KEYINPUT119), .C2(new_n559), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n559), .A2(KEYINPUT119), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1136), .A2(new_n1137), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1035), .A2(new_n829), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1021), .A2(new_n1023), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(G1348), .B1(new_n1056), .B2(new_n1032), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1072), .A2(G2067), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1145), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1139), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n612), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1143), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(new_n1153), .A3(new_n1148), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n599), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1153), .B(new_n612), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1150), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1150), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1160), .B2(new_n1142), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1072), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1024), .B2(G1996), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n546), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(KEYINPUT59), .A3(new_n546), .ZN(new_n1168));
  AND4_X1   g743(.A1(new_n1158), .A2(new_n1161), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1152), .B1(new_n1157), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1037), .A2(KEYINPUT122), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1021), .A2(KEYINPUT53), .A3(new_n822), .A4(new_n1023), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1035), .A2(new_n1173), .A3(new_n1036), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1171), .A2(new_n1025), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1174), .A2(new_n1172), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1178), .A2(KEYINPUT123), .A3(new_n1025), .A4(new_n1171), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1179), .A3(G171), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1038), .A2(new_n602), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1060), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1175), .A2(new_n602), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1182), .B1(new_n1186), .B2(new_n1039), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1184), .A2(new_n1123), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1124), .B(new_n1135), .C1(new_n1170), .C2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1123), .A2(new_n1067), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1051), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1191), .A2(new_n1061), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1039), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT124), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(G288), .A2(G1976), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1196), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1107), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1081), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1084), .A2(new_n1128), .A3(new_n1087), .A4(new_n1121), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT118), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT118), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1195), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1019), .B1(new_n1189), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1009), .B1(new_n1010), .B2(new_n784), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1009), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT46), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1009), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(G1996), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1206), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(new_n1211), .B(KEYINPUT47), .Z(new_n1212));
  OR2_X1    g787(.A1(new_n1015), .A2(KEYINPUT125), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1015), .A2(KEYINPUT125), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1213), .A2(new_n1011), .A3(new_n1012), .A4(new_n1214), .ZN(new_n1215));
  OR2_X1    g790(.A1(new_n773), .A2(G2067), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1209), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1209), .A2(G1986), .A3(G290), .ZN(new_n1218));
  XOR2_X1   g793(.A(new_n1218), .B(KEYINPUT126), .Z(new_n1219));
  INV_X1    g794(.A(KEYINPUT48), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1221), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1223));
  AOI211_X1 g798(.A(new_n1212), .B(new_n1217), .C1(new_n1222), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1205), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g800(.A1(new_n710), .A2(new_n714), .ZN(new_n1227));
  NAND3_X1  g801(.A1(new_n672), .A2(G319), .A3(new_n673), .ZN(new_n1228));
  XNOR2_X1  g802(.A(new_n1228), .B(KEYINPUT127), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1229), .B1(new_n653), .B2(new_n654), .ZN(new_n1230));
  AND2_X1   g804(.A1(new_n1230), .A2(new_n904), .ZN(new_n1231));
  AND3_X1   g805(.A1(new_n1227), .A2(new_n988), .A3(new_n1231), .ZN(G308));
  NAND4_X1  g806(.A1(new_n988), .A2(new_n1231), .A3(new_n714), .A4(new_n710), .ZN(G225));
endmodule


