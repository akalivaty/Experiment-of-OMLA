//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1253, new_n1254, new_n1255, new_n1256;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n463), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n463), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n489), .A2(new_n490), .A3(G138), .A4(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n463), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n496), .A2(new_n500), .B1(new_n480), .B2(G126), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n492), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT71), .B(G88), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(G62), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT72), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n518), .A2(new_n519), .A3(new_n508), .A4(new_n507), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(G166));
  NOR2_X1   g096(.A1(new_n511), .A2(new_n512), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n504), .A2(KEYINPUT73), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n530));
  AND3_X1   g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n505), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n512), .A2(new_n511), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n532), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n529), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n524), .A2(new_n525), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  AOI22_X1  g122(.A1(G52), .A2(new_n533), .B1(new_n538), .B2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n505), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n552), .B1(new_n537), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n544), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n554), .B1(new_n557), .B2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n533), .A2(new_n564), .A3(G53), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n551), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n522), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(G651), .A2(new_n571), .B1(new_n538), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G166), .ZN(G303));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n551), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n505), .A2(KEYINPUT76), .A3(G49), .A4(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n538), .A2(G87), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n524), .B2(new_n525), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n510), .C2(new_n581), .ZN(G288));
  OAI21_X1  g157(.A(G61), .B1(new_n511), .B2(new_n512), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n510), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT77), .B1(new_n537), .B2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n504), .A2(new_n505), .A3(new_n588), .A4(G86), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n533), .A2(G48), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n551), .A2(new_n598), .B1(new_n537), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G60), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n544), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n600), .B1(new_n603), .B2(G651), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n538), .A2(G92), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n522), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(new_n533), .B2(G54), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n606), .B1(new_n615), .B2(G868), .ZN(G321));
  AND2_X1   g192(.A1(new_n568), .A2(new_n572), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n618), .B2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  MUX2_X1   g195(.A(KEYINPUT79), .B(new_n619), .S(new_n620), .Z(G297));
  MUX2_X1   g196(.A(KEYINPUT79), .B(new_n619), .S(new_n620), .Z(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n623), .B2(G860), .ZN(G148));
  NOR2_X1   g199(.A1(new_n614), .A2(G559), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  OR3_X1    g201(.A1(new_n625), .A2(KEYINPUT80), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n625), .B2(new_n626), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n627), .B(new_n628), .C1(G868), .C2(new_n558), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g205(.A1(new_n475), .A2(G2105), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n489), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n478), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n480), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n463), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT81), .Z(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n635), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g221(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  XOR2_X1   g223(.A(G2443), .B(G2446), .Z(new_n649));
  XOR2_X1   g224(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  INV_X1    g227(.A(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2430), .Z(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2451), .B(G2454), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n651), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(new_n650), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1341), .B(G1348), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(G14), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT87), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n666), .A2(new_n670), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n675), .B1(new_n676), .B2(new_n671), .ZN(new_n677));
  AOI211_X1 g252(.A(KEYINPUT87), .B(new_n672), .C1(new_n666), .C2(new_n670), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G401));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT17), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n681), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G2100), .ZN(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n684), .B2(KEYINPUT18), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G2096), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1956), .B(G2474), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n696), .B1(new_n701), .B2(KEYINPUT89), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(KEYINPUT89), .B2(new_n701), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT20), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n696), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n705), .B(new_n696), .S(new_n706), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT90), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n704), .A2(new_n710), .A3(new_n707), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n715), .B1(new_n712), .B2(new_n716), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n694), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n719), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n721), .A2(new_n693), .A3(new_n717), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(G229));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G32), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n631), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n480), .A2(G129), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n478), .A2(G139), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n489), .A2(G127), .ZN(new_n738));
  NAND2_X1  g313(.A1(G115), .A2(G2104), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n463), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(new_n724), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n724), .B2(G33), .ZN(new_n743));
  INV_X1    g318(.A(G2072), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n733), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G160), .B2(new_n724), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n745), .B1(new_n744), .B2(new_n743), .C1(G2084), .C2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G16), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G20), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT23), .Z(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G299), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n751), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n615), .B2(G16), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NOR2_X1   g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G28), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n724), .B1(new_n766), .B2(G28), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n640), .A2(new_n724), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n765), .B1(new_n767), .B2(new_n768), .C1(new_n769), .C2(KEYINPUT96), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(KEYINPUT96), .B2(new_n769), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n731), .A2(new_n732), .B1(new_n750), .B2(G2084), .ZN(new_n772));
  AND3_X1   g347(.A1(new_n762), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n724), .A2(G26), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT28), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n478), .A2(G140), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT92), .ZN(new_n777));
  OAI21_X1  g352(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n778));
  INV_X1    g353(.A(G116), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(G2105), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n489), .A2(G2105), .ZN(new_n781));
  INV_X1    g356(.A(G128), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT93), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n480), .A2(new_n784), .A3(G128), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n775), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n752), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n558), .B2(new_n752), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NAND4_X1  g367(.A1(new_n758), .A2(new_n773), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n752), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n752), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT94), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G1966), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT95), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n724), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n724), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n752), .A2(G5), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G171), .B2(new_n752), .ZN(new_n804));
  INV_X1    g379(.A(G1961), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n724), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n724), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT29), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n802), .B(new_n806), .C1(new_n809), .C2(G2090), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(G2090), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n796), .B2(G1966), .ZN(new_n812));
  NOR4_X1   g387(.A1(new_n793), .A2(new_n798), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n596), .A2(G16), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G6), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n752), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n752), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1971), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n752), .A2(G23), .ZN(new_n825));
  INV_X1    g400(.A(G288), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n752), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT33), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1976), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n752), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n752), .B2(G24), .ZN(new_n832));
  INV_X1    g407(.A(G1986), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n724), .A2(G25), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n478), .A2(G131), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n480), .A2(G119), .ZN(new_n838));
  OR2_X1    g413(.A1(G95), .A2(G2105), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n839), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n836), .B1(new_n842), .B2(new_n724), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT35), .B(G1991), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n843), .B(new_n845), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n834), .A2(new_n835), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n830), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n824), .B1(new_n823), .B2(new_n829), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT36), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n851), .A2(new_n830), .A3(new_n852), .A4(new_n847), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n814), .B1(new_n850), .B2(new_n853), .ZN(G311));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n813), .ZN(G150));
  NAND3_X1  g431(.A1(new_n524), .A2(new_n525), .A3(G67), .ZN(new_n857));
  NAND2_X1  g432(.A1(G80), .A2(G543), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n510), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI22_X1  g436(.A1(new_n551), .A2(new_n860), .B1(new_n537), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G860), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT37), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n615), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n857), .A2(new_n858), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G651), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT97), .ZN(new_n871));
  INV_X1    g446(.A(new_n862), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT97), .B1(new_n859), .B2(new_n862), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n873), .A2(new_n558), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n558), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n868), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n864), .B1(new_n879), .B2(KEYINPUT39), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n866), .B1(new_n880), .B2(new_n881), .ZN(G145));
  XOR2_X1   g457(.A(new_n502), .B(KEYINPUT98), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n777), .A2(new_n885), .A3(new_n786), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n777), .B2(new_n786), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n887), .A2(new_n888), .A3(new_n741), .ZN(new_n889));
  INV_X1    g464(.A(new_n741), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n787), .A2(new_n730), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(new_n886), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n884), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n478), .A2(G142), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n480), .A2(G130), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n463), .A2(G118), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n633), .B(new_n898), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n841), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n741), .B1(new_n887), .B2(new_n888), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n891), .A2(new_n890), .A3(new_n886), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n883), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n893), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT99), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n893), .A2(new_n900), .A3(new_n906), .A4(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n899), .B(new_n842), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n901), .A2(new_n883), .A3(new_n902), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n883), .B1(new_n901), .B2(new_n902), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n640), .B(G160), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n485), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT100), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g493(.A(KEYINPUT100), .B(new_n909), .C1(new_n910), .C2(new_n911), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n908), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g500(.A1(G290), .A2(G303), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n826), .B1(new_n594), .B2(new_n595), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n604), .A2(G166), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(G288), .A3(new_n593), .ZN(new_n930));
  AND4_X1   g505(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n927), .A2(new_n930), .B1(new_n926), .B2(new_n928), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  INV_X1    g511(.A(new_n558), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n859), .A2(KEYINPUT97), .A3(new_n862), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n873), .A2(new_n558), .A3(new_n874), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(new_n625), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n614), .A2(G299), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n618), .A2(new_n609), .A3(new_n613), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n936), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n942), .A2(new_n625), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n942), .A2(new_n625), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n936), .B(new_n947), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT41), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n614), .A2(G299), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n618), .B1(new_n609), .B2(new_n613), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n944), .A2(KEYINPUT41), .A3(new_n945), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n943), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n934), .B(new_n935), .C1(new_n948), .C2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n935), .B1(new_n959), .B2(new_n948), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n959), .A2(new_n948), .A3(new_n935), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n931), .A2(new_n932), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G868), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(G868), .B2(new_n863), .ZN(G295));
  OAI21_X1  g543(.A(new_n967), .B1(G868), .B2(new_n863), .ZN(G331));
  INV_X1    g544(.A(G37), .ZN(new_n970));
  AND4_X1   g545(.A1(new_n529), .A2(new_n547), .A3(new_n540), .A4(new_n548), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n529), .A2(new_n540), .B1(new_n547), .B2(new_n548), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n942), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G286), .A2(G301), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n529), .A2(new_n547), .A3(new_n540), .A4(new_n548), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n941), .A3(new_n940), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n957), .B1(new_n975), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(KEYINPUT104), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n946), .B1(new_n877), .B2(new_n978), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n942), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n986), .A3(new_n963), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n974), .A2(new_n979), .A3(new_n947), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n982), .A2(new_n979), .A3(new_n985), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n957), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n970), .B(new_n987), .C1(new_n990), .C2(new_n963), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT105), .B1(new_n991), .B2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n987), .A2(new_n970), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n989), .A2(new_n957), .ZN(new_n995));
  INV_X1    g570(.A(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n933), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT105), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n994), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n963), .B1(new_n981), .B2(new_n986), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT43), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n992), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n993), .A2(new_n1002), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n991), .A2(new_n1000), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1006), .A2(new_n1010), .ZN(G397));
  AOI21_X1  g586(.A(G1384), .B1(new_n492), .B2(new_n501), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1013));
  INV_X1    g588(.A(G125), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n476), .B2(new_n477), .ZN(new_n1015));
  INV_X1    g590(.A(new_n467), .ZN(new_n1016));
  OAI21_X1  g591(.A(G2105), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n470), .B1(new_n478), .B2(G137), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT106), .B(G40), .Z(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(G160), .A2(KEYINPUT107), .A3(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1013), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(G1996), .A3(new_n730), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT108), .ZN(new_n1028));
  INV_X1    g603(.A(G2067), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n787), .B(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(G1996), .B2(new_n730), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1028), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n842), .A2(new_n844), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n841), .A2(new_n845), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1026), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n604), .B(new_n833), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1026), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n591), .B1(new_n586), .B2(new_n537), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1039), .B2(new_n585), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT115), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1981), .B1(new_n533), .B2(G48), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n590), .A2(KEYINPUT114), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n590), .B2(new_n1043), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1040), .B(new_n1042), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n587), .A2(new_n589), .ZN(new_n1050));
  INV_X1    g625(.A(new_n585), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1043), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n590), .A2(KEYINPUT114), .A3(new_n1043), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1042), .B1(new_n1056), .B2(new_n1040), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT116), .B1(new_n1049), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1040), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1059), .A2(KEYINPUT115), .A3(new_n1041), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1048), .A4(new_n1046), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1384), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n502), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1024), .A3(new_n1068), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT109), .B(G1971), .Z(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1072));
  AOI22_X1  g647(.A1(new_n1023), .A2(new_n1022), .B1(new_n1012), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1065), .A2(KEYINPUT50), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1071), .B1(G2090), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n516), .A2(new_n520), .A3(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n516), .A2(new_n520), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(KEYINPUT111), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1076), .A2(G8), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n581), .A2(new_n510), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(G1976), .A3(new_n579), .A4(new_n580), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1087), .B1(new_n1048), .B2(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT112), .B(G1976), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(G288), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1048), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT113), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1048), .A2(new_n1095), .A3(new_n1092), .A4(new_n1089), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1063), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1023), .A2(new_n1022), .B1(new_n1012), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G2090), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1072), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1065), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1071), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1047), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1071), .A2(KEYINPUT117), .A3(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1081), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1098), .A2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(G301), .B(KEYINPUT54), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n805), .B2(new_n1075), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1069), .B2(G2078), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1018), .A2(KEYINPUT53), .A3(G40), .A4(new_n801), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(KEYINPUT125), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n463), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(KEYINPUT125), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT126), .Z(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT107), .B1(G160), .B2(new_n1019), .ZN(new_n1124));
  AND4_X1   g699(.A1(KEYINPUT107), .A2(new_n1017), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1066), .B(G1384), .C1(new_n492), .C2(new_n501), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1126), .A2(new_n1013), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT53), .A3(new_n801), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1075), .A2(new_n805), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(new_n1114), .A3(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1115), .A2(new_n1123), .B1(new_n1111), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  INV_X1    g708(.A(G2084), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1012), .A2(new_n1072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1074), .A2(new_n1024), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1966), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1069), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1073), .A2(KEYINPUT118), .A3(new_n1134), .A4(new_n1074), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(G168), .A4(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1142), .A2(G8), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G286), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1133), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1142), .A2(G8), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(KEYINPUT51), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1110), .B(new_n1132), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n1151));
  INV_X1    g726(.A(G1996), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1067), .A2(new_n1024), .A3(new_n1152), .A4(new_n1068), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1012), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT58), .B(G1341), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1156), .A3(KEYINPUT122), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1151), .B1(new_n1161), .B2(new_n558), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1153), .A2(new_n1156), .A3(KEYINPUT122), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT122), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1151), .B(new_n558), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT56), .B(G2072), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1067), .A2(new_n1024), .A3(new_n1068), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(G1956), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1168), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1012), .A2(new_n1099), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1103), .A2(new_n1024), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n756), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1176), .A2(KEYINPUT121), .A3(new_n1170), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1178));
  XNOR2_X1  g753(.A(G299), .B(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1173), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1128), .A2(new_n1169), .B1(new_n1175), .B2(new_n756), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1179), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1183), .B1(new_n1176), .B2(new_n1170), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1171), .A2(new_n1172), .A3(new_n1179), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1150), .B1(new_n1167), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n558), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(KEYINPUT59), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1165), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(KEYINPUT124), .A3(new_n1185), .A4(new_n1189), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1154), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1075), .A2(new_n761), .B1(new_n1196), .B2(new_n1029), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1197), .A2(KEYINPUT60), .A3(new_n614), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n614), .B1(new_n1197), .B2(KEYINPUT60), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n1198), .A2(new_n1199), .B1(KEYINPUT60), .B2(new_n1197), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1191), .A2(new_n1195), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1180), .ZN(new_n1202));
  NOR3_X1   g777(.A1(new_n1188), .A2(new_n614), .A3(new_n1197), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1149), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1063), .A2(new_n1086), .A3(new_n1097), .ZN(new_n1206));
  NOR2_X1   g781(.A1(G286), .A2(new_n1047), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1144), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT119), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n1207), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1076), .A2(G8), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1082), .ZN(new_n1214));
  NAND4_X1  g789(.A1(new_n1206), .A2(KEYINPUT63), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  AND3_X1   g790(.A1(new_n1144), .A2(KEYINPUT119), .A3(new_n1207), .ZN(new_n1216));
  AOI21_X1  g791(.A(KEYINPUT119), .B1(new_n1144), .B2(new_n1207), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NOR3_X1   g793(.A1(new_n1218), .A2(new_n1098), .A3(new_n1109), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1215), .B1(new_n1219), .B2(KEYINPUT63), .ZN(new_n1220));
  OAI21_X1  g795(.A(KEYINPUT62), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1221));
  INV_X1    g796(.A(new_n1145), .ZN(new_n1222));
  OAI21_X1  g797(.A(KEYINPUT51), .B1(new_n1222), .B2(new_n1147), .ZN(new_n1223));
  INV_X1    g798(.A(new_n1148), .ZN(new_n1224));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1223), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1131), .A2(G171), .ZN(new_n1227));
  NOR3_X1   g802(.A1(new_n1098), .A2(new_n1109), .A3(new_n1227), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1221), .A2(new_n1226), .A3(new_n1228), .ZN(new_n1229));
  AOI211_X1 g804(.A(G1976), .B(G288), .C1(new_n1058), .C2(new_n1062), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1056), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1048), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1063), .A2(new_n1097), .ZN(new_n1233));
  OR2_X1    g808(.A1(new_n1233), .A2(new_n1086), .ZN(new_n1234));
  AND2_X1   g809(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1220), .A2(new_n1229), .A3(new_n1235), .ZN(new_n1236));
  OAI21_X1  g811(.A(new_n1038), .B1(new_n1205), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1025), .B1(new_n1030), .B2(new_n885), .ZN(new_n1238));
  OAI21_X1  g813(.A(KEYINPUT46), .B1(new_n1025), .B2(G1996), .ZN(new_n1239));
  OR3_X1    g814(.A1(new_n1025), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1240));
  AOI21_X1  g815(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  XNOR2_X1  g816(.A(new_n1241), .B(KEYINPUT47), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n777), .A2(new_n786), .A3(new_n1029), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1025), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1036), .ZN(new_n1246));
  NOR3_X1   g821(.A1(new_n1025), .A2(G1986), .A3(G290), .ZN(new_n1247));
  XNOR2_X1  g822(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1248));
  XNOR2_X1  g823(.A(new_n1247), .B(new_n1248), .ZN(new_n1249));
  AOI211_X1 g824(.A(new_n1242), .B(new_n1245), .C1(new_n1246), .C2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1237), .A2(new_n1250), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g826(.A1(G227), .A2(new_n461), .ZN(new_n1253));
  NAND4_X1  g827(.A1(new_n679), .A2(new_n722), .A3(new_n720), .A4(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g828(.A(new_n920), .B(new_n921), .ZN(new_n1255));
  AOI21_X1  g829(.A(new_n1254), .B1(new_n1255), .B2(new_n916), .ZN(new_n1256));
  AND2_X1   g830(.A1(new_n1256), .A2(new_n1004), .ZN(G308));
  NAND2_X1  g831(.A1(new_n1256), .A2(new_n1004), .ZN(G225));
endmodule


