

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(n532), .A2(n627), .ZN(n642) );
  AND2_X1 U556 ( .A1(G125), .A2(n870), .ZN(n520) );
  XNOR2_X1 U557 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n727) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n766), .ZN(n746) );
  INV_X1 U559 ( .A(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U560 ( .A1(n770), .A2(n685), .ZN(n733) );
  NOR2_X1 U561 ( .A1(G651), .A2(n627), .ZN(n636) );
  NOR2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n521) );
  NOR2_X1 U563 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U564 ( .A1(n526), .A2(n520), .ZN(n527) );
  AND2_X1 U565 ( .A1(n528), .A2(n527), .ZN(G160) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n521), .Z(n865) );
  NAND2_X1 U567 ( .A1(G137), .A2(n865), .ZN(n528) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n868) );
  NAND2_X1 U569 ( .A1(n868), .A2(G113), .ZN(n524) );
  INV_X1 U570 ( .A(G2105), .ZN(n525) );
  AND2_X1 U571 ( .A1(n525), .A2(G2104), .ZN(n864) );
  NAND2_X1 U572 ( .A1(G101), .A2(n864), .ZN(n522) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n526) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n525), .ZN(n870) );
  AND2_X1 U576 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U577 ( .A(G132), .ZN(G219) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n638) );
  NAND2_X1 U579 ( .A1(G88), .A2(n638), .ZN(n531) );
  INV_X1 U580 ( .A(G651), .ZN(n532) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n529) );
  XNOR2_X1 U582 ( .A(KEYINPUT64), .B(n529), .ZN(n627) );
  NAND2_X1 U583 ( .A1(G75), .A2(n642), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n537) );
  NAND2_X1 U585 ( .A1(G50), .A2(n636), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n533), .Z(n639) );
  NAND2_X1 U588 ( .A1(G62), .A2(n639), .ZN(n534) );
  NAND2_X1 U589 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n537), .A2(n536), .ZN(G166) );
  NAND2_X1 U591 ( .A1(n639), .A2(G64), .ZN(n538) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n538), .Z(n540) );
  NAND2_X1 U593 ( .A1(n636), .A2(G52), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U595 ( .A(KEYINPUT66), .B(n541), .ZN(n547) );
  NAND2_X1 U596 ( .A1(G90), .A2(n638), .ZN(n543) );
  NAND2_X1 U597 ( .A1(G77), .A2(n642), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(n544), .ZN(n545) );
  XNOR2_X1 U600 ( .A(KEYINPUT9), .B(n545), .ZN(n546) );
  NOR2_X1 U601 ( .A1(n547), .A2(n546), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G51), .A2(n636), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G63), .A2(n639), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U605 ( .A(KEYINPUT6), .B(n550), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n642), .A2(G76), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n551), .B(KEYINPUT76), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n638), .A2(G89), .ZN(n552) );
  XNOR2_X1 U609 ( .A(KEYINPUT4), .B(n552), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U611 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT7), .B(n558), .Z(n559) );
  XOR2_X1 U613 ( .A(KEYINPUT77), .B(n559), .Z(G168) );
  XOR2_X1 U614 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n560) );
  XNOR2_X1 U616 ( .A(n560), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U617 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n562) );
  INV_X1 U618 ( .A(G223), .ZN(n821) );
  NAND2_X1 U619 ( .A1(G567), .A2(n821), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n562), .B(n561), .ZN(G234) );
  INV_X1 U621 ( .A(G860), .ZN(n614) );
  INV_X1 U622 ( .A(KEYINPUT74), .ZN(n574) );
  NAND2_X1 U623 ( .A1(n638), .A2(G81), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT12), .B(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n642), .A2(G68), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT73), .B(n564), .Z(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G43), .A2(n636), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n639), .A2(G56), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U634 ( .A(n574), .B(n573), .ZN(n932) );
  OR2_X1 U635 ( .A1(n614), .A2(n932), .ZN(G153) );
  INV_X1 U636 ( .A(G171), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U638 ( .A1(n639), .A2(G66), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G79), .A2(n642), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G54), .A2(n636), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G92), .A2(n638), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT75), .B(n577), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n582), .Z(n917) );
  INV_X1 U647 ( .A(G868), .ZN(n593) );
  NAND2_X1 U648 ( .A1(n917), .A2(n593), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G78), .A2(n642), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(KEYINPUT68), .ZN(n592) );
  NAND2_X1 U652 ( .A1(G91), .A2(n638), .ZN(n587) );
  NAND2_X1 U653 ( .A1(G53), .A2(n636), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G65), .A2(n639), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT69), .B(n588), .ZN(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n593), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n594), .B(KEYINPUT78), .ZN(n596) );
  NOR2_X1 U661 ( .A1(G299), .A2(G868), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n614), .A2(G559), .ZN(n597) );
  INV_X1 U664 ( .A(n917), .ZN(n612) );
  NAND2_X1 U665 ( .A1(n597), .A2(n612), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(n932), .A2(G868), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G868), .A2(n612), .ZN(n599) );
  NOR2_X1 U669 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G123), .A2(n870), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G111), .A2(n868), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT79), .B(n603), .Z(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G99), .A2(n864), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G135), .A2(n865), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n998) );
  XNOR2_X1 U680 ( .A(n998), .B(G2096), .ZN(n611) );
  INV_X1 U681 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U683 ( .A1(G559), .A2(n612), .ZN(n613) );
  XOR2_X1 U684 ( .A(n932), .B(n613), .Z(n655) );
  NAND2_X1 U685 ( .A1(n614), .A2(n655), .ZN(n623) );
  NAND2_X1 U686 ( .A1(G55), .A2(n636), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G67), .A2(n639), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n638), .A2(G93), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n617), .B(KEYINPUT80), .ZN(n619) );
  NAND2_X1 U691 ( .A1(G80), .A2(n642), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n620), .Z(n621) );
  NOR2_X1 U694 ( .A1(n622), .A2(n621), .ZN(n659) );
  XOR2_X1 U695 ( .A(n623), .B(n659), .Z(G145) );
  NAND2_X1 U696 ( .A1(G49), .A2(n636), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U699 ( .A1(n639), .A2(n626), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G87), .A2(n627), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(G288) );
  AND2_X1 U702 ( .A1(n636), .A2(G47), .ZN(n633) );
  NAND2_X1 U703 ( .A1(G85), .A2(n638), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G72), .A2(n642), .ZN(n630) );
  NAND2_X1 U705 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U707 ( .A1(n639), .A2(G60), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U709 ( .A1(G48), .A2(n636), .ZN(n637) );
  XNOR2_X1 U710 ( .A(n637), .B(KEYINPUT82), .ZN(n647) );
  NAND2_X1 U711 ( .A1(G86), .A2(n638), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n642), .A2(G73), .ZN(n643) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U718 ( .A(KEYINPUT83), .B(n648), .Z(G305) );
  XNOR2_X1 U719 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n650) );
  INV_X1 U720 ( .A(G299), .ZN(n925) );
  XNOR2_X1 U721 ( .A(G288), .B(n925), .ZN(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n659), .B(n651), .ZN(n653) );
  XNOR2_X1 U724 ( .A(G290), .B(G166), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(G305), .ZN(n890) );
  XNOR2_X1 U727 ( .A(n890), .B(KEYINPUT85), .ZN(n656) );
  XNOR2_X1 U728 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U729 ( .A1(G868), .A2(n657), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT86), .ZN(n661) );
  OR2_X1 U731 ( .A1(n659), .A2(G868), .ZN(n660) );
  NAND2_X1 U732 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XOR2_X1 U738 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U739 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U741 ( .A1(G108), .A2(G120), .ZN(n666) );
  NOR2_X1 U742 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U743 ( .A1(G69), .A2(n667), .ZN(n912) );
  NAND2_X1 U744 ( .A1(G567), .A2(n912), .ZN(n673) );
  NOR2_X1 U745 ( .A1(G219), .A2(G220), .ZN(n669) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(KEYINPUT87), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U748 ( .A1(n670), .A2(G218), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G96), .A2(n671), .ZN(n913) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n913), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U752 ( .A(KEYINPUT88), .B(n674), .Z(G319) );
  INV_X1 U753 ( .A(G319), .ZN(n676) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U755 ( .A1(n676), .A2(n675), .ZN(n824) );
  NAND2_X1 U756 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(n864), .A2(G102), .ZN(n679) );
  NAND2_X1 U758 ( .A1(G114), .A2(n868), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT89), .B(n677), .Z(n678) );
  NAND2_X1 U760 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G138), .A2(n865), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G126), .A2(n870), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n683), .A2(n682), .ZN(G164) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U766 ( .A(G1981), .B(KEYINPUT99), .ZN(n684) );
  XNOR2_X1 U767 ( .A(n684), .B(G305), .ZN(n922) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n770) );
  AND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n685) );
  NAND2_X1 U770 ( .A1(G8), .A2(n733), .ZN(n766) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n915) );
  INV_X1 U772 ( .A(n915), .ZN(n686) );
  NOR2_X1 U773 ( .A1(n766), .A2(n686), .ZN(n687) );
  NOR2_X1 U774 ( .A1(KEYINPUT33), .A2(n687), .ZN(n691) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n752) );
  NAND2_X1 U776 ( .A1(KEYINPUT33), .A2(n752), .ZN(n688) );
  XNOR2_X1 U777 ( .A(KEYINPUT98), .B(n688), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n766), .A2(n689), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n692) );
  AND2_X1 U780 ( .A1(n922), .A2(n692), .ZN(n756) );
  XNOR2_X1 U781 ( .A(G2078), .B(KEYINPUT25), .ZN(n954) );
  NOR2_X1 U782 ( .A1(n733), .A2(n954), .ZN(n694) );
  INV_X1 U783 ( .A(n733), .ZN(n705) );
  INV_X1 U784 ( .A(G1961), .ZN(n978) );
  NOR2_X1 U785 ( .A1(n705), .A2(n978), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n720) );
  AND2_X1 U787 ( .A1(G171), .A2(n720), .ZN(n695) );
  XNOR2_X1 U788 ( .A(n695), .B(KEYINPUT93), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n705), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U791 ( .A(G1956), .ZN(n965) );
  NOR2_X1 U792 ( .A1(n965), .A2(n705), .ZN(n697) );
  NOR2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n925), .A2(n700), .ZN(n699) );
  XOR2_X1 U795 ( .A(n699), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U796 ( .A1(n925), .A2(n700), .ZN(n714) );
  INV_X1 U797 ( .A(G1996), .ZN(n948) );
  NOR2_X1 U798 ( .A1(n733), .A2(n948), .ZN(n701) );
  XOR2_X1 U799 ( .A(n701), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U800 ( .A1(n733), .A2(G1341), .ZN(n702) );
  NAND2_X1 U801 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U802 ( .A1(n932), .A2(n704), .ZN(n709) );
  NAND2_X1 U803 ( .A1(G1348), .A2(n733), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n705), .A2(G2067), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n917), .A2(n710), .ZN(n708) );
  OR2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n917), .A2(n710), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U812 ( .A(KEYINPUT29), .B(n717), .Z(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n730) );
  NOR2_X1 U814 ( .A1(G171), .A2(n720), .ZN(n726) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n733), .ZN(n743) );
  NOR2_X1 U816 ( .A1(n746), .A2(n743), .ZN(n721) );
  XNOR2_X1 U817 ( .A(n721), .B(KEYINPUT94), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n722), .A2(G8), .ZN(n723) );
  XNOR2_X1 U819 ( .A(n723), .B(KEYINPUT30), .ZN(n724) );
  NOR2_X1 U820 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U822 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n731), .B(KEYINPUT96), .ZN(n744) );
  NAND2_X1 U825 ( .A1(n744), .A2(G286), .ZN(n740) );
  INV_X1 U826 ( .A(G8), .ZN(n738) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n766), .ZN(n732) );
  XNOR2_X1 U828 ( .A(KEYINPUT97), .B(n732), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U830 ( .A1(G166), .A2(n734), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U834 ( .A(n742), .B(n741), .ZN(n750) );
  NAND2_X1 U835 ( .A1(G8), .A2(n743), .ZN(n748) );
  INV_X1 U836 ( .A(n744), .ZN(n745) );
  NOR2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n759) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n916) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n753) );
  AND2_X1 U843 ( .A1(n916), .A2(n753), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n759), .A2(n754), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n762) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n760), .A2(n766), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(n763), .B(KEYINPUT100), .ZN(n768) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U853 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n774) );
  NAND2_X1 U856 ( .A1(G160), .A2(G40), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n817) );
  NOR2_X1 U858 ( .A1(G1986), .A2(G290), .ZN(n805) );
  INV_X1 U859 ( .A(n805), .ZN(n920) );
  NAND2_X1 U860 ( .A1(G1986), .A2(G290), .ZN(n930) );
  NAND2_X1 U861 ( .A1(n920), .A2(n930), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n817), .A2(n771), .ZN(n772) );
  XOR2_X1 U863 ( .A(KEYINPUT90), .B(n772), .Z(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n803) );
  NAND2_X1 U865 ( .A1(G117), .A2(n868), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G129), .A2(n870), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n864), .A2(G105), .ZN(n777) );
  XOR2_X1 U869 ( .A(KEYINPUT38), .B(n777), .Z(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U871 ( .A1(n865), .A2(G141), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n854) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n854), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G107), .A2(n868), .ZN(n783) );
  NAND2_X1 U875 ( .A1(G119), .A2(n870), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G95), .A2(n864), .ZN(n785) );
  NAND2_X1 U878 ( .A1(G131), .A2(n865), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n879) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n879), .ZN(n788) );
  NAND2_X1 U882 ( .A1(n789), .A2(n788), .ZN(n1001) );
  NAND2_X1 U883 ( .A1(n817), .A2(n1001), .ZN(n790) );
  XOR2_X1 U884 ( .A(KEYINPUT92), .B(n790), .Z(n808) );
  INV_X1 U885 ( .A(n808), .ZN(n801) );
  XOR2_X1 U886 ( .A(G2067), .B(KEYINPUT37), .Z(n816) );
  NAND2_X1 U887 ( .A1(G104), .A2(n864), .ZN(n792) );
  NAND2_X1 U888 ( .A1(G140), .A2(n865), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U890 ( .A(KEYINPUT34), .B(n793), .ZN(n799) );
  NAND2_X1 U891 ( .A1(G116), .A2(n868), .ZN(n795) );
  NAND2_X1 U892 ( .A1(G128), .A2(n870), .ZN(n794) );
  NAND2_X1 U893 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U894 ( .A(KEYINPUT35), .B(n796), .ZN(n797) );
  XNOR2_X1 U895 ( .A(KEYINPUT91), .B(n797), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U897 ( .A(KEYINPUT36), .B(n800), .Z(n886) );
  AND2_X1 U898 ( .A1(n816), .A2(n886), .ZN(n1019) );
  NAND2_X1 U899 ( .A1(n1019), .A2(n817), .ZN(n804) );
  AND2_X1 U900 ( .A1(n801), .A2(n804), .ZN(n802) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n815) );
  INV_X1 U902 ( .A(n804), .ZN(n813) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n854), .ZN(n1005) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n879), .ZN(n999) );
  NOR2_X1 U905 ( .A1(n999), .A2(n805), .ZN(n806) );
  XOR2_X1 U906 ( .A(KEYINPUT101), .B(n806), .Z(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n1005), .A2(n809), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n810), .B(KEYINPUT39), .ZN(n811) );
  NAND2_X1 U910 ( .A1(n811), .A2(n817), .ZN(n812) );
  OR2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  AND2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n816), .A2(n886), .ZN(n1015) );
  NAND2_X1 U914 ( .A1(n1015), .A2(n817), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U922 ( .A(G2100), .B(G2096), .Z(n826) );
  XNOR2_X1 U923 ( .A(KEYINPUT42), .B(G2678), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT43), .B(G2090), .Z(n828) );
  XNOR2_X1 U926 ( .A(G2067), .B(G2072), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U928 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U929 ( .A(G2078), .B(G2084), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(G227) );
  XOR2_X1 U931 ( .A(G1966), .B(G1981), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n844) );
  XOR2_X1 U934 ( .A(KEYINPUT41), .B(G2474), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1956), .B(KEYINPUT104), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(G1961), .B(G1971), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1976), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G124), .A2(n870), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U946 ( .A1(G112), .A2(n868), .ZN(n846) );
  XOR2_X1 U947 ( .A(KEYINPUT107), .B(n846), .Z(n847) );
  NAND2_X1 U948 ( .A1(n848), .A2(n847), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G100), .A2(n864), .ZN(n850) );
  NAND2_X1 U950 ( .A1(G136), .A2(n865), .ZN(n849) );
  NAND2_X1 U951 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(G162) );
  XOR2_X1 U953 ( .A(G162), .B(n998), .Z(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n863) );
  NAND2_X1 U955 ( .A1(G118), .A2(n868), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G130), .A2(n870), .ZN(n855) );
  NAND2_X1 U957 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G106), .A2(n864), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G142), .A2(n865), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(KEYINPUT45), .B(n859), .Z(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n863), .B(n862), .Z(n878) );
  NAND2_X1 U964 ( .A1(G103), .A2(n864), .ZN(n867) );
  NAND2_X1 U965 ( .A1(G139), .A2(n865), .ZN(n866) );
  NAND2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n876) );
  NAND2_X1 U967 ( .A1(n868), .A2(G115), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n869), .B(KEYINPUT108), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G127), .A2(n870), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(KEYINPUT109), .B(n873), .ZN(n874) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n874), .ZN(n875) );
  NOR2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n1010) );
  XNOR2_X1 U974 ( .A(G164), .B(n1010), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n888) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U979 ( .A(n882), .B(KEYINPUT110), .Z(n884) );
  XNOR2_X1 U980 ( .A(G160), .B(KEYINPUT111), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n886), .B(n885), .Z(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n889) );
  NOR2_X1 U984 ( .A1(G37), .A2(n889), .ZN(G395) );
  XNOR2_X1 U985 ( .A(n890), .B(KEYINPUT113), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n917), .B(G171), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U988 ( .A(G286), .B(n932), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G397) );
  XNOR2_X1 U991 ( .A(G2451), .B(G2427), .ZN(n905) );
  XOR2_X1 U992 ( .A(G2430), .B(G2443), .Z(n897) );
  XNOR2_X1 U993 ( .A(KEYINPUT103), .B(G2438), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n899) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2446), .B(KEYINPUT102), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U1002 ( .A1(n906), .A2(G14), .ZN(n914) );
  NAND2_X1 U1003 ( .A1(n914), .A2(G319), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(G225) );
  XOR2_X1 U1009 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  INV_X1 U1017 ( .A(n914), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G16), .B(KEYINPUT56), .Z(n942) );
  NAND2_X1 U1019 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G1348), .B(n917), .ZN(n918) );
  NOR2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n939) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G168), .ZN(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(n924), .B(KEYINPUT57), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(G1956), .B(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(G1971), .A2(G303), .ZN(n926) );
  NAND2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G1961), .B(G301), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n932), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT118), .B(n933), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT119), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n996) );
  XOR2_X1 U1039 ( .A(G2090), .B(G35), .Z(n945) );
  XOR2_X1 U1040 ( .A(KEYINPUT54), .B(G34), .Z(n943) );
  XNOR2_X1 U1041 ( .A(G2084), .B(n943), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n959) );
  XNOR2_X1 U1043 ( .A(G2067), .B(G26), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G32), .B(n948), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n949), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G25), .B(G1991), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n956) );
  XOR2_X1 U1051 ( .A(G27), .B(n954), .Z(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT53), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT55), .B(n960), .ZN(n962) );
  INV_X1 U1056 ( .A(G29), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(G11), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT117), .ZN(n994) );
  XOR2_X1 U1060 ( .A(G16), .B(KEYINPUT120), .Z(n992) );
  XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(KEYINPUT124), .ZN(n990) );
  XNOR2_X1 U1062 ( .A(G20), .B(n965), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G6), .ZN(n967) );
  XNOR2_X1 U1064 ( .A(G1341), .B(G19), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1066 ( .A(KEYINPUT121), .B(n968), .Z(n969) );
  NAND2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n971) );
  XNOR2_X1 U1069 ( .A(G4), .B(n971), .ZN(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1071 ( .A(KEYINPUT60), .B(n974), .Z(n976) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G21), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(KEYINPUT122), .B(n977), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n978), .B(G5), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n988) );
  XOR2_X1 U1077 ( .A(G1986), .B(G24), .Z(n984) );
  XNOR2_X1 U1078 ( .A(G1976), .B(G23), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n981) );
  NOR2_X1 U1080 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1082 ( .A(KEYINPUT123), .B(n985), .Z(n986) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(n986), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(n990), .B(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT125), .B(n997), .ZN(n1026) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(G160), .B(G2084), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G2090), .B(G162), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT115), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT51), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1017) );
  XOR2_X1 U1099 ( .A(G2072), .B(n1010), .Z(n1012) );
  XOR2_X1 U1100 ( .A(G164), .B(G2078), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1013), .Z(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1020), .ZN(n1022) );
  INV_X1 U1107 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(n1024), .B(KEYINPUT116), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .Z(n1028) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(n1028), .Z(G311) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

