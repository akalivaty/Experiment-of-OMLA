//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(G250), .B1(G257), .B2(G264), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(KEYINPUT0), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT64), .B(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  OR3_X1    g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n231), .A2(new_n232), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n212), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n225), .B(new_n240), .C1(KEYINPUT1), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT2), .B(G226), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G13), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n258), .A2(new_n210), .A3(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n222), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n209), .A2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(new_n267), .B2(KEYINPUT75), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(KEYINPUT75), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(new_n269), .B1(new_n259), .B2(new_n264), .ZN(new_n270));
  INV_X1    g0070(.A(new_n261), .ZN(new_n271));
  AND2_X1   g0071(.A1(G58), .A2(G68), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n272), .B2(new_n201), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G159), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n277), .B1(new_n282), .B2(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT64), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G20), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(KEYINPUT7), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n227), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n277), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT73), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT3), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT7), .B1(new_n293), .B2(G20), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n276), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n271), .B1(new_n295), .B2(KEYINPUT16), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n279), .A2(new_n281), .A3(new_n292), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT7), .A4(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n301), .A2(new_n277), .A3(G20), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n298), .A2(new_n300), .B1(new_n302), .B2(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G68), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n276), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT7), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n221), .B(new_n308), .C1(new_n282), .C2(KEYINPUT3), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n290), .A2(new_n210), .A3(new_n299), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n227), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT74), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT16), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n270), .B1(new_n297), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT76), .ZN(new_n317));
  INV_X1    g0117(.A(G223), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n283), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G87), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n293), .A2(G226), .A3(G1698), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n292), .B1(new_n279), .B2(new_n281), .ZN(new_n324));
  OAI211_X1 g0124(.A(KEYINPUT76), .B(new_n319), .C1(new_n324), .C2(new_n277), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n321), .A2(new_n322), .A3(new_n323), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G41), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G1), .A3(G13), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(G274), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT68), .ZN(new_n333));
  NOR2_X1   g0133(.A1(G41), .A2(G45), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(G1), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n209), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT69), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n334), .B2(G1), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n209), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n328), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n338), .B1(new_n243), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n343), .B1(new_n326), .B2(new_n329), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT77), .ZN(new_n349));
  AOI21_X1  g0149(.A(G200), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G190), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n316), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT17), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT77), .B1(new_n330), .B2(new_n344), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n346), .B(new_n343), .C1(new_n326), .C2(new_n329), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n348), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n315), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT18), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT18), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n360), .A2(new_n315), .A3(new_n365), .A4(new_n362), .ZN(new_n366));
  INV_X1    g0166(.A(G200), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n358), .B2(new_n359), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n315), .B1(new_n368), .B2(new_n352), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT17), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n356), .A2(new_n364), .A3(new_n366), .A4(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n221), .A2(G33), .A3(G77), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n227), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n271), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n374), .A2(KEYINPUT11), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n262), .A2(G68), .A3(new_n266), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n376), .B(KEYINPUT71), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n259), .A2(new_n227), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT12), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(KEYINPUT11), .ZN(new_n380));
  AND4_X1   g0180(.A1(new_n375), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT72), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT14), .ZN(new_n383));
  INV_X1    g0183(.A(G1698), .ZN(new_n384));
  OAI211_X1 g0184(.A(G226), .B(new_n384), .C1(new_n301), .C2(new_n277), .ZN(new_n385));
  OAI211_X1 g0185(.A(G232), .B(G1698), .C1(new_n301), .C2(new_n277), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(new_n329), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n340), .A2(new_n328), .A3(G238), .A4(new_n341), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n338), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT13), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n340), .A2(new_n328), .A3(new_n341), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(G238), .B1(new_n332), .B2(new_n337), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n388), .A2(new_n329), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n383), .B(G169), .C1(new_n392), .C2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n389), .B2(new_n391), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n393), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(G179), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n399), .A2(new_n400), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n383), .B1(new_n403), .B2(G169), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n382), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(G169), .B1(new_n392), .B2(new_n397), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT14), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(KEYINPUT72), .A3(new_n401), .A4(new_n398), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n381), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n266), .A2(G77), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n263), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n229), .B2(new_n259), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n221), .A2(G33), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n274), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n229), .A2(new_n221), .B1(new_n264), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n261), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n290), .A2(new_n299), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G232), .A3(new_n384), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(G1698), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n421), .B1(new_n206), .B2(new_n420), .C1(new_n422), .C2(new_n228), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n329), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n338), .B1(new_n230), .B2(new_n342), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT70), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT70), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n338), .B(new_n427), .C1(new_n230), .C2(new_n342), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n419), .B1(new_n429), .B2(G200), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n351), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n357), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n419), .C1(G179), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n420), .A2(G222), .A3(new_n384), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n436), .B1(new_n229), .B2(new_n420), .C1(new_n422), .C2(new_n318), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n329), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n394), .A2(G226), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n338), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n274), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n442), .B1(new_n413), .B2(new_n264), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n261), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n266), .A2(G50), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n262), .A2(new_n446), .B1(new_n202), .B2(new_n259), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT9), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n438), .A2(G190), .A3(new_n338), .A4(new_n439), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT9), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n441), .A2(new_n450), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT10), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n450), .A2(new_n453), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT10), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n451), .A4(new_n441), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n440), .A2(G179), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n440), .A2(new_n357), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n448), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n435), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n403), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G190), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n465), .B(new_n381), .C1(new_n367), .C2(new_n464), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NOR4_X1   g0267(.A1(new_n371), .A2(new_n409), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT21), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n258), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n278), .A2(G1), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n259), .A2(new_n261), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(G116), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n260), .A2(new_n222), .B1(G20), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n278), .A2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n287), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n221), .A2(new_n479), .A3(new_n478), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n475), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G169), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n328), .A3(G274), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n328), .ZN(new_n493));
  INV_X1    g0293(.A(G270), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(G257), .B(new_n384), .C1(new_n324), .C2(new_n277), .ZN(new_n496));
  OAI211_X1 g0296(.A(G264), .B(G1698), .C1(new_n324), .C2(new_n277), .ZN(new_n497));
  INV_X1    g0297(.A(new_n420), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G303), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n495), .B1(new_n500), .B2(new_n329), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n469), .B1(new_n487), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n329), .ZN(new_n503));
  INV_X1    g0303(.A(new_n495), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n481), .A2(new_n482), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n477), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n357), .B1(new_n508), .B2(new_n475), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(KEYINPUT21), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(G179), .A3(new_n486), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n501), .A2(G190), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n486), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n501), .B2(new_n367), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT85), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n487), .A2(new_n501), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n361), .B(new_n495), .C1(new_n329), .C2(new_n500), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n519), .A2(KEYINPUT21), .B1(new_n520), .B2(new_n486), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT85), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n513), .B(new_n515), .C1(new_n367), .C2(new_n501), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n502), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT4), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n230), .A2(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n283), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(KEYINPUT4), .C1(new_n277), .C2(new_n301), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(G1698), .C1(new_n301), .C2(new_n277), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n479), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n328), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G257), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n491), .B1(new_n493), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n357), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n206), .A2(G97), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G97), .A2(G107), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n207), .A2(new_n539), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n287), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n274), .A2(G77), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n206), .B1(new_n309), .B2(new_n311), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n261), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n471), .A2(G97), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n474), .B2(G97), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT4), .B1(new_n293), .B2(new_n527), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n329), .B1(new_n555), .B2(new_n532), .ZN(new_n556));
  INV_X1    g0356(.A(new_n536), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n361), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n537), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT80), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT80), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n537), .A2(new_n554), .A3(new_n561), .A4(new_n558), .ZN(new_n562));
  INV_X1    g0362(.A(new_n553), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n303), .A2(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(new_n548), .A3(new_n547), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n565), .B2(new_n261), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n534), .A2(G190), .A3(new_n536), .ZN(new_n568));
  AOI21_X1  g0368(.A(G200), .B1(new_n556), .B2(new_n557), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n556), .A2(new_n351), .A3(new_n557), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n529), .A2(new_n533), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n536), .B1(new_n573), .B2(new_n329), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n572), .B1(new_n574), .B2(G200), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n567), .B1(new_n575), .B2(new_n566), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n560), .B(new_n562), .C1(new_n571), .C2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n284), .B(new_n286), .C1(new_n578), .C2(new_n387), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n205), .A3(new_n206), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n284), .A2(new_n286), .A3(G33), .A4(G97), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n579), .A2(new_n581), .B1(new_n582), .B2(new_n578), .ZN(new_n583));
  OAI211_X1 g0383(.A(G68), .B(new_n221), .C1(new_n324), .C2(new_n277), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n261), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n414), .A2(new_n259), .ZN(new_n587));
  INV_X1    g0387(.A(new_n414), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n474), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT83), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n586), .A2(new_n592), .A3(new_n587), .A4(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(G244), .B(G1698), .C1(new_n324), .C2(new_n277), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT82), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT82), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n293), .A2(new_n597), .A3(G244), .A4(G1698), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n282), .A2(G116), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n293), .A2(G238), .A3(new_n384), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n329), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n328), .A2(G274), .A3(new_n490), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT81), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(G250), .B1(new_n489), .B2(G1), .ZN(new_n607));
  OAI22_X1  g0407(.A1(new_n605), .A2(new_n606), .B1(new_n329), .B2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n357), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n601), .B2(new_n329), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n361), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n594), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT84), .B1(new_n474), .B2(G87), .ZN(new_n615));
  INV_X1    g0415(.A(new_n474), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n616), .A2(new_n617), .A3(new_n580), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n586), .B(new_n587), .C1(new_n615), .C2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(G190), .B2(new_n612), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n610), .A2(G200), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g0423(.A(G257), .B(G1698), .C1(new_n324), .C2(new_n277), .ZN(new_n624));
  OAI211_X1 g0424(.A(G250), .B(new_n384), .C1(new_n324), .C2(new_n277), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n282), .A2(G294), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n329), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n492), .A2(G264), .A3(new_n328), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n491), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n367), .ZN(new_n631));
  INV_X1    g0431(.A(new_n629), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n627), .B2(new_n329), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n351), .A3(new_n491), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT25), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n471), .B2(G107), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n637), .B(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n206), .B2(new_n616), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n293), .A2(KEYINPUT22), .A3(G87), .A4(new_n221), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n420), .A2(new_n221), .A3(G87), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT22), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n282), .A2(new_n210), .A3(G116), .ZN(new_n646));
  NOR2_X1   g0446(.A1(KEYINPUT23), .A2(G107), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n206), .A2(G20), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n287), .A2(new_n647), .B1(KEYINPUT23), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n642), .A2(new_n645), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(KEYINPUT24), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n649), .A2(new_n646), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT24), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n642), .A3(new_n653), .A4(new_n645), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n641), .B1(new_n655), .B2(new_n261), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n635), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n630), .A2(new_n357), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n633), .A2(new_n361), .A3(new_n491), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n271), .B1(new_n651), .B2(new_n654), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n658), .B(new_n659), .C1(new_n660), .C2(new_n641), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n577), .A2(new_n623), .A3(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n468), .A2(new_n525), .A3(new_n663), .ZN(G372));
  AOI22_X1  g0464(.A1(new_n591), .A2(new_n593), .B1(new_n361), .B2(new_n612), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT87), .B1(new_n610), .B2(new_n357), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n612), .A2(new_n667), .A3(G169), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n665), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n665), .B(new_n671), .C1(new_n666), .C2(new_n668), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n661), .A2(new_n502), .A3(new_n521), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n574), .A2(new_n361), .B1(new_n551), .B2(new_n553), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n561), .B1(new_n674), .B2(new_n537), .ZN(new_n675));
  INV_X1    g0475(.A(new_n562), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT79), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n570), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n673), .A2(new_n677), .A3(new_n680), .A4(new_n657), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n669), .A2(new_n622), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n670), .B(new_n672), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n560), .A2(new_n562), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n614), .A3(KEYINPUT26), .A4(new_n622), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n559), .B(KEYINPUT89), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n688), .A2(new_n669), .A3(new_n622), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n686), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n468), .B1(new_n683), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n369), .B(new_n355), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n433), .B(KEYINPUT90), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n467), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n692), .B1(new_n694), .B2(new_n409), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n364), .A2(new_n366), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n459), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(new_n462), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n691), .A2(new_n700), .ZN(G369));
  NAND2_X1  g0501(.A1(new_n221), .A2(new_n470), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT27), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(G213), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n512), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n662), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n661), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n710), .A2(new_n515), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n518), .B2(new_n524), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n715), .A2(new_n512), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  OAI211_X1 g0521(.A(new_n657), .B(new_n661), .C1(new_n656), .C2(new_n710), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n713), .A2(new_n709), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n714), .B1(new_n721), .B2(new_n725), .ZN(G399));
  NOR2_X1   g0526(.A1(new_n214), .A2(G41), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n209), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n581), .A2(G116), .ZN(new_n729));
  INV_X1    g0529(.A(new_n220), .ZN(new_n730));
  AOI22_X1  g0530(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n727), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT28), .Z(new_n732));
  AND4_X1   g0532(.A1(new_n614), .A2(new_n622), .A3(new_n657), .A4(new_n661), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n684), .B1(new_n679), .B2(new_n570), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n733), .A2(new_n734), .A3(new_n525), .A4(new_n710), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n663), .A2(KEYINPUT94), .A3(new_n525), .A4(new_n710), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(G179), .B1(new_n556), .B2(new_n557), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n610), .A2(new_n505), .A3(new_n630), .A4(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT93), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n574), .A2(new_n633), .A3(new_n501), .A4(G179), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(new_n610), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n574), .A2(new_n633), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(KEYINPUT30), .A3(new_n520), .A4(new_n612), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n574), .A2(new_n501), .A3(G179), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(KEYINPUT93), .A3(new_n610), .A4(new_n630), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n743), .A2(new_n746), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n709), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT31), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n748), .A2(new_n746), .A3(new_n741), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n739), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n710), .B1(new_n690), .B2(new_n683), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT29), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n687), .B1(new_n623), .B2(new_n677), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n688), .A2(new_n669), .A3(KEYINPUT26), .A4(new_n622), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT29), .B(new_n710), .C1(new_n765), .C2(new_n683), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT95), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n670), .A2(new_n672), .ZN(new_n769));
  AND4_X1   g0569(.A1(new_n677), .A2(new_n673), .A3(new_n680), .A4(new_n657), .ZN(new_n770));
  INV_X1    g0570(.A(new_n682), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n764), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n773), .A2(KEYINPUT95), .A3(KEYINPUT29), .A4(new_n710), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n758), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n732), .B1(new_n776), .B2(G1), .ZN(G364));
  NOR2_X1   g0577(.A1(new_n287), .A2(new_n258), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G45), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n728), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n718), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n721), .B(new_n780), .C1(G330), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n780), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n213), .A2(new_n420), .ZN(new_n784));
  INV_X1    g0584(.A(G355), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n785), .B1(G116), .B2(new_n213), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n253), .A2(new_n489), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n283), .A2(new_n213), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n489), .B2(new_n730), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n222), .B1(G20), .B2(new_n357), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n783), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n221), .A2(new_n361), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n351), .A2(G200), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n367), .A2(G179), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n804), .A2(new_n210), .A3(new_n351), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n420), .B(new_n802), .C1(G303), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G326), .ZN(new_n807));
  INV_X1    g0607(.A(new_n798), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(new_n351), .A3(new_n367), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n808), .A2(G190), .A3(new_n367), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XOR2_X1   g0612(.A(KEYINPUT33), .B(G317), .Z(new_n813));
  OAI221_X1 g0613(.A(new_n806), .B1(new_n807), .B2(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n221), .B1(new_n361), .B2(new_n799), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n221), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(G294), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n221), .A2(new_n804), .A3(G190), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G190), .A2(G200), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n798), .A2(new_n823), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n818), .B1(new_n819), .B2(new_n821), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n817), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  OR3_X1    g0627(.A1(new_n826), .A2(KEYINPUT32), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT32), .B1(new_n826), .B2(new_n827), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n227), .C2(new_n812), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n821), .A2(new_n206), .ZN(new_n831));
  INV_X1    g0631(.A(new_n805), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n832), .A2(new_n580), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n831), .A2(new_n833), .A3(new_n498), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n815), .A2(new_n205), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n800), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G58), .A2(new_n837), .B1(new_n838), .B2(G77), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n809), .A2(G50), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n834), .A2(new_n836), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n814), .A2(new_n825), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n797), .B1(new_n842), .B2(new_n794), .ZN(new_n843));
  INV_X1    g0643(.A(new_n793), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n781), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n782), .A2(new_n845), .ZN(G396));
  NAND2_X1  g0646(.A1(new_n709), .A2(new_n419), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n435), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n693), .B2(new_n847), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n759), .A2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(KEYINPUT97), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(KEYINPUT97), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n434), .A2(new_n709), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n689), .A2(new_n687), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n685), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n772), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n780), .B1(new_n860), .B2(new_n758), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n855), .B1(new_n690), .B2(new_n683), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n758), .B(new_n862), .C1(new_n852), .C2(new_n853), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n794), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n792), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n783), .B1(G77), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT96), .ZN(new_n869));
  AOI22_X1  g0669(.A1(G143), .A2(new_n837), .B1(new_n838), .B2(G159), .ZN(new_n870));
  INV_X1    g0670(.A(G150), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n870), .B1(new_n812), .B2(new_n871), .C1(new_n872), .C2(new_n810), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT34), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n820), .A2(G68), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n283), .B1(G50), .B2(new_n805), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n816), .A2(G58), .B1(new_n817), .B2(G132), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n498), .B1(new_n832), .B2(new_n206), .ZN(new_n879));
  AOI211_X1 g0679(.A(new_n835), .B(new_n879), .C1(G303), .C2(new_n809), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n838), .A2(G116), .B1(G87), .B2(new_n820), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n837), .A2(G294), .B1(G311), .B2(new_n817), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n811), .A2(G283), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n869), .B1(new_n885), .B2(new_n866), .C1(new_n792), .C2(new_n849), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n865), .A2(new_n886), .ZN(G384));
  NOR3_X1   g0687(.A1(new_n221), .A2(new_n476), .A3(new_n222), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n544), .A2(new_n546), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT35), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n889), .ZN(new_n892));
  XNOR2_X1  g0692(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n892), .B(new_n893), .ZN(new_n894));
  OR3_X1    g0694(.A1(new_n220), .A2(new_n229), .A3(new_n272), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n202), .A2(G68), .ZN(new_n896));
  AOI211_X1 g0696(.A(new_n209), .B(G13), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n463), .A2(new_n409), .A3(new_n467), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n696), .A3(new_n692), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n759), .B2(new_n760), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n699), .B1(new_n775), .B2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(new_n707), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n315), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n354), .A2(new_n906), .A3(new_n363), .A4(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n295), .A2(KEYINPUT16), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n270), .B1(new_n297), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n360), .A2(new_n362), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT101), .B1(new_n913), .B2(new_n369), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT101), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n360), .A2(new_n362), .A3(new_n912), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n354), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n907), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n910), .B1(new_n919), .B2(KEYINPUT37), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n918), .B1(new_n692), .B2(new_n696), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n908), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n371), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n363), .A2(new_n908), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT37), .B1(new_n926), .B2(new_n369), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n909), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n905), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n409), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n709), .ZN(new_n932));
  INV_X1    g0732(.A(new_n918), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n371), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n354), .A2(new_n916), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(KEYINPUT101), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n906), .B1(new_n936), .B2(new_n917), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT38), .B(new_n934), .C1(new_n937), .C2(new_n910), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n922), .B1(new_n920), .B2(new_n921), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT39), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n930), .A2(new_n932), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT99), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n433), .A2(new_n709), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n859), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n862), .A2(KEYINPUT99), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n405), .A2(new_n466), .A3(new_n408), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT100), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n710), .A2(new_n381), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(KEYINPUT100), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n409), .A2(new_n467), .A3(new_n950), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n938), .A2(new_n939), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n947), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n696), .A2(new_n907), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n941), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n904), .B(new_n961), .Z(new_n962));
  OAI211_X1 g0762(.A(new_n849), .B(new_n951), .C1(new_n953), .C2(new_n954), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n754), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n739), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n923), .B2(new_n929), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n965), .B1(new_n737), .B2(new_n738), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n969), .A2(KEYINPUT40), .A3(new_n963), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(KEYINPUT40), .B1(new_n957), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n969), .A2(new_n900), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n971), .B1(new_n900), .B2(new_n969), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(G330), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n962), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n209), .B2(new_n778), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n962), .A2(new_n976), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n898), .B1(new_n978), .B2(new_n979), .ZN(G367));
  XOR2_X1   g0780(.A(new_n727), .B(KEYINPUT41), .Z(new_n981));
  OAI21_X1  g0781(.A(new_n734), .B1(new_n566), .B2(new_n710), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n559), .B2(new_n710), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n714), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT45), .Z(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n714), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT105), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n721), .A2(new_n725), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n725), .A2(new_n711), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT106), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT106), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(new_n995), .C1(new_n662), .C2(new_n711), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n721), .B(new_n996), .Z(new_n997));
  NAND3_X1  g0797(.A1(new_n992), .A2(new_n776), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n981), .B1(new_n998), .B2(new_n776), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n779), .A2(G1), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n709), .A2(new_n619), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n682), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n769), .B2(new_n1002), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT43), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n983), .A2(new_n712), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT42), .Z(new_n1008));
  AND2_X1   g0808(.A1(new_n983), .A2(new_n713), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n710), .B1(new_n1009), .B2(new_n684), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1006), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n991), .A2(new_n983), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1013), .B(new_n1014), .Z(new_n1015));
  AND2_X1   g0815(.A1(new_n1001), .A2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n795), .B1(new_n213), .B2(new_n414), .C1(new_n249), .C2(new_n788), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n809), .A2(G143), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n820), .A2(G77), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n498), .B1(new_n805), .B2(G58), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G159), .B2(new_n811), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n816), .A2(G68), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n817), .A2(G137), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G50), .A2(new_n838), .B1(new_n837), .B2(G150), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n837), .A2(G303), .B1(G317), .B2(new_n817), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n820), .A2(G97), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n819), .C2(new_n824), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n283), .B1(new_n815), .B2(new_n206), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n809), .B2(G311), .ZN(new_n1031));
  INV_X1    g0831(.A(G294), .ZN(new_n1032));
  AOI21_X1  g0832(.A(KEYINPUT107), .B1(new_n805), .B2(G116), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(KEYINPUT46), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(KEYINPUT46), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1031), .B1(new_n812), .B2(new_n1032), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1026), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT47), .Z(new_n1039));
  OAI211_X1 g0839(.A(new_n783), .B(new_n1017), .C1(new_n1039), .C2(new_n866), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1004), .B2(new_n793), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1016), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(G387));
  OAI22_X1  g0843(.A1(new_n784), .A2(new_n729), .B1(G107), .B2(new_n213), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n246), .A2(new_n489), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n729), .ZN(new_n1046));
  AOI211_X1 g0846(.A(G45), .B(new_n1046), .C1(G68), .C2(G77), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n264), .A2(G50), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n788), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1044), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(KEYINPUT108), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT108), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n795), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n783), .B1(new_n1052), .B2(new_n1054), .C1(new_n724), .C2(new_n844), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1028), .B(new_n293), .C1(new_n229), .C2(new_n832), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n265), .B2(new_n811), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n816), .A2(new_n588), .B1(new_n817), .B2(G150), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G50), .A2(new_n837), .B1(new_n838), .B2(G68), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n809), .A2(G159), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n816), .A2(G283), .B1(G294), .B2(new_n805), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G303), .A2(new_n838), .B1(new_n837), .B2(G317), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n812), .B2(new_n822), .C1(new_n801), .C2(new_n810), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT109), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n283), .B1(new_n821), .B2(new_n476), .C1(new_n807), .C2(new_n826), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT110), .Z(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT49), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1061), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT111), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1055), .B1(new_n1075), .B2(new_n794), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n997), .B2(new_n1000), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n997), .A2(new_n776), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n727), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n997), .A2(new_n776), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(KEYINPUT112), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n989), .B1(new_n991), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n991), .A2(new_n1082), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1085), .A2(KEYINPUT113), .B1(G1), .B2(new_n779), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(KEYINPUT113), .B2(new_n1085), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n795), .B1(new_n205), .B2(new_n213), .C1(new_n256), .C2(new_n788), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n783), .A2(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n809), .A2(G317), .B1(G311), .B2(new_n837), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n826), .A2(new_n801), .B1(new_n476), .B2(new_n815), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G294), .B2(new_n838), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n498), .B1(new_n832), .B2(new_n819), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1094), .B(new_n831), .C1(G303), .C2(new_n811), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n809), .A2(G150), .B1(G159), .B2(new_n837), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n293), .B1(new_n832), .B2(new_n227), .C1(new_n821), .C2(new_n580), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G50), .B2(new_n811), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n816), .A2(G77), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n838), .A2(new_n265), .B1(G143), .B2(new_n817), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1096), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n1104), .B2(new_n794), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n983), .B2(new_n844), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1085), .A2(new_n1078), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n998), .A2(new_n727), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1087), .B(new_n1106), .C1(new_n1107), .C2(new_n1108), .ZN(G390));
  NAND2_X1  g0909(.A1(new_n739), .A2(new_n966), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(G330), .A3(new_n468), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n973), .A2(KEYINPUT114), .A3(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1115), .A2(KEYINPUT115), .A3(new_n902), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n902), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n850), .A2(new_n719), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1110), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n955), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n956), .B1(new_n757), .B2(new_n1119), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n947), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n955), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n709), .B1(new_n772), .B2(new_n764), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n943), .B1(new_n1125), .B2(new_n849), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n757), .A2(new_n956), .A3(new_n1119), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1118), .A2(new_n1129), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n859), .A2(new_n942), .A3(new_n943), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT99), .B1(new_n862), .B2(new_n945), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n956), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n932), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(new_n1134), .B1(new_n930), .B2(new_n940), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1126), .A2(new_n955), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1137), .A2(new_n909), .B1(new_n371), .B2(new_n933), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n929), .B1(new_n1138), .B2(KEYINPUT38), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1136), .A2(new_n1139), .A3(new_n932), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1121), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1134), .B1(new_n923), .B2(new_n929), .C1(new_n955), .C2(new_n1126), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n955), .B1(new_n944), .B2(new_n946), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1143), .A2(new_n932), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT39), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n929), .ZN(new_n1146));
  AOI21_X1  g0946(.A(KEYINPUT39), .B1(new_n938), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1142), .B(new_n1127), .C1(new_n1144), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1141), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1130), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1118), .A2(new_n1149), .A3(new_n1141), .A4(new_n1129), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n727), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1141), .A2(new_n1149), .A3(new_n1000), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n783), .B1(new_n265), .B2(new_n867), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT54), .B(G143), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n826), .A2(new_n1156), .B1(new_n824), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n498), .B(new_n1158), .C1(G50), .C2(new_n820), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n809), .B1(new_n811), .B2(G137), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n805), .A2(G150), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G132), .B2(new_n837), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n827), .B2(new_n815), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n875), .B1(new_n826), .B2(new_n1032), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT116), .Z(new_n1167));
  AOI22_X1  g0967(.A1(G107), .A2(new_n811), .B1(new_n809), .B2(G283), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n833), .A2(new_n420), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G97), .A2(new_n838), .B1(new_n837), .B2(G116), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n1101), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1161), .A2(new_n1165), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1155), .B1(new_n1172), .B2(new_n794), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1148), .B2(new_n792), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1153), .A2(new_n1154), .A3(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(new_n1129), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1118), .B1(new_n1150), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT119), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n963), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1110), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT40), .B1(new_n1139), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n957), .A2(new_n970), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n719), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n961), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n959), .B1(new_n1143), .B2(new_n957), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n941), .C1(new_n971), .C2(new_n719), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n459), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n462), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n707), .A2(new_n449), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n449), .B(new_n707), .C1(new_n459), .C2(new_n462), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1193), .B(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT118), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1187), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1184), .A2(new_n1186), .A3(new_n1197), .A4(new_n1196), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT119), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1118), .C1(new_n1150), .C2(new_n1176), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1178), .A2(KEYINPUT57), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1204), .A2(new_n727), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT57), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1202), .B1(new_n1152), .B2(new_n1118), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT120), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1178), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1206), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1205), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1196), .A2(new_n791), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n783), .B1(G50), .B2(new_n867), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n826), .A2(new_n819), .B1(new_n206), .B2(new_n800), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n588), .B2(new_n838), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n816), .A2(G68), .B1(G77), .B2(new_n805), .ZN(new_n1219));
  INV_X1    g1019(.A(G41), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n283), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G58), .B2(new_n820), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G97), .A2(new_n811), .B1(new_n809), .B2(G116), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1218), .A2(new_n1219), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT58), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G50), .B1(new_n278), .B2(new_n1220), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1224), .A2(new_n1225), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n810), .A2(new_n1156), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1157), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n816), .A2(G150), .B1(new_n805), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G128), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1230), .B1(new_n800), .B2(new_n1231), .C1(new_n872), .C2(new_n824), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1228), .B(new_n1232), .C1(G132), .C2(new_n811), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT59), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(KEYINPUT117), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n278), .B(new_n1220), .C1(new_n821), .C2(new_n827), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G124), .B2(new_n817), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT117), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1238), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1227), .B1(new_n1225), .B2(new_n1224), .C1(new_n1236), .C2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1216), .B1(new_n1241), .B2(new_n794), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n1201), .A2(new_n1000), .B1(new_n1215), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1214), .A2(new_n1243), .ZN(G375));
  AOI21_X1  g1044(.A(new_n981), .B1(new_n1118), .B2(new_n1129), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1118), .B2(new_n1129), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n206), .A2(new_n824), .B1(new_n800), .B2(new_n819), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n816), .A2(new_n588), .B1(G97), .B2(new_n805), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n812), .B2(new_n476), .C1(new_n1032), .C2(new_n810), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1247), .B(new_n1249), .C1(G303), .C2(new_n817), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1019), .A2(new_n498), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT121), .Z(new_n1252));
  OAI22_X1  g1052(.A1(new_n826), .A2(new_n1231), .B1(new_n872), .B2(new_n800), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n824), .A2(new_n871), .B1(new_n815), .B2(new_n202), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n820), .A2(G58), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n283), .B1(G159), .B2(new_n805), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1257), .C1(new_n812), .C2(new_n1157), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G132), .B2(new_n809), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1250), .A2(new_n1252), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n783), .B1(G68), .B2(new_n867), .C1(new_n1260), .C2(new_n866), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n955), .B2(new_n791), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1129), .B2(new_n1000), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1246), .A2(new_n1263), .ZN(G381));
  AND2_X1   g1064(.A1(new_n1214), .A2(new_n1243), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT122), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1042), .A2(new_n1267), .A3(new_n1263), .A4(new_n1246), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1266), .A2(new_n1268), .A3(G378), .ZN(G407));
  NAND2_X1  g1069(.A1(new_n708), .A2(G213), .ZN(new_n1270));
  OR3_X1    g1070(.A1(new_n1266), .A2(G378), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(new_n1271), .A3(G213), .ZN(G409));
  OAI211_X1 g1072(.A(KEYINPUT123), .B(new_n886), .C1(new_n861), .C2(new_n864), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1273), .A2(new_n1263), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1118), .A2(new_n1129), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1176), .B(KEYINPUT60), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n727), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT123), .B1(new_n865), .B2(new_n886), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1280), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1274), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1283));
  INV_X1    g1083(.A(G2897), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1270), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1281), .A2(new_n1288), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1270), .B1(KEYINPUT124), .B2(new_n1284), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(KEYINPUT124), .B2(new_n1284), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1214), .A2(G378), .A3(new_n1243), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1243), .B1(new_n1211), .B2(new_n981), .ZN(new_n1298));
  INV_X1    g1098(.A(G378), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1270), .ZN(new_n1302));
  AOI21_X1  g1102(.A(KEYINPUT61), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1291), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1304), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1042), .A2(G390), .ZN(new_n1307));
  XOR2_X1   g1107(.A(G393), .B(G396), .Z(new_n1308));
  INV_X1    g1108(.A(G390), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1016), .B2(new_n1041), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1270), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1297), .B2(new_n1300), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1303), .A2(new_n1306), .A3(new_n1313), .A4(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1315), .A2(new_n1318), .A3(new_n1291), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1315), .B2(new_n1295), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1315), .B2(new_n1291), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1323), .B2(new_n1313), .ZN(G405));
  NOR3_X1   g1124(.A1(new_n1305), .A2(KEYINPUT126), .A3(KEYINPUT127), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1326), .B1(new_n1291), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G375), .A2(new_n1299), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1297), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1330), .B(new_n1297), .C1(new_n1325), .C2(new_n1328), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1334), .B(new_n1313), .ZN(G402));
endmodule


