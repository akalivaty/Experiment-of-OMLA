//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G325));
  XOR2_X1   g032(.A(G325), .B(KEYINPUT68), .Z(G261));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n455), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  AND2_X1   g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n466), .A2(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n463), .A2(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT72), .Z(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT73), .ZN(G162));
  NAND3_X1  g059(.A1(new_n463), .A2(G138), .A3(new_n470), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n463), .A2(G126), .A3(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G164));
  AND2_X1   g068(.A1(KEYINPUT74), .A2(G651), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT74), .A2(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G62), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  XNOR2_X1  g076(.A(new_n501), .B(KEYINPUT78), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT74), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT74), .A2(G651), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT6), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n494), .A2(new_n495), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT75), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(G88), .A3(new_n499), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n508), .B2(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT74), .B(G651), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n516), .B2(new_n508), .ZN(new_n517));
  AOI211_X1 g092(.A(KEYINPUT76), .B(new_n514), .C1(new_n517), .C2(new_n507), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n519));
  INV_X1    g094(.A(new_n514), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n519), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n513), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT77), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n524), .B(new_n513), .C1(new_n518), .C2(new_n521), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n503), .B1(new_n523), .B2(new_n525), .ZN(G166));
  INV_X1    g101(.A(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n517), .B2(new_n507), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT7), .ZN(new_n532));
  AND2_X1   g107(.A1(G63), .A2(G651), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(new_n532), .B1(new_n499), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n499), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n517), .B2(new_n507), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n537), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n528), .A2(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n496), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n537), .A2(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n512), .A2(G43), .A3(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n536), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(new_n516), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n497), .B2(new_n498), .ZN(new_n562));
  AND2_X1   g137(.A1(G78), .A2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n510), .B1(new_n564), .B2(KEYINPUT80), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n566), .B1(new_n562), .B2(new_n563), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n567), .B1(new_n537), .B2(G91), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n528), .A2(new_n569), .A3(G53), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n569), .B1(new_n528), .B2(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(G299));
  INV_X1    g148(.A(new_n503), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n512), .A2(new_n520), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n512), .A2(new_n519), .A3(new_n520), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n524), .B1(new_n578), .B2(new_n513), .ZN(new_n579));
  INV_X1    g154(.A(new_n525), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(G303));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n510), .B1(new_n536), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(G49), .A2(G543), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n511), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n585));
  INV_X1    g160(.A(new_n507), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n512), .A2(new_n589), .A3(new_n584), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n583), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n512), .A2(G87), .A3(new_n499), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n537), .A2(KEYINPUT81), .A3(G87), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G61), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n536), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n528), .A2(G48), .B1(new_n516), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n537), .A2(G86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G305));
  AOI22_X1  g178(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(new_n496), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n512), .A2(G85), .A3(new_n499), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n512), .A2(G47), .A3(G543), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n536), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n528), .A2(G54), .B1(G651), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(KEYINPUT10), .B1(new_n537), .B2(G92), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n615), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n621), .B(new_n615), .C1(new_n617), .C2(new_n618), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n611), .B1(new_n623), .B2(new_n610), .ZN(G284));
  AOI21_X1  g199(.A(new_n611), .B1(new_n623), .B2(new_n610), .ZN(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n610), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n610), .ZN(G280));
  XNOR2_X1  g202(.A(G280), .B(KEYINPUT84), .ZN(G297));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(new_n629), .B2(G860), .ZN(G148));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n463), .A2(new_n471), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n475), .A2(G123), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  INV_X1    g216(.A(G111), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(G2105), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(G135), .B2(new_n469), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(G2100), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(G2096), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n639), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT85), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(new_n665), .A3(G14), .ZN(G401));
  XOR2_X1   g241(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  INV_X1    g249(.A(new_n667), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1971), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n687), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT87), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G35), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT94), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G162), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT29), .Z(new_n702));
  INV_X1    g277(.A(G2090), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G20), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT23), .Z(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G299), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1956), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n702), .B2(new_n703), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT96), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(new_n711), .C1(new_n702), .C2(new_n703), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n707), .A2(G21), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G286), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  NOR2_X1   g296(.A1(G27), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G164), .B2(G29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2078), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n698), .A2(G33), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n463), .A2(G127), .ZN(new_n726));
  AND2_X1   g301(.A1(G115), .A2(G2104), .ZN(new_n727));
  OAI21_X1  g302(.A(G2105), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n729));
  NAND2_X1  g304(.A1(G103), .A2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n470), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n469), .A2(G139), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n725), .B1(new_n734), .B2(new_n698), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G2072), .Z(new_n736));
  OR2_X1    g311(.A1(KEYINPUT30), .A2(G28), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT30), .A2(G28), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT31), .B(G11), .Z(new_n740));
  AOI211_X1 g315(.A(new_n739), .B(new_n740), .C1(new_n645), .C2(G29), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n698), .B1(new_n742), .B2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G160), .B2(G29), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n736), .B(new_n741), .C1(G2084), .C2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G1961), .ZN(new_n747));
  NAND2_X1  g322(.A1(G171), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G5), .B2(G16), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n724), .B(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n554), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G16), .B2(G19), .ZN(new_n752));
  INV_X1    g327(.A(G1341), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n749), .A2(new_n747), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n718), .A2(new_n719), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n752), .A2(new_n753), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n754), .A2(new_n755), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n698), .A2(G32), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n475), .A2(G129), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n471), .A2(G105), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(G141), .C2(new_n469), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n698), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT27), .B(G1996), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n745), .A2(G2084), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT92), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n698), .A2(G26), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n475), .A2(G128), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(G116), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G140), .B2(new_n469), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(G29), .ZN(new_n781));
  INV_X1    g356(.A(G2067), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n769), .A2(new_n771), .A3(new_n783), .ZN(new_n784));
  AND4_X1   g359(.A1(new_n721), .A2(new_n750), .A3(new_n758), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G4), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n623), .B2(G16), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT90), .B(G1348), .Z(new_n788));
  XOR2_X1   g363(.A(new_n787), .B(new_n788), .Z(new_n789));
  NAND4_X1  g364(.A1(new_n706), .A2(new_n716), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G22), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G166), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1971), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G16), .A2(G23), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT89), .Z(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G288), .B2(new_n707), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT33), .B(G1976), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n528), .A2(G48), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n600), .A2(new_n516), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n602), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G6), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n805), .A2(G1981), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(G1981), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n794), .B(new_n799), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  NOR2_X1   g385(.A1(G25), .A2(G29), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n475), .A2(G119), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G131), .B2(new_n469), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n811), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT88), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n608), .A2(G16), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G16), .B2(G24), .ZN(new_n824));
  INV_X1    g399(.A(G1986), .ZN(new_n825));
  AND2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n824), .A2(new_n825), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n809), .A2(new_n810), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT36), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT36), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n809), .A2(new_n831), .A3(new_n810), .A4(new_n828), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n790), .B1(new_n830), .B2(new_n832), .ZN(G311));
  NAND2_X1  g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n790), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  NAND2_X1  g411(.A1(new_n623), .A2(G559), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT38), .Z(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT97), .B(G93), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n512), .A2(new_n499), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n512), .A2(G55), .A3(G543), .ZN(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n536), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(new_n516), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n553), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n553), .A2(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n838), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  XNOR2_X1  g431(.A(new_n765), .B(new_n492), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n780), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n734), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT99), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n780), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n857), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n475), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n470), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n469), .B2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n636), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n818), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(KEYINPUT101), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n867), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n867), .A2(new_n876), .ZN(new_n878));
  XNOR2_X1  g453(.A(G162), .B(G160), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n881), .A2(new_n645), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n645), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n877), .B(new_n878), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n881), .A2(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n646), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n645), .A3(new_n882), .ZN(new_n888));
  INV_X1    g463(.A(new_n875), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n867), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n866), .A2(new_n862), .A3(new_n875), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n888), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n885), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g470(.A(new_n849), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n623), .B2(new_n629), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n629), .A3(new_n623), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(G651), .A3(new_n567), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n537), .A2(G91), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n528), .A2(G53), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT9), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(new_n570), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n619), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n528), .A2(G54), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n614), .A2(G651), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n537), .A2(G92), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT10), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(new_n616), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(G299), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n907), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n898), .A2(new_n899), .A3(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT41), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n907), .B2(new_n915), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n899), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n897), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n591), .A2(new_n596), .A3(new_n608), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n608), .B1(new_n591), .B2(new_n596), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n523), .A2(new_n525), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n802), .B1(new_n931), .B2(new_n574), .ZN(new_n932));
  AOI211_X1 g507(.A(new_n503), .B(G305), .C1(new_n523), .C2(new_n525), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n927), .B(new_n930), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G303), .A2(G305), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n928), .B2(new_n929), .ZN(new_n936));
  NAND2_X1  g511(.A1(G288), .A2(G290), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n591), .A2(new_n596), .A3(new_n608), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n927), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n574), .A3(new_n802), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(new_n936), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT103), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n926), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n925), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT103), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT103), .B1(new_n934), .B2(new_n941), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n947), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n924), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n610), .B1(new_n948), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n846), .A2(new_n610), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n954), .A2(KEYINPUT104), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n951), .A2(new_n924), .A3(new_n952), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(G868), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n961), .B2(new_n955), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n957), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n955), .ZN(G331));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n548), .A2(new_n552), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n528), .A2(G55), .B1(new_n516), .B2(new_n844), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n547), .A4(new_n840), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n553), .A2(new_n846), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(G301), .ZN(new_n970));
  AOI21_X1  g545(.A(G301), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n970), .A2(new_n971), .A3(G286), .ZN(new_n972));
  OAI21_X1  g547(.A(G171), .B1(new_n847), .B2(new_n848), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n969), .A3(G301), .ZN(new_n974));
  AOI21_X1  g549(.A(G168), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n916), .B(new_n965), .C1(new_n972), .C2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(G286), .B1(new_n970), .B2(new_n971), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(G168), .A3(new_n974), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(new_n978), .C1(new_n919), .C2(new_n920), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n978), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n965), .B1(new_n981), .B2(new_n916), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n949), .A2(new_n950), .ZN(new_n984));
  AOI21_X1  g559(.A(G37), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n916), .B1(new_n972), .B2(new_n975), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n979), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(KEYINPUT106), .C1(new_n949), .C2(new_n950), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n949), .B2(new_n950), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AND4_X1   g566(.A1(KEYINPUT43), .A2(new_n985), .A3(new_n988), .A4(new_n991), .ZN(new_n992));
  OAI22_X1  g567(.A1(new_n980), .A2(new_n982), .B1(new_n949), .B2(new_n950), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT43), .B1(new_n985), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n976), .A2(new_n979), .ZN(new_n996));
  INV_X1    g571(.A(new_n982), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n945), .A3(new_n997), .A4(new_n944), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(new_n893), .A3(new_n993), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n985), .A2(new_n1001), .A3(new_n988), .A4(new_n991), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n995), .A2(new_n1005), .ZN(G397));
  INV_X1    g581(.A(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n492), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n466), .A2(G40), .A3(new_n472), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n817), .B(new_n820), .ZN(new_n1013));
  XOR2_X1   g588(.A(new_n1013), .B(KEYINPUT108), .Z(new_n1014));
  XNOR2_X1  g589(.A(new_n780), .B(new_n782), .ZN(new_n1015));
  INV_X1    g590(.A(G1996), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n765), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n608), .A2(new_n825), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT107), .Z(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n825), .B2(new_n608), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1012), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n492), .A2(new_n1026), .A3(new_n1007), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT114), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n492), .A2(new_n1029), .A3(new_n1026), .A4(new_n1007), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT109), .B(G2090), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1011), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1011), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1010), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n793), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  OAI211_X1 g615(.A(G303), .B(G8), .C1(KEYINPUT111), .C2(KEYINPUT55), .ZN(new_n1041));
  INV_X1    g616(.A(G8), .ZN(new_n1042));
  AND2_X1   g617(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1043));
  NOR2_X1   g618(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1044));
  OAI22_X1  g619(.A1(G166), .A2(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1027), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1026), .B1(new_n492), .B2(new_n1007), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1011), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1051), .A2(new_n1032), .B1(new_n1037), .B2(new_n793), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1032), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1038), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT110), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1045), .ZN(new_n1059));
  NOR3_X1   g634(.A1(G166), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1054), .B(new_n1058), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n591), .A2(new_n596), .A3(G1976), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT112), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1042), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1062), .B2(KEYINPUT112), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n601), .A2(new_n1069), .A3(new_n602), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n601), .B2(new_n602), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT113), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT49), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT113), .B(new_n1074), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1066), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1062), .A2(KEYINPUT112), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(new_n1063), .A3(new_n1066), .A4(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1068), .A2(new_n1076), .A3(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT115), .A4(new_n1045), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1048), .A2(new_n1061), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1065), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1051), .A2(G1348), .B1(G2067), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1085), .A2(new_n623), .A3(KEYINPUT60), .ZN(new_n1086));
  INV_X1    g661(.A(new_n622), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n913), .A2(new_n616), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n621), .B1(new_n1088), .B2(new_n615), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G1348), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n1056), .A2(new_n1091), .B1(new_n1065), .B2(new_n782), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n623), .A2(KEYINPUT60), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n571), .B2(new_n572), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n905), .A2(KEYINPUT119), .A3(new_n570), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n568), .A3(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n906), .A2(KEYINPUT57), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  XOR2_X1   g678(.A(KEYINPUT117), .B(G1956), .Z(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1011), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1106));
  XNOR2_X1  g681(.A(KEYINPUT56), .B(G2072), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1106), .A2(new_n1035), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1094), .A2(new_n1095), .B1(new_n1110), .B2(KEYINPUT61), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1010), .A2(new_n1036), .A3(new_n1016), .A4(new_n1035), .ZN(new_n1116));
  XOR2_X1   g691(.A(KEYINPUT58), .B(G1341), .Z(new_n1117));
  AOI22_X1  g692(.A1(new_n1116), .A2(KEYINPUT121), .B1(new_n1084), .B2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1010), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1016), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT59), .B1(new_n1122), .B2(new_n554), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  AOI211_X1 g699(.A(new_n1124), .B(new_n553), .C1(new_n1118), .C2(new_n1121), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1111), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1109), .B1(new_n1128), .B2(new_n1103), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1101), .A2(KEYINPUT120), .A3(new_n1102), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1085), .A2(new_n623), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1129), .A2(new_n1130), .B1(new_n1110), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT124), .B1(G168), .B2(new_n1042), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n1135));
  NAND3_X1  g710(.A1(G286), .A2(new_n1135), .A3(G8), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT116), .B(G2084), .Z(new_n1140));
  AND3_X1   g715(.A1(new_n1033), .A2(new_n1027), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1966), .B1(new_n1106), .B2(new_n1035), .ZN(new_n1142));
  OAI21_X1  g717(.A(G8), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1033), .A2(new_n1027), .A3(new_n1140), .ZN(new_n1147));
  OAI211_X1 g722(.A(KEYINPUT123), .B(new_n1147), .C1(new_n1119), .C2(G1966), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n1148), .A3(G8), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1149), .A2(new_n1138), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1137), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT125), .B(KEYINPUT51), .Z(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1144), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1037), .A2(G2078), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1155), .A2(new_n1156), .B1(new_n747), .B2(new_n1056), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(KEYINPUT126), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1037), .A2(G2078), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(KEYINPUT53), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G301), .B(KEYINPUT54), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n1159), .B2(KEYINPUT53), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1157), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1154), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1133), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1154), .A2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(KEYINPUT62), .B(new_n1144), .C1(new_n1150), .C2(new_n1153), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1162), .A2(G171), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1083), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n1143), .A2(G286), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1083), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(new_n1045), .A3(new_n1041), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1177), .A2(new_n1176), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1061), .A4(new_n1081), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1076), .A2(new_n1078), .A3(new_n596), .A4(new_n591), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(G1981), .B2(G305), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1061), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1066), .A2(new_n1185), .B1(new_n1186), .B2(new_n1081), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1025), .B1(new_n1175), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1022), .A2(new_n1012), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1020), .A2(new_n1012), .B1(KEYINPUT48), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(KEYINPUT48), .B2(new_n1191), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1012), .A2(new_n1016), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT46), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT127), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1015), .A2(new_n766), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1198), .A2(new_n1012), .B1(new_n1195), .B2(new_n1194), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT47), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n818), .A2(new_n820), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1018), .A2(new_n1202), .B1(G2067), .B2(new_n780), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1012), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1193), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1189), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G319), .ZN(new_n1208));
  NOR4_X1   g782(.A1(G229), .A2(new_n1208), .A3(G401), .A4(G227), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n1003), .A2(new_n1209), .A3(new_n894), .ZN(G225));
  INV_X1    g784(.A(G225), .ZN(G308));
endmodule


