

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(n434), .B(KEYINPUT55), .ZN(n435) );
  XNOR2_X1 U326 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U327 ( .A(n411), .B(KEYINPUT54), .ZN(n412) );
  XNOR2_X1 U328 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U329 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U330 ( .A(n436), .B(n435), .ZN(n454) );
  XNOR2_X1 U331 ( .A(n363), .B(n362), .ZN(n563) );
  XNOR2_X1 U332 ( .A(n456), .B(G176GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  XOR2_X1 U334 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n294) );
  XNOR2_X1 U335 ( .A(KEYINPUT5), .B(KEYINPUT6), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n311) );
  XOR2_X1 U337 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n296) );
  XNOR2_X1 U338 ( .A(KEYINPUT91), .B(KEYINPUT88), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U340 ( .A(n297), .B(G57GAT), .Z(n299) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G148GAT), .Z(n314) );
  XNOR2_X1 U342 ( .A(n314), .B(G85GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n304) );
  XOR2_X1 U344 ( .A(G113GAT), .B(KEYINPUT0), .Z(n442) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(G127GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n300), .B(G155GAT), .ZN(n341) );
  XOR2_X1 U347 ( .A(n442), .B(n341), .Z(n302) );
  NAND2_X1 U348 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U350 ( .A(n304), .B(n303), .Z(n309) );
  XOR2_X1 U351 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n306) );
  XNOR2_X1 U352 ( .A(G141GAT), .B(G162GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n425) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(KEYINPUT77), .ZN(n352) );
  XNOR2_X1 U356 ( .A(n425), .B(n352), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U358 ( .A(n311), .B(n310), .Z(n466) );
  XOR2_X1 U359 ( .A(KEYINPUT92), .B(n466), .Z(n522) );
  INV_X1 U360 ( .A(n522), .ZN(n504) );
  XOR2_X1 U361 ( .A(KEYINPUT13), .B(KEYINPUT69), .Z(n313) );
  XNOR2_X1 U362 ( .A(G71GAT), .B(G57GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n333) );
  XOR2_X1 U364 ( .A(n314), .B(n333), .Z(n316) );
  NAND2_X1 U365 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n330) );
  XOR2_X1 U367 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n318) );
  XNOR2_X1 U368 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n320) );
  XNOR2_X1 U371 ( .A(G78GAT), .B(KEYINPUT73), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U373 ( .A(n322), .B(n321), .Z(n328) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n404) );
  XOR2_X1 U377 ( .A(KEYINPUT71), .B(G85GAT), .Z(n326) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n361) );
  XNOR2_X1 U380 ( .A(n404), .B(n361), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U382 ( .A(n330), .B(n329), .Z(n575) );
  INV_X1 U383 ( .A(KEYINPUT45), .ZN(n366) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n332) );
  XNOR2_X1 U385 ( .A(G15GAT), .B(G64GAT), .ZN(n331) );
  XOR2_X1 U386 ( .A(n332), .B(n331), .Z(n345) );
  XOR2_X1 U387 ( .A(G22GAT), .B(G78GAT), .Z(n418) );
  XOR2_X1 U388 ( .A(n333), .B(n418), .Z(n335) );
  NAND2_X1 U389 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U391 ( .A(KEYINPUT80), .B(KEYINPUT15), .Z(n337) );
  XNOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT81), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U394 ( .A(n339), .B(n338), .Z(n343) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n340), .B(G211GAT), .ZN(n400) );
  XNOR2_X1 U397 ( .A(n341), .B(n400), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U399 ( .A(n345), .B(n344), .ZN(n580) );
  XNOR2_X1 U400 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n364) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n347) );
  XOR2_X1 U402 ( .A(G50GAT), .B(G218GAT), .Z(n421) );
  XOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  XNOR2_X1 U404 ( .A(n421), .B(n399), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(n348), .B(KEYINPUT9), .Z(n355) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  INV_X1 U408 ( .A(KEYINPUT10), .ZN(n349) );
  XNOR2_X1 U409 ( .A(G162GAT), .B(n353), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT64), .B(KEYINPUT75), .Z(n357) );
  XNOR2_X1 U412 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n358) );
  XNOR2_X1 U414 ( .A(n359), .B(n358), .ZN(n363) );
  XNOR2_X1 U415 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n360), .B(KEYINPUT7), .ZN(n373) );
  XOR2_X1 U417 ( .A(n373), .B(n361), .Z(n362) );
  XNOR2_X1 U418 ( .A(n364), .B(n563), .ZN(n486) );
  NOR2_X1 U419 ( .A1(n580), .A2(n486), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  NOR2_X1 U421 ( .A1(n575), .A2(n367), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n368), .B(KEYINPUT112), .ZN(n387) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n370) );
  XNOR2_X1 U424 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n376) );
  XOR2_X1 U427 ( .A(G1GAT), .B(G113GAT), .Z(n372) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G15GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n378), .B(n377), .ZN(n386) );
  NAND2_X1 U433 ( .A1(G229GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X1 U434 ( .A(G141GAT), .B(G197GAT), .Z(n380) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(G22GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n382) );
  XOR2_X1 U437 ( .A(G29GAT), .B(G50GAT), .Z(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n501) );
  INV_X1 U441 ( .A(n501), .ZN(n570) );
  NAND2_X1 U442 ( .A1(n387), .A2(n570), .ZN(n394) );
  XOR2_X1 U443 ( .A(KEYINPUT110), .B(n580), .Z(n560) );
  XNOR2_X1 U444 ( .A(n575), .B(KEYINPUT41), .ZN(n548) );
  NOR2_X1 U445 ( .A1(n570), .A2(n548), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n388), .B(KEYINPUT111), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  INV_X1 U448 ( .A(n563), .ZN(n555) );
  NAND2_X1 U449 ( .A1(n390), .A2(n555), .ZN(n391) );
  NOR2_X1 U450 ( .A1(n560), .A2(n391), .ZN(n392) );
  XNOR2_X1 U451 ( .A(KEYINPUT47), .B(n392), .ZN(n393) );
  NAND2_X1 U452 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n395), .B(KEYINPUT48), .ZN(n531) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n397) );
  XNOR2_X1 U455 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U457 ( .A(G169GAT), .B(n398), .Z(n449) );
  XOR2_X1 U458 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n403), .B(KEYINPUT94), .Z(n406) );
  XNOR2_X1 U462 ( .A(n404), .B(KEYINPUT95), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U464 ( .A(n407), .B(KEYINPUT93), .Z(n409) );
  XOR2_X1 U465 ( .A(G197GAT), .B(KEYINPUT21), .Z(n417) );
  XNOR2_X1 U466 ( .A(G218GAT), .B(n417), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U468 ( .A(n449), .B(n410), .Z(n524) );
  INV_X1 U469 ( .A(n524), .ZN(n508) );
  NAND2_X1 U470 ( .A1(n531), .A2(n508), .ZN(n413) );
  XOR2_X1 U471 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n411) );
  NOR2_X1 U472 ( .A1(n504), .A2(n414), .ZN(n567) );
  XOR2_X1 U473 ( .A(KEYINPUT87), .B(KEYINPUT85), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n433) );
  XOR2_X1 U476 ( .A(G211GAT), .B(G106GAT), .Z(n420) );
  XNOR2_X1 U477 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n431) );
  XOR2_X1 U480 ( .A(G204GAT), .B(G148GAT), .Z(n424) );
  XNOR2_X1 U481 ( .A(KEYINPUT86), .B(KEYINPUT23), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U483 ( .A(G155GAT), .B(n425), .Z(n427) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n468) );
  NAND2_X1 U489 ( .A1(n567), .A2(n468), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n434) );
  XOR2_X1 U491 ( .A(KEYINPUT82), .B(G183GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(G71GAT), .B(G176GAT), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n453) );
  XOR2_X1 U494 ( .A(G99GAT), .B(G190GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(G134GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U497 ( .A(n441), .B(G120GAT), .Z(n444) );
  XNOR2_X1 U498 ( .A(G15GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U500 ( .A(KEYINPUT83), .B(G127GAT), .Z(n446) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U503 ( .A(n448), .B(n447), .Z(n451) );
  XNOR2_X1 U504 ( .A(n449), .B(KEYINPUT20), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U506 ( .A(n453), .B(n452), .Z(n532) );
  INV_X1 U507 ( .A(n532), .ZN(n512) );
  NAND2_X1 U508 ( .A1(n454), .A2(n512), .ZN(n455) );
  XOR2_X1 U509 ( .A(n455), .B(KEYINPUT120), .Z(n564) );
  INV_X1 U510 ( .A(n564), .ZN(n557) );
  NOR2_X1 U511 ( .A1(n557), .A2(n548), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n575), .A2(n570), .ZN(n490) );
  NAND2_X1 U514 ( .A1(n512), .A2(n508), .ZN(n459) );
  NAND2_X1 U515 ( .A1(n468), .A2(n459), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n460), .B(KEYINPUT25), .ZN(n464) );
  XNOR2_X1 U517 ( .A(KEYINPUT27), .B(n524), .ZN(n469) );
  NOR2_X1 U518 ( .A1(n512), .A2(n468), .ZN(n462) );
  XNOR2_X1 U519 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n461) );
  XOR2_X1 U520 ( .A(n462), .B(n461), .Z(n568) );
  NOR2_X1 U521 ( .A1(n469), .A2(n568), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n472) );
  XOR2_X1 U524 ( .A(KEYINPUT28), .B(KEYINPUT65), .Z(n467) );
  XOR2_X1 U525 ( .A(n468), .B(n467), .Z(n515) );
  INV_X1 U526 ( .A(n515), .ZN(n535) );
  NOR2_X1 U527 ( .A1(n522), .A2(n469), .ZN(n530) );
  NAND2_X1 U528 ( .A1(n535), .A2(n530), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n470), .A2(n512), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n487) );
  NOR2_X1 U531 ( .A1(n580), .A2(n563), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U533 ( .A1(n487), .A2(n474), .ZN(n502) );
  NAND2_X1 U534 ( .A1(n490), .A2(n502), .ZN(n483) );
  NOR2_X1 U535 ( .A1(n522), .A2(n483), .ZN(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U537 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U539 ( .A1(n524), .A2(n483), .ZN(n479) );
  XNOR2_X1 U540 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n478) );
  XNOR2_X1 U541 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n532), .A2(n483), .ZN(n482) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n535), .A2(n483), .ZN(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT100), .B(n484), .Z(n485) );
  XNOR2_X1 U548 ( .A(G22GAT), .B(n485), .ZN(G1327GAT) );
  XOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .Z(n493) );
  NOR2_X1 U550 ( .A1(n486), .A2(n487), .ZN(n488) );
  NAND2_X1 U551 ( .A1(n580), .A2(n488), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT37), .B(n489), .ZN(n521) );
  NAND2_X1 U553 ( .A1(n490), .A2(n521), .ZN(n491) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(n491), .Z(n499) );
  NAND2_X1 U555 ( .A1(n499), .A2(n504), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n508), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT102), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G36GAT), .B(n495), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n497) );
  NAND2_X1 U561 ( .A1(n499), .A2(n512), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n515), .A2(n499), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n506) );
  NOR2_X1 U567 ( .A1(n501), .A2(n548), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n520), .A2(n502), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(n503), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n516), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U572 ( .A(G57GAT), .B(n507), .Z(G1332GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U574 ( .A1(n516), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n511), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n516), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT108), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  NAND2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U585 ( .A1(n522), .A2(n527), .ZN(n523) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n524), .A2(n527), .ZN(n525) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n525), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n532), .A2(n527), .ZN(n526) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U591 ( .A1(n535), .A2(n527), .ZN(n528) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(n528), .Z(n529) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n546) );
  NOR2_X1 U595 ( .A1(n532), .A2(n546), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT113), .B(n533), .Z(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n539) );
  NOR2_X1 U598 ( .A1(n570), .A2(n539), .ZN(n536) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n548), .A2(n539), .ZN(n538) );
  XNOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  INV_X1 U603 ( .A(n539), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n542), .A2(n560), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n563), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  OR2_X1 U611 ( .A1(n546), .A2(n568), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n570), .A2(n554), .ZN(n547) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U614 ( .A1(n554), .A2(n548), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT115), .Z(n550) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n580), .A2(n554), .ZN(n553) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n556), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n570), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n564), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(n562), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  INV_X1 U632 ( .A(n567), .ZN(n569) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n576) );
  INV_X1 U634 ( .A(n576), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n570), .A2(n584), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n582) );
  OR2_X1 U645 ( .A1(n584), .A2(n580), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n486), .A2(n584), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

