//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT75), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n192), .A2(KEYINPUT75), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n190), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(KEYINPUT16), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n187), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(KEYINPUT75), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n189), .B2(KEYINPUT75), .ZN(new_n199));
  OAI211_X1 g013(.A(G146), .B(new_n197), .C1(new_n199), .C2(new_n188), .ZN(new_n200));
  NOR2_X1   g014(.A1(G237), .A2(G953), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G214), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT89), .A3(G143), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT89), .A2(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT89), .A2(G143), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n204), .A2(G214), .A3(new_n201), .A4(new_n205), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT17), .A4(G131), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(new_n200), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n206), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n211), .B(G131), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n196), .A2(KEYINPUT90), .A3(new_n200), .A4(new_n207), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G113), .B(G122), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n189), .A2(new_n187), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n199), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n187), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT18), .A4(G131), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n211), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n224), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n216), .A2(new_n219), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n211), .B(new_n227), .ZN(new_n231));
  MUX2_X1   g045(.A(new_n189), .B(new_n199), .S(KEYINPUT19), .Z(new_n232));
  OAI211_X1 g046(.A(new_n231), .B(new_n200), .C1(new_n232), .C2(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n219), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(G475), .A2(G902), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n241));
  INV_X1    g055(.A(new_n238), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n242), .B1(new_n230), .B2(new_n236), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT92), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT20), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n237), .B(new_n247), .C1(new_n246), .C2(new_n242), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n230), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n219), .B1(new_n216), .B2(new_n229), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G475), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G478), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT15), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT78), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G107), .ZN(new_n260));
  INV_X1    g074(.A(G107), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT78), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XOR2_X1   g077(.A(G116), .B(G122), .Z(new_n264));
  OR2_X1    g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G116), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT14), .A3(G122), .ZN(new_n267));
  OAI211_X1 g081(.A(G107), .B(new_n267), .C1(new_n264), .C2(KEYINPUT14), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G128), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT93), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G143), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n272), .B1(new_n271), .B2(new_n274), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n265), .B(new_n268), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT95), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n275), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(KEYINPUT95), .A3(new_n265), .A4(new_n268), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n263), .B(new_n264), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n272), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n271), .A2(new_n274), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n271), .B2(new_n274), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT94), .B(new_n285), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT9), .B(G234), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G217), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(G953), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n294), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n298), .B1(new_n284), .B2(new_n294), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n250), .B(new_n258), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n284), .A2(new_n294), .ZN(new_n304));
  INV_X1    g118(.A(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n299), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n258), .B1(new_n307), .B2(new_n250), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n255), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  INV_X1    g125(.A(G137), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n311), .B1(new_n312), .B2(G134), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n272), .A2(KEYINPUT66), .A3(G137), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT11), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(new_n272), .B2(G137), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(KEYINPUT11), .A3(G134), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G131), .B1(new_n315), .B2(new_n319), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n312), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT11), .B1(new_n312), .B2(G134), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n313), .A2(new_n314), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n227), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n327), .B(G104), .C1(new_n260), .C2(new_n262), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n261), .A2(G104), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n261), .A2(G104), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(KEYINPUT3), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n261), .A2(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n259), .A2(G107), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n334), .A2(new_n335), .A3(new_n218), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n218), .B2(G107), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n261), .A2(KEYINPUT79), .A3(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G101), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n273), .A2(KEYINPUT1), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n187), .A2(G143), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n269), .A2(G146), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n269), .A2(KEYINPUT1), .A3(G146), .ZN(new_n346));
  XNOR2_X1  g160(.A(G143), .B(G146), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n345), .B(new_n346), .C1(G128), .C2(new_n347), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n333), .A2(new_n341), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n333), .B2(new_n341), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT81), .B(new_n326), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n326), .C1(new_n349), .C2(new_n350), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT12), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT3), .B(new_n218), .C1(new_n334), .C2(new_n335), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(G104), .B2(new_n261), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT0), .A2(G128), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT64), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(KEYINPUT0), .A3(G128), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n343), .A2(new_n344), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT0), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n273), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n343), .A2(new_n344), .B1(new_n370), .B2(new_n273), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT65), .A3(new_n368), .ZN(new_n376));
  INV_X1    g190(.A(new_n364), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n374), .A2(new_n376), .B1(new_n347), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G101), .C1(new_n359), .C2(new_n361), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n363), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AND4_X1   g195(.A1(new_n227), .A2(new_n324), .A3(new_n317), .A4(new_n318), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n227), .B1(new_n323), .B2(new_n324), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n349), .A2(KEYINPUT10), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n333), .A2(new_n341), .A3(new_n348), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT10), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n358), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G140), .ZN(new_n394));
  INV_X1    g208(.A(G953), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(G227), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n394), .B(new_n396), .Z(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n381), .A2(new_n385), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(KEYINPUT80), .A3(new_n384), .A4(new_n388), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n389), .A2(new_n390), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n381), .A2(new_n388), .A3(new_n385), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n403), .A2(new_n326), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n393), .A2(new_n398), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G469), .B1(new_n406), .B2(G902), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n404), .B1(new_n400), .B2(new_n401), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n397), .B1(new_n391), .B2(new_n392), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n353), .A2(new_n355), .A3(new_n357), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n397), .A2(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(KEYINPUT83), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n411), .A2(new_n250), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n266), .A2(G119), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT67), .B(G119), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n421), .B2(new_n266), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT2), .B(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n425), .B(new_n420), .C1(new_n266), .C2(new_n421), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n363), .A2(new_n427), .A3(new_n380), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT5), .B(new_n420), .C1(new_n421), .C2(new_n266), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT5), .ZN(new_n430));
  INV_X1    g244(.A(G119), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n431), .A2(KEYINPUT67), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(KEYINPUT67), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(G116), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(G113), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n435), .A2(new_n426), .A3(new_n333), .A4(new_n341), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(KEYINPUT8), .ZN(new_n439));
  INV_X1    g253(.A(new_n436), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n435), .A2(new_n426), .B1(new_n333), .B2(new_n341), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n348), .A2(G125), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n347), .A2(new_n377), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n375), .A2(KEYINPUT65), .A3(new_n368), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT65), .B1(new_n375), .B2(new_n368), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n444), .B1(new_n451), .B2(G125), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n447), .B1(new_n452), .B2(new_n446), .ZN(new_n453));
  INV_X1    g267(.A(G224), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(new_n454), .B2(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n447), .B(new_n455), .C1(new_n452), .C2(new_n446), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n443), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n419), .B1(new_n459), .B2(G902), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n438), .A2(new_n442), .ZN(new_n461));
  INV_X1    g275(.A(G125), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n445), .B1(new_n378), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT86), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n455), .B1(new_n464), .B2(new_n447), .ZN(new_n465));
  INV_X1    g279(.A(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT87), .A3(new_n250), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n428), .A2(new_n436), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n437), .B(KEYINPUT84), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(KEYINPUT85), .A2(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n436), .A4(new_n437), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n469), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n454), .A2(G953), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n453), .B(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n460), .A2(new_n468), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT88), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n482), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n460), .A2(new_n468), .A3(new_n479), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G234), .A2(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(G952), .A3(new_n395), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(G902), .A3(G953), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G214), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n486), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n310), .A2(new_n418), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n196), .A2(new_n200), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n421), .A2(new_n273), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(G119), .B2(new_n273), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT24), .B(G110), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n421), .A2(new_n273), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT73), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n421), .A2(new_n506), .A3(new_n273), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT23), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n505), .B(new_n507), .C1(new_n508), .C2(new_n499), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n273), .A2(KEYINPUT23), .A3(G119), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n503), .B1(new_n511), .B2(G110), .ZN(new_n512));
  INV_X1    g326(.A(G110), .ZN(new_n513));
  AOI211_X1 g327(.A(KEYINPUT74), .B(new_n513), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n498), .B(new_n502), .C1(new_n512), .C2(new_n514), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n511), .A2(G110), .B1(new_n500), .B2(new_n501), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n200), .A3(new_n222), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n395), .A2(G221), .A3(G234), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(G137), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT77), .B(KEYINPUT22), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n515), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n515), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n250), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT25), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n297), .B1(G234), .B2(new_n250), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n250), .C1(new_n522), .C2(new_n523), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n524), .A2(new_n526), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n201), .A2(G210), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT26), .B(G101), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n374), .A2(new_n376), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n326), .A3(new_n448), .ZN(new_n543));
  INV_X1    g357(.A(new_n427), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n272), .A2(G137), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n312), .A2(G134), .ZN(new_n546));
  OAI21_X1  g360(.A(G131), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n325), .A2(new_n348), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n544), .B1(new_n543), .B2(new_n548), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT28), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n541), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n548), .B1(new_n451), .B2(new_n384), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT30), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n559), .B(new_n548), .C1(new_n451), .C2(new_n384), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n550), .B1(new_n561), .B2(new_n427), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n556), .B1(new_n562), .B2(new_n541), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT70), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n555), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n560), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n559), .B1(new_n543), .B2(new_n548), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n427), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n568), .A2(new_n556), .A3(new_n549), .A4(new_n541), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n564), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n549), .A3(new_n541), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT31), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT71), .B(new_n534), .C1(new_n565), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n575));
  INV_X1    g389(.A(new_n555), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(new_n564), .A3(KEYINPUT31), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n578), .B2(new_n533), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n532), .B1(new_n574), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n534), .B1(new_n565), .B2(new_n573), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n552), .A2(new_n541), .A3(new_n554), .ZN(new_n582));
  INV_X1    g396(.A(new_n541), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n544), .B1(new_n558), .B2(new_n560), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n550), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT72), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n582), .A2(new_n586), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n582), .A2(new_n585), .A3(new_n590), .A4(new_n586), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n589), .A3(new_n250), .A4(new_n591), .ZN(new_n592));
  AOI22_X1  g406(.A1(KEYINPUT32), .A2(new_n581), .B1(new_n592), .B2(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n531), .B1(new_n580), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n497), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  INV_X1    g410(.A(KEYINPUT96), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n483), .A2(new_n597), .A3(new_n485), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n485), .A2(new_n597), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n598), .A2(new_n493), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n304), .B2(KEYINPUT97), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n299), .A3(new_n306), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n284), .B2(new_n294), .ZN(new_n605));
  OAI22_X1  g419(.A1(new_n300), .A2(new_n301), .B1(new_n605), .B2(new_n601), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n256), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n307), .A2(new_n256), .A3(new_n250), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n256), .A2(new_n250), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n249), .A2(new_n254), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n491), .A4(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n598), .A2(new_n599), .A3(new_n491), .A4(new_n493), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n613), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n531), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n578), .B2(new_n250), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n578), .A2(new_n533), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT71), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n581), .A2(new_n575), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n417), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n407), .B2(new_n415), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n619), .A2(new_n620), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  AND3_X1   g446(.A1(new_n243), .A2(KEYINPUT100), .A3(new_n244), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT100), .B1(new_n243), .B2(new_n244), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT91), .B1(new_n239), .B2(KEYINPUT20), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n243), .A2(new_n241), .A3(new_n244), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n240), .A2(KEYINPUT99), .A3(new_n245), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n303), .A2(new_n308), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n254), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n617), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n620), .A3(new_n629), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NAND2_X1  g462(.A1(new_n515), .A2(new_n517), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n250), .C1(new_n297), .C2(G234), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n529), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n497), .A2(new_n626), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  NAND2_X1  g470(.A1(new_n580), .A2(new_n593), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n493), .A2(new_n598), .A3(new_n653), .A4(new_n599), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n488), .B1(new_n490), .B2(G900), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n641), .A2(new_n643), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n658), .A3(new_n661), .A4(new_n628), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n418), .B1(new_n580), .B2(new_n593), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n661), .A4(new_n658), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G128), .ZN(G30));
  XOR2_X1   g482(.A(new_n659), .B(KEYINPUT39), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n418), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT104), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n653), .B1(new_n671), .B2(KEYINPUT40), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n623), .A2(new_n532), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n624), .A2(new_n625), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(new_n532), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n550), .A2(new_n551), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n541), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n562), .B2(new_n541), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n682), .B2(G902), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT102), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n486), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n309), .B1(new_n249), .B2(new_n254), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n494), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n672), .A2(new_n676), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G143), .ZN(G45));
  NOR2_X1   g507(.A1(new_n613), .A2(new_n660), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n657), .A2(new_n658), .A3(new_n628), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n664), .A2(KEYINPUT105), .A3(new_n658), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NAND2_X1  g514(.A1(new_n411), .A2(new_n250), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n417), .A3(new_n415), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n531), .B(new_n703), .C1(new_n580), .C2(new_n593), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n619), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n645), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND4_X1  g523(.A1(new_n598), .A2(new_n653), .A3(new_n599), .A4(new_n493), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n710), .A2(new_n492), .A3(new_n703), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n310), .B1(new_n580), .B2(new_n593), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  NAND2_X1  g528(.A1(new_n576), .A2(new_n572), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n569), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n715), .A2(KEYINPUT106), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n533), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n622), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n620), .A2(new_n719), .A3(new_n720), .A4(new_n491), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n688), .A2(new_n598), .A3(new_n493), .A4(new_n599), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n721), .A2(new_n722), .A3(new_n703), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(G122), .Z(G24));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n720), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n703), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n658), .A3(new_n694), .A4(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT107), .B(G125), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G27));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n416), .B2(new_n417), .ZN(new_n732));
  AOI211_X1 g546(.A(KEYINPUT108), .B(new_n627), .C1(new_n407), .C2(new_n415), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n483), .A2(new_n485), .A3(new_n493), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n613), .A2(new_n660), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n594), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n594), .A2(new_n734), .A3(KEYINPUT109), .A4(new_n736), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n743));
  INV_X1    g557(.A(new_n732), .ZN(new_n744));
  INV_X1    g558(.A(new_n733), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n736), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n581), .A2(KEYINPUT32), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n531), .B1(new_n748), .B2(new_n593), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n743), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n740), .B(new_n531), .C1(new_n593), .C2(new_n748), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(KEYINPUT110), .A3(new_n736), .A4(new_n734), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n742), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  INV_X1    g570(.A(new_n735), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n594), .A2(new_n734), .A3(new_n661), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n255), .A2(new_n611), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n255), .A2(KEYINPUT43), .A3(new_n611), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT112), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n653), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n626), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT44), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n406), .B2(KEYINPUT45), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n406), .A2(KEYINPUT45), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT111), .B(G469), .C1(new_n406), .C2(KEYINPUT45), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n627), .B1(new_n781), .B2(new_n415), .ZN(new_n782));
  INV_X1    g596(.A(new_n669), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n765), .A2(KEYINPUT44), .A3(new_n770), .A4(new_n767), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n757), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n771), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G137), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(G39));
  INV_X1    g603(.A(new_n736), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n657), .A2(new_n620), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  AOI21_X1  g610(.A(new_n418), .B1(new_n679), .B2(new_n683), .ZN(new_n797));
  INV_X1    g611(.A(new_n722), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n769), .A3(new_n659), .A4(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n667), .A2(new_n699), .A3(new_n728), .A4(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n666), .A2(new_n663), .B1(new_n697), .B2(new_n698), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT52), .A3(new_n728), .A4(new_n799), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n734), .A2(new_n614), .A3(new_n726), .ZN(new_n806));
  INV_X1    g620(.A(new_n641), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n664), .A2(new_n254), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n808), .B2(new_n642), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n653), .A3(new_n659), .A4(new_n757), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n755), .A2(new_n758), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n723), .B1(new_n619), .B2(new_n704), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n704), .A2(new_n645), .B1(new_n711), .B2(new_n712), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n813), .B1(new_n812), .B2(new_n814), .ZN(new_n816));
  INV_X1    g630(.A(new_n496), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT115), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n614), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n496), .B2(new_n613), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n629), .A2(new_n819), .A3(new_n820), .A4(new_n620), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n612), .A2(new_n309), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n629), .A2(new_n620), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n823), .A3(new_n595), .A4(new_n654), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n815), .A2(new_n816), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n805), .A2(new_n811), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT53), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n814), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n829));
  INV_X1    g643(.A(new_n824), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n755), .A2(new_n758), .A3(new_n810), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n800), .A2(new_n836), .A3(new_n801), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT116), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n827), .A2(new_n839), .A3(KEYINPUT54), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n835), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  AND4_X1   g656(.A1(KEYINPUT53), .A2(new_n755), .A3(new_n758), .A4(new_n810), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n828), .A2(new_n824), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n843), .A3(new_n837), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n488), .B1(new_n762), .B2(new_n763), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n725), .A2(new_n531), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n791), .A2(new_n792), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n702), .A2(new_n415), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n417), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n757), .B(new_n851), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n703), .A2(new_n735), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n849), .A2(new_n653), .A3(new_n726), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n684), .A2(new_n488), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n620), .A3(new_n856), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n611), .A2(new_n612), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n851), .A2(new_n494), .A3(new_n727), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n862), .A2(new_n863), .A3(new_n687), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n863), .B1(new_n862), .B2(new_n687), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n848), .A2(new_n855), .A3(KEYINPUT51), .A4(new_n866), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n855), .A2(new_n866), .B1(new_n848), .B2(KEYINPUT51), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n848), .A2(KEYINPUT51), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n849), .A2(new_n749), .A3(new_n856), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n851), .A2(new_n600), .A3(new_n727), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n871), .B(new_n872), .C1(new_n613), .C2(new_n859), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n847), .A2(new_n874), .A3(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(G952), .A3(new_n395), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n847), .A2(new_n874), .ZN(new_n877));
  OAI21_X1  g691(.A(G953), .B1(new_n877), .B2(KEYINPUT118), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n684), .A2(new_n627), .A3(new_n494), .A4(new_n760), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n531), .B1(new_n853), .B2(KEYINPUT49), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(KEYINPUT49), .B2(new_n853), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n687), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n878), .A3(new_n883), .ZN(G75));
  NAND2_X1  g698(.A1(new_n841), .A2(new_n845), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G902), .A3(new_n482), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n476), .B(new_n478), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n886), .A2(new_n887), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n886), .B2(new_n887), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n395), .A2(G952), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(G51));
  XNOR2_X1  g708(.A(new_n778), .B(KEYINPUT119), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT57), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n841), .A2(new_n842), .A3(new_n845), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n842), .B1(new_n841), .B2(new_n845), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(KEYINPUT120), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n411), .A3(new_n902), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n837), .A2(new_n838), .A3(new_n843), .A4(new_n844), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n834), .B2(new_n805), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n906), .A2(new_n250), .A3(new_n777), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n893), .B1(new_n903), .B2(new_n907), .ZN(G54));
  NOR2_X1   g722(.A1(new_n906), .A2(new_n250), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n230), .A3(new_n236), .ZN(new_n911));
  INV_X1    g725(.A(new_n893), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(new_n237), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G60));
  XNOR2_X1  g728(.A(new_n610), .B(KEYINPUT59), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n840), .B2(new_n846), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n603), .A2(new_n606), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n912), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n915), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n897), .C2(new_n898), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT122), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n847), .B2(new_n915), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n912), .A4(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n885), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n522), .A2(new_n523), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n893), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n885), .A2(new_n651), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT61), .B1(new_n935), .B2(KEYINPUT123), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n934), .B(new_n935), .C1(KEYINPUT123), .C2(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n395), .B1(new_n489), .B2(G224), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n832), .B2(new_n395), .ZN(new_n942));
  INV_X1    g756(.A(G898), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n476), .B1(new_n943), .B2(G953), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n942), .B(new_n944), .ZN(G69));
  XOR2_X1   g759(.A(new_n561), .B(new_n232), .Z(new_n946));
  AOI21_X1  g760(.A(new_n787), .B1(new_n793), .B2(new_n794), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n667), .A2(new_n699), .A3(new_n728), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n798), .A2(new_n749), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n755), .B(new_n758), .C1(new_n784), .C2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n946), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n948), .A2(new_n692), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n613), .B1(new_n612), .B2(new_n309), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n594), .A2(new_n670), .A3(new_n757), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n947), .A3(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n952), .B(new_n395), .C1(new_n946), .C2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n946), .A2(G227), .A3(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT124), .ZN(new_n962));
  AOI21_X1  g776(.A(G227), .B1(new_n946), .B2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g777(.A(G900), .ZN(new_n964));
  OAI21_X1  g778(.A(G953), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(G72));
  XNOR2_X1  g780(.A(new_n562), .B(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n955), .A2(new_n947), .A3(new_n825), .A4(new_n957), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n621), .A2(new_n250), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n967), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n541), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n949), .A2(new_n832), .A3(new_n951), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n583), .B(new_n967), .C1(new_n975), .C2(new_n971), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n971), .B1(new_n585), .B2(new_n571), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n827), .A2(new_n839), .A3(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n974), .A2(new_n912), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n893), .B1(new_n973), .B2(new_n541), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n982), .A2(KEYINPUT127), .A3(new_n976), .A4(new_n978), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(G57));
endmodule


