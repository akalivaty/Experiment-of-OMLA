//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT75), .B1(new_n188), .B2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n190), .A2(new_n191), .A3(new_n187), .A4(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G125), .B(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT74), .B1(new_n194), .B2(KEYINPUT16), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G140), .ZN(new_n197));
  AND4_X1   g011(.A1(KEYINPUT74), .A2(new_n188), .A3(new_n197), .A4(KEYINPUT16), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n193), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n193), .C1(new_n195), .C2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT17), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n205));
  INV_X1    g019(.A(G237), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G214), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n206), .A2(new_n207), .A3(G143), .A4(G214), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n205), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(new_n211), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT86), .A3(G131), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n204), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT87), .B1(new_n203), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n213), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT86), .B1(new_n215), .B2(G131), .ZN(new_n222));
  AOI211_X1 g036(.A(new_n205), .B(new_n213), .C1(new_n210), .C2(new_n211), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT17), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT87), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n224), .A2(new_n225), .A3(new_n201), .A4(new_n202), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT76), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n194), .B(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n200), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(new_n200), .B2(new_n194), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT18), .A2(G131), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n215), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n240));
  NOR2_X1   g054(.A1(G475), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT19), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n194), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n229), .B2(new_n242), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n200), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(new_n202), .A3(new_n220), .ZN(new_n246));
  INV_X1    g060(.A(new_n238), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n234), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n239), .A2(new_n240), .A3(new_n241), .A4(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT88), .ZN(new_n250));
  INV_X1    g064(.A(new_n248), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(new_n235), .B2(new_n238), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT88), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n240), .A4(new_n241), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n239), .A2(new_n241), .A3(new_n248), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n250), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT90), .ZN(new_n259));
  OR2_X1    g073(.A1(new_n238), .A2(KEYINPUT89), .ZN(new_n260));
  AOI21_X1  g074(.A(G902), .B1(new_n235), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n260), .B2(new_n235), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G475), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n259), .B1(new_n258), .B2(new_n263), .ZN(new_n265));
  NAND2_X1  g079(.A1(G234), .A2(G237), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n266), .A2(G952), .A3(new_n207), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n266), .A2(G902), .A3(G953), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT21), .B(G898), .Z(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT93), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n264), .A2(new_n265), .A3(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT9), .B(G234), .Z(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G221), .B1(new_n277), .B2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G101), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT78), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G107), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n284), .A3(G104), .ZN(new_n285));
  NOR2_X1   g099(.A1(G104), .A2(G107), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT3), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n281), .A2(KEYINPUT3), .A3(G104), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n280), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT78), .B(G107), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n286), .B1(new_n292), .B2(G104), .ZN(new_n293));
  OAI211_X1 g107(.A(G101), .B(new_n289), .C1(new_n293), .C2(KEYINPUT3), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n294), .A3(KEYINPUT4), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n200), .A2(G143), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n209), .A2(G146), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT0), .A2(G128), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G143), .B(G146), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT0), .A3(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n288), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n307), .A3(G101), .A4(new_n289), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n295), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT11), .ZN(new_n310));
  INV_X1    g124(.A(G134), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(G137), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(G137), .ZN(new_n313));
  INV_X1    g127(.A(G137), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT11), .A3(G134), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G131), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n312), .A2(new_n315), .A3(new_n213), .A4(new_n313), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT80), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n292), .A2(new_n237), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n281), .A2(G104), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n280), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n289), .B1(new_n293), .B2(KEYINPUT3), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n280), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT64), .ZN(new_n327));
  OAI21_X1  g141(.A(G128), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT64), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n298), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n302), .A2(new_n331), .A3(G128), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n325), .A2(KEYINPUT10), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n323), .ZN(new_n335));
  INV_X1    g149(.A(G128), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n296), .B2(KEYINPUT1), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n332), .B1(new_n337), .B2(new_n302), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n291), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n309), .A2(new_n320), .A3(new_n334), .A4(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n339), .B1(new_n325), .B2(new_n333), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n317), .A2(new_n318), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n344), .B2(KEYINPUT81), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n343), .B2(new_n344), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n207), .A2(G227), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n342), .A2(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n309), .A2(new_n334), .A3(new_n341), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n344), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n354), .A2(KEYINPUT82), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT82), .B1(new_n354), .B2(new_n358), .ZN(new_n360));
  OAI21_X1  g174(.A(G469), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G469), .ZN(new_n362));
  INV_X1    g176(.A(G902), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n357), .A2(new_n342), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n344), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n345), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n364), .B1(new_n372), .B2(new_n362), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n279), .B1(new_n361), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G119), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  INV_X1    g191(.A(G116), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n378), .A2(KEYINPUT66), .A3(G119), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT66), .B1(new_n378), .B2(G119), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G113), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT2), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G113), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT66), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n376), .B2(G116), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n378), .A2(KEYINPUT66), .A3(G119), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n377), .A3(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(KEYINPUT67), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n392), .A2(new_n377), .A3(new_n386), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n386), .B1(new_n392), .B2(new_n377), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n295), .A2(new_n394), .A3(new_n398), .A4(new_n308), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n392), .A3(new_n377), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(G113), .C1(new_n377), .C2(new_n400), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n325), .A2(new_n393), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(G110), .B(G122), .Z(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n405), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(new_n410), .A3(new_n405), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n304), .A2(G125), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n333), .B2(G125), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n207), .A2(G224), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT7), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n413), .B(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n392), .A2(KEYINPUT5), .A3(new_n377), .ZN(new_n420));
  OAI21_X1  g234(.A(G113), .B1(new_n400), .B2(new_n377), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n393), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n325), .A2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n405), .B(KEYINPUT8), .Z(new_n424));
  NAND2_X1  g238(.A1(new_n402), .A2(new_n393), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n423), .B(new_n424), .C1(new_n325), .C2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n408), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n363), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G210), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n416), .A2(new_n363), .A3(new_n429), .A4(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT84), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G214), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n435), .A3(new_n430), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n375), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G122), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G116), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT91), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n441), .A2(KEYINPUT14), .B1(G116), .B2(new_n439), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(KEYINPUT14), .B2(new_n441), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G107), .ZN(new_n444));
  INV_X1    g258(.A(new_n292), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(G116), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G128), .B(G143), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(new_n311), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n311), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(KEYINPUT13), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n209), .A2(G128), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n454), .B(G134), .C1(KEYINPUT13), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n447), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n445), .B1(new_n441), .B2(new_n446), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n453), .B(new_n456), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n277), .A2(new_n460), .A3(G953), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n452), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n452), .B2(new_n459), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G902), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(KEYINPUT15), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n465), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n275), .A2(new_n438), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT71), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n396), .A2(new_n397), .A3(new_n395), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT67), .B1(new_n388), .B2(new_n393), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n313), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n311), .A2(G137), .ZN(new_n476));
  OAI21_X1  g290(.A(G131), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n318), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n333), .A2(new_n479), .B1(new_n305), .B2(new_n344), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n398), .A2(KEYINPUT68), .A3(new_n394), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n474), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n480), .A4(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n304), .B1(new_n318), .B2(new_n317), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n478), .B1(new_n330), .B2(new_n332), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT30), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(KEYINPUT65), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n326), .A2(new_n327), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n296), .A2(KEYINPUT64), .A3(KEYINPUT1), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(G128), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n298), .A2(new_n336), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n494), .A2(new_n298), .B1(new_n495), .B2(new_n331), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n491), .B1(new_n496), .B2(new_n478), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n305), .A2(new_n344), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n489), .B1(new_n499), .B2(new_n488), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n472), .A2(new_n473), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n484), .A2(new_n485), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(G101), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n206), .A2(new_n207), .A3(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n470), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n482), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n484), .A2(new_n485), .B1(new_n501), .B2(new_n499), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n509), .B(new_n506), .C1(new_n510), .C2(new_n508), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n484), .A2(new_n485), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n499), .A2(new_n501), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT28), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n516), .A2(new_n470), .A3(new_n509), .A4(new_n506), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT29), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n480), .B1(new_n474), .B2(new_n481), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n484), .B2(new_n485), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n509), .B1(new_n521), .B2(new_n508), .ZN(new_n522));
  INV_X1    g336(.A(new_n506), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n518), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n363), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n499), .A2(new_n488), .ZN(new_n530));
  INV_X1    g344(.A(new_n489), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n501), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n513), .A2(new_n506), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n535));
  NAND4_X1  g349(.A1(new_n513), .A2(new_n532), .A3(new_n506), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n509), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n534), .B(new_n536), .C1(new_n538), .C2(new_n506), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n528), .A2(G472), .B1(new_n529), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n506), .B1(new_n516), .B2(new_n509), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n536), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT32), .B(new_n540), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n539), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n540), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT24), .B(G110), .Z(new_n551));
  XNOR2_X1  g365(.A(G119), .B(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n336), .A2(G119), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT23), .B1(new_n376), .B2(G128), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT23), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n336), .A3(G119), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n554), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G110), .B1(new_n558), .B2(KEYINPUT73), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n560), .B(new_n554), .C1(new_n555), .C2(new_n557), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n553), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n562), .B1(new_n201), .B2(new_n202), .ZN(new_n563));
  INV_X1    g377(.A(G110), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n552), .B2(new_n551), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n230), .A2(new_n566), .A3(new_n202), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT77), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n562), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n203), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT77), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n230), .A2(new_n566), .A3(new_n202), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT22), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(G137), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n568), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n570), .A2(new_n572), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(KEYINPUT77), .A3(new_n576), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT25), .B1(new_n581), .B2(G902), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n460), .B1(G234), .B2(new_n363), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT25), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n363), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n582), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n583), .A2(G902), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n550), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n469), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n280), .ZN(G3));
  OR3_X1    g408(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT33), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n462), .B2(new_n463), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(G478), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n465), .A2(new_n466), .ZN(new_n598));
  NAND2_X1  g412(.A1(G478), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n258), .A2(new_n263), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT90), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n258), .A2(new_n259), .A3(new_n263), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT96), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n431), .A2(new_n606), .A3(new_n432), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n428), .A2(KEYINPUT96), .A3(new_n430), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n434), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n605), .A2(new_n274), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n539), .A2(new_n363), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT94), .A3(G472), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n613));
  INV_X1    g427(.A(G472), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n539), .B(new_n363), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n612), .A2(new_n374), .A3(new_n591), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT97), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n618), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(new_n467), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n465), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n255), .B(new_n256), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n263), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n609), .A2(new_n625), .A3(new_n274), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n617), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT98), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n579), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n588), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n587), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n631), .B1(new_n587), .B2(new_n634), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n612), .B(new_n615), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n638), .A2(new_n275), .A3(new_n438), .A4(new_n468), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT37), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n564), .ZN(G12));
  NOR2_X1   g455(.A1(new_n635), .A2(new_n636), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n542), .B2(new_n549), .ZN(new_n643));
  INV_X1    g457(.A(new_n609), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n269), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n625), .B1(new_n268), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n643), .A2(new_n374), .A3(new_n644), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n587), .A2(new_n634), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n646), .A2(new_n268), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT39), .Z(new_n652));
  OR2_X1    g466(.A1(new_n375), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT40), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n547), .A2(new_n548), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n529), .B2(new_n541), .ZN(new_n656));
  INV_X1    g470(.A(new_n533), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n521), .A2(new_n506), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n363), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G472), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n433), .A2(new_n436), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT38), .Z(new_n663));
  AOI21_X1  g477(.A(new_n468), .B1(new_n602), .B2(new_n603), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n434), .A3(new_n664), .ZN(new_n665));
  OR4_X1    g479(.A1(new_n650), .A2(new_n654), .A3(new_n661), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  OR2_X1    g481(.A1(new_n635), .A2(new_n636), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n550), .A2(new_n374), .A3(new_n644), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n600), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n651), .C1(new_n264), .C2(new_n265), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(KEYINPUT100), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n643), .A2(new_n374), .A3(new_n644), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n675), .B2(new_n671), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI21_X1  g492(.A(new_n590), .B1(new_n542), .B2(new_n549), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n372), .A2(new_n680), .A3(new_n362), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n362), .ZN(new_n682));
  AOI211_X1 g496(.A(G902), .B(new_n682), .C1(new_n366), .C2(new_n371), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n681), .A2(new_n683), .A3(new_n279), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n610), .A2(new_n679), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND3_X1  g501(.A1(new_n679), .A2(new_n626), .A3(new_n684), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT102), .B(G116), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G18));
  NOR2_X1   g504(.A1(new_n681), .A2(new_n683), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n278), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n642), .A2(new_n692), .A3(new_n609), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(new_n550), .A3(new_n468), .A4(new_n275), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  INV_X1    g509(.A(new_n540), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n506), .B1(new_n522), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n697), .B2(new_n522), .ZN(new_n699));
  INV_X1    g513(.A(new_n544), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n614), .B1(new_n539), .B2(new_n363), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n590), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n703), .A2(new_n684), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n664), .A2(new_n705), .A3(new_n644), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n705), .B1(new_n664), .B2(new_n644), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n273), .B(new_n704), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT105), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(new_n702), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n699), .A2(new_n700), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n712), .B(new_n650), .C1(new_n713), .C2(new_n696), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n671), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n692), .A2(new_n609), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(KEYINPUT106), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n650), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n701), .A2(new_n718), .A3(new_n702), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n604), .A2(new_n716), .A3(new_n651), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  AOI21_X1  g538(.A(new_n352), .B1(new_n370), .B2(new_n342), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n357), .A2(new_n342), .A3(new_n352), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n279), .B1(new_n373), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n662), .A2(new_n434), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n604), .A2(new_n730), .A3(new_n651), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n542), .A2(new_n545), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(new_n591), .ZN(new_n734));
  AOI211_X1 g548(.A(KEYINPUT107), .B(new_n590), .C1(new_n542), .C2(new_n545), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n731), .B(KEYINPUT42), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n672), .A2(new_n679), .A3(new_n730), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  NAND4_X1  g555(.A1(new_n550), .A2(new_n730), .A3(new_n647), .A4(new_n591), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(new_n434), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n433), .B2(new_n436), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n602), .A2(new_n603), .A3(new_n670), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n612), .A2(new_n615), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n650), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n745), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n750), .A2(new_n751), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT108), .B(new_n745), .C1(new_n750), .C2(new_n751), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n727), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n364), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT46), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n362), .B2(new_n372), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n278), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n652), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n754), .A2(new_n769), .A3(new_n755), .A4(new_n756), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(new_n745), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n767), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(KEYINPUT47), .A3(new_n278), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n671), .B(new_n773), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n542), .A3(new_n549), .A4(new_n590), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  INV_X1    g593(.A(new_n691), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n590), .B1(new_n780), .B2(KEYINPUT49), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(KEYINPUT49), .B2(new_n780), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n663), .A2(new_n782), .A3(new_n279), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n746), .A2(new_n744), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n661), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n748), .A2(new_n267), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n663), .A2(new_n692), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n744), .A3(new_n703), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT50), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n789), .A2(KEYINPUT50), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(KEYINPUT50), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n775), .B(new_n776), .C1(new_n278), .C2(new_n780), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n786), .A2(new_n703), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n745), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n773), .A2(new_n692), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n661), .A2(new_n591), .A3(new_n267), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n602), .A2(new_n603), .A3(new_n600), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n786), .A2(new_n798), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n719), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n797), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g618(.A(G952), .B(new_n207), .C1(new_n794), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n790), .A2(new_n793), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n790), .A2(KEYINPUT118), .A3(new_n793), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n803), .A3(new_n797), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n278), .A2(new_n651), .ZN(new_n814));
  INV_X1    g628(.A(new_n708), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n706), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n373), .A2(new_n728), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n650), .B(new_n818), .C1(new_n656), .C2(new_n660), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n813), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT106), .B1(new_n715), .B2(new_n716), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n684), .A2(new_n608), .A3(new_n434), .A4(new_n607), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n671), .A2(new_n714), .A3(new_n822), .A4(new_n721), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n648), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT112), .B1(new_n723), .B2(new_n648), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n677), .B(new_n820), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n816), .A2(new_n819), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n717), .A2(new_n722), .B1(new_n669), .B2(new_n647), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n677), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n694), .A2(new_n688), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n685), .A2(new_n740), .A3(new_n709), .A4(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n604), .A2(new_n730), .A3(new_n651), .A4(new_n719), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n742), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n539), .A2(new_n540), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT29), .B1(new_n507), .B2(new_n511), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n526), .B1(new_n841), .B2(new_n517), .ZN(new_n842));
  OAI22_X1  g656(.A1(new_n840), .A2(KEYINPUT32), .B1(new_n842), .B2(new_n614), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n374), .B(new_n668), .C1(new_n655), .C2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n468), .A2(new_n263), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n745), .A2(new_n845), .A3(new_n624), .A4(new_n651), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT111), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n846), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n643), .A3(new_n374), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n742), .A4(new_n838), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n616), .ZN(new_n854));
  INV_X1    g668(.A(new_n437), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n855), .A3(new_n273), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n856), .A2(new_n605), .B1(new_n469), .B2(new_n592), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n264), .A2(new_n265), .A3(new_n468), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n859), .A3(new_n855), .A4(new_n273), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n639), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT110), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n639), .A2(new_n860), .A3(KEYINPUT110), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n858), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n829), .A2(new_n677), .A3(new_n813), .A4(new_n830), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n837), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT53), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT54), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n853), .B2(new_n865), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n639), .A2(new_n860), .A3(KEYINPUT110), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT110), .B1(new_n639), .B2(new_n860), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n877), .A3(new_n857), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n848), .A2(new_n852), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n878), .A2(KEYINPUT114), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n875), .A2(KEYINPUT53), .A3(new_n837), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n673), .A2(new_n676), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n824), .A2(new_n825), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n723), .A2(KEYINPUT112), .A3(new_n648), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n885), .A2(new_n820), .B1(new_n831), .B2(new_n832), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n873), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n880), .A2(new_n837), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n878), .A2(new_n879), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n835), .B1(new_n889), .B2(new_n874), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n834), .A3(KEYINPUT115), .A4(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n835), .B1(new_n869), .B2(new_n870), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n891), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n812), .A2(new_n872), .A3(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n734), .A2(new_n735), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n802), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT48), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n799), .A2(new_n605), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n796), .A2(new_n716), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT119), .Z(new_n902));
  NOR4_X1   g716(.A1(new_n896), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(G952), .A2(G953), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n785), .B1(new_n903), .B2(new_n904), .ZN(G75));
  NOR2_X1   g719(.A1(new_n207), .A2(G952), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT122), .Z(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n887), .A2(new_n894), .A3(new_n891), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G210), .A3(G902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n409), .A2(new_n411), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n415), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT120), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT55), .Z(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n912), .B2(new_n913), .ZN(new_n919));
  INV_X1    g733(.A(new_n918), .ZN(new_n920));
  AOI211_X1 g734(.A(KEYINPUT121), .B(new_n920), .C1(new_n910), .C2(new_n911), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n914), .A2(new_n919), .A3(new_n921), .ZN(G51));
  NAND2_X1  g736(.A1(new_n909), .A2(new_n892), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n923), .A2(KEYINPUT123), .A3(new_n895), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n909), .A2(new_n925), .A3(new_n892), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n364), .B(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n366), .A2(new_n371), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n761), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n909), .A2(G902), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n906), .B1(new_n930), .B2(new_n932), .ZN(G54));
  AND2_X1   g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(KEYINPUT124), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n909), .A2(G902), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n252), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n906), .ZN(G60));
  NAND2_X1  g755(.A1(new_n595), .A2(new_n596), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n895), .A2(new_n872), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n599), .B(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(new_n907), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n924), .A2(new_n942), .A3(new_n926), .A4(new_n944), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT60), .Z(new_n950));
  NAND3_X1  g764(.A1(new_n909), .A2(new_n633), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n909), .A2(new_n950), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n908), .B(new_n951), .C1(new_n952), .C2(new_n584), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G66));
  NAND4_X1  g769(.A1(new_n878), .A2(new_n685), .A3(new_n709), .A4(new_n836), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n207), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT126), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n207), .B1(new_n271), .B2(G224), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n915), .B1(G898), .B2(new_n207), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  OAI211_X1 g778(.A(new_n768), .B(new_n897), .C1(new_n707), .C2(new_n708), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n771), .A2(new_n778), .A3(new_n885), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n740), .A2(new_n742), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n966), .A2(G953), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n500), .B(new_n244), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n645), .A2(new_n207), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n885), .A2(new_n666), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT62), .Z(new_n976));
  OAI21_X1  g790(.A(new_n679), .B1(new_n604), .B2(new_n859), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n977), .A2(new_n653), .A3(new_n773), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n976), .A2(new_n771), .A3(new_n778), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n969), .B1(new_n979), .B2(new_n207), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n972), .A2(new_n974), .A3(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n973), .B1(new_n983), .B2(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(G72));
  INV_X1    g799(.A(new_n906), .ZN(new_n986));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n979), .B2(new_n957), .ZN(new_n989));
  INV_X1    g803(.A(new_n502), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n506), .A3(new_n990), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n966), .A2(new_n957), .A3(new_n967), .ZN(new_n992));
  INV_X1    g806(.A(new_n988), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n523), .B(new_n502), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n502), .B(new_n506), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n867), .A2(new_n871), .A3(new_n988), .A4(new_n995), .ZN(new_n996));
  AND4_X1   g810(.A1(new_n986), .A2(new_n991), .A3(new_n994), .A4(new_n996), .ZN(G57));
endmodule


