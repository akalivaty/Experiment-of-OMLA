//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(KEYINPUT65), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT3), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g047(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(KEYINPUT65), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n462), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n478), .A2(KEYINPUT3), .B1(new_n469), .B2(new_n471), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n479), .A2(KEYINPUT67), .A3(G137), .A4(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI22_X1  g060(.A1(new_n485), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n486), .A2(new_n467), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n478), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G101), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT68), .Z(G160));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n466), .A2(new_n472), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT69), .A3(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT69), .B1(new_n493), .B2(new_n467), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G124), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(KEYINPUT70), .A3(G124), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n493), .A2(G2105), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(new_n501), .B1(G136), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(G100), .A2(G2105), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(G162));
  NAND4_X1  g081(.A1(new_n466), .A2(G138), .A3(new_n467), .A4(new_n472), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n482), .A2(new_n483), .A3(G138), .A4(new_n467), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR3_X1    g086(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT72), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n467), .A2(G102), .A3(G2104), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT65), .B(G2104), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n472), .B(G126), .C1(new_n470), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G114), .A2(G2104), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n514), .B1(new_n518), .B2(G2105), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G164));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT6), .B(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  INV_X1    g107(.A(G50), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(G543), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n529), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  INV_X1    g112(.A(new_n534), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(G51), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n531), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT73), .B(G89), .Z(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n523), .A2(new_n525), .ZN(new_n547));
  INV_X1    g122(.A(G63), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  INV_X1    g128(.A(G52), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n531), .A2(new_n553), .B1(new_n554), .B2(new_n534), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n555), .B1(G651), .B2(new_n557), .ZN(G171));
  AOI22_X1  g133(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n528), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  INV_X1    g136(.A(G43), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n531), .A2(new_n561), .B1(new_n562), .B2(new_n534), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  AND3_X1   g140(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G36), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G188));
  XOR2_X1   g145(.A(KEYINPUT75), .B(G65), .Z(new_n571));
  AOI22_X1  g146(.A1(new_n526), .A2(new_n571), .B1(G78), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n528), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n531), .A2(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n538), .A2(G53), .A3(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n534), .A2(new_n579), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  NAND2_X1  g160(.A1(new_n542), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n538), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n531), .A2(new_n590), .B1(new_n591), .B2(new_n534), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n526), .A2(KEYINPUT76), .A3(G61), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n547), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n593), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n592), .B1(G651), .B2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n538), .A2(G47), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI221_X1 g178(.A(new_n601), .B1(new_n602), .B2(new_n531), .C1(new_n528), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n542), .A2(G92), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT10), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n528), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n538), .A2(G54), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n605), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n583), .ZN(G297));
  XNOR2_X1  g192(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n613), .B1(new_n619), .B2(G860), .ZN(G148));
  NOR2_X1   g195(.A1(new_n564), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n497), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n502), .A2(G135), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(KEYINPUT80), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(KEYINPUT80), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G111), .C2(new_n467), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n488), .A2(new_n485), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  NAND2_X1  g210(.A1(KEYINPUT79), .A2(G2100), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT13), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n633), .B(new_n638), .C1(KEYINPUT79), .C2(G2100), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2067), .B(G2678), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT17), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n662), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT82), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(KEYINPUT18), .B2(new_n658), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n665), .B(new_n668), .Z(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n671), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n675), .A2(KEYINPUT20), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n671), .A3(new_n674), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n678), .B(new_n680), .C1(KEYINPUT20), .C2(new_n675), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT84), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G23), .ZN(new_n690));
  INV_X1    g265(.A(G288), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT33), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1976), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n689), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT89), .B(G1971), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n689), .A2(G6), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n599), .B2(new_n689), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT88), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n694), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G24), .B(G290), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT86), .B(G1986), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G25), .ZN(new_n711));
  INV_X1    g286(.A(G119), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n495), .B2(new_n496), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n479), .A2(new_n467), .ZN(new_n715));
  INV_X1    g290(.A(G131), .ZN(new_n716));
  NOR2_X1   g291(.A1(G95), .A2(G2105), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n718));
  OAI22_X1  g293(.A1(new_n715), .A2(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OR3_X1    g294(.A1(new_n713), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n714), .B1(new_n713), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n711), .B1(new_n723), .B2(new_n710), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT35), .B(G1991), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n706), .A2(new_n709), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT36), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n689), .A2(G4), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n613), .B2(new_n689), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1348), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n632), .A2(new_n710), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(G1348), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n689), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n564), .B2(new_n689), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G1341), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n732), .A2(new_n733), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n710), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n710), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2078), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G5), .B2(G16), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n742), .A2(G5), .A3(G16), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n743), .B(new_n744), .C1(G301), .C2(new_n689), .ZN(new_n745));
  INV_X1    g320(.A(G1961), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G11), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n745), .A2(new_n746), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n710), .B1(new_n750), .B2(G28), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT94), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n750), .A2(G28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  NOR3_X1   g332(.A1(new_n738), .A2(new_n741), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(G160), .A2(G29), .B1(KEYINPUT92), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT92), .B2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2084), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n758), .B(new_n765), .C1(G1341), .C2(new_n736), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT93), .B1(G16), .B2(G21), .ZN(new_n767));
  NAND2_X1  g342(.A1(G168), .A2(G16), .ZN(new_n768));
  MUX2_X1   g343(.A(KEYINPUT93), .B(new_n767), .S(new_n768), .Z(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT95), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n689), .A2(G20), .ZN(new_n773));
  OAI211_X1 g348(.A(KEYINPUT23), .B(new_n773), .C1(new_n583), .C2(new_n689), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT23), .B2(new_n773), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n710), .A2(G33), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(new_n467), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n502), .A2(G139), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(new_n710), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT91), .Z(new_n787));
  AOI21_X1  g362(.A(new_n777), .B1(G2072), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n496), .ZN(new_n789));
  OAI21_X1  g364(.A(G129), .B1(new_n789), .B2(new_n494), .ZN(new_n790));
  NAND3_X1  g365(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT26), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n488), .A2(G105), .ZN(new_n794));
  INV_X1    g369(.A(G141), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n715), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n790), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G32), .B(new_n798), .S(G29), .Z(new_n799));
  XOR2_X1   g374(.A(KEYINPUT27), .B(G1996), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n769), .A2(new_n770), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n787), .A2(G2072), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n772), .A2(new_n788), .A3(new_n801), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G140), .ZN(new_n806));
  NOR2_X1   g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n715), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n497), .B2(G128), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n710), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n710), .A2(G26), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT28), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(KEYINPUT28), .B2(new_n812), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT90), .B(G2067), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n766), .A2(new_n805), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n710), .A2(G35), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G162), .B2(new_n710), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT29), .B(G2090), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n729), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(G311));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n822), .B(new_n824), .ZN(G150));
  NAND2_X1  g400(.A1(new_n542), .A2(G93), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT98), .B(G55), .Z(new_n828));
  OAI221_X1 g403(.A(new_n826), .B1(new_n528), .B2(new_n827), .C1(new_n534), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n613), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n829), .B(new_n564), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT39), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n831), .B1(new_n836), .B2(G860), .ZN(G145));
  XNOR2_X1  g412(.A(G160), .B(new_n632), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G162), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n520), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n798), .A2(new_n810), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n798), .A2(new_n810), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n798), .A2(new_n810), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n520), .A2(new_n842), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT99), .B1(new_n513), .B2(new_n519), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n851), .A3(new_n844), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n847), .A2(KEYINPUT100), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT100), .B1(new_n847), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n784), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n784), .B1(new_n847), .B2(new_n852), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n841), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n845), .A2(new_n843), .A3(new_n846), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n851), .B1(new_n848), .B2(new_n844), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n847), .A2(new_n852), .A3(KEYINPUT100), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n785), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n502), .A2(G142), .ZN(new_n866));
  INV_X1    g441(.A(G130), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT102), .B1(new_n498), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n497), .A2(new_n869), .A3(G130), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n467), .A2(G118), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n720), .A2(new_n635), .A3(new_n721), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n635), .B1(new_n720), .B2(new_n721), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n635), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n722), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n873), .ZN(new_n880));
  AOI211_X1 g455(.A(new_n880), .B(new_n866), .C1(new_n868), .C2(new_n870), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n720), .A2(new_n635), .A3(new_n721), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n877), .A2(new_n883), .A3(KEYINPUT103), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n877), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n858), .A2(new_n865), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n877), .A2(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n877), .A2(new_n883), .A3(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT101), .B1(new_n864), .B2(new_n856), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n855), .A2(new_n841), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n840), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n892), .A3(new_n894), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n858), .A2(new_n865), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(new_n839), .C1(new_n899), .C2(new_n888), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT104), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n896), .A2(new_n900), .A3(new_n903), .A4(new_n897), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n902), .A2(KEYINPUT40), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT40), .B1(new_n902), .B2(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(G395));
  INV_X1    g482(.A(G868), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n829), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n612), .B(G299), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT41), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n622), .B(new_n834), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  XNOR2_X1  g490(.A(G305), .B(G303), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n691), .B(G290), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(KEYINPUT105), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(KEYINPUT105), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT106), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n915), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n909), .B1(new_n922), .B2(new_n908), .ZN(G295));
  OAI21_X1  g498(.A(new_n909), .B1(new_n922), .B2(new_n908), .ZN(G331));
  XNOR2_X1  g499(.A(new_n834), .B(G286), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G301), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n911), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n910), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n920), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n897), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(KEYINPUT107), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n933), .A2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT44), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n934), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n931), .A2(KEYINPUT43), .A3(new_n897), .A4(new_n932), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(KEYINPUT44), .B2(new_n941), .ZN(G397));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n851), .B2(G1384), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n481), .A2(new_n487), .A3(G40), .A4(new_n489), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(KEYINPUT108), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G2067), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n810), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT109), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(new_n954), .A3(new_n951), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n798), .B(G1996), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n953), .A2(new_n955), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n722), .A2(new_n725), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n723), .A2(new_n726), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n949), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(G290), .B(G1986), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n949), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  NOR2_X1   g539(.A1(G168), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n520), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT111), .B1(new_n967), .B2(new_n945), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n513), .B2(new_n519), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT45), .ZN(new_n970));
  INV_X1    g545(.A(new_n945), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(new_n972), .C1(KEYINPUT45), .C2(new_n969), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n770), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n520), .A2(new_n977), .A3(new_n966), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n971), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n969), .B2(new_n977), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n520), .A2(new_n966), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G2084), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n975), .A2(new_n976), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n976), .B1(new_n975), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n965), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT118), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n991), .B(new_n965), .C1(new_n987), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT62), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n770), .A2(new_n974), .B1(new_n984), .B2(new_n985), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT119), .B1(new_n995), .B2(new_n964), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n975), .A2(new_n986), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n965), .A2(KEYINPUT51), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n987), .A2(new_n988), .A3(G286), .ZN(new_n1002));
  NAND2_X1  g577(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n993), .A2(new_n994), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT121), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G2078), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n974), .A2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT120), .B(G1961), .Z(new_n1011));
  NOR2_X1   g586(.A1(new_n984), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1006), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n983), .A2(new_n981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n945), .B1(new_n969), .B2(new_n977), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1011), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(KEYINPUT121), .C1(new_n974), .C2(new_n1009), .ZN(new_n1019));
  OR2_X1    g594(.A1(KEYINPUT122), .A2(KEYINPUT53), .ZN(new_n1020));
  NAND2_X1  g595(.A1(KEYINPUT122), .A2(KEYINPUT53), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT45), .B(new_n966), .C1(new_n849), .C2(new_n850), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n967), .A2(new_n945), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1020), .B(new_n1021), .C1(new_n1024), .C2(G2078), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1013), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1026), .A2(G171), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n982), .A2(new_n945), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n964), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  NOR2_X1   g606(.A1(G288), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n599), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(KEYINPUT49), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1029), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1029), .B(new_n1041), .C1(new_n1031), .C2(G288), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1033), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT55), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2090), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n984), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1050));
  OAI211_X1 g625(.A(G8), .B(new_n1046), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1015), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2090), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1045), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1043), .A2(new_n1051), .A3(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1027), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1005), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1005), .B2(new_n1058), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n994), .B1(new_n993), .B2(new_n1004), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n1065));
  OAI21_X1  g640(.A(G8), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1045), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n997), .A2(G8), .A3(G168), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1068), .A2(KEYINPUT112), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(KEYINPUT112), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1064), .B(new_n1067), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1057), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1065), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1068), .B(KEYINPUT112), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(KEYINPUT113), .A3(new_n1064), .A4(new_n1067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1040), .A2(new_n1031), .A3(new_n691), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1030), .B1(new_n1079), .B2(new_n1036), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1051), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n1043), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT56), .B(G2072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1022), .A2(new_n1023), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n573), .B2(new_n575), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT114), .ZN(new_n1086));
  OAI221_X1 g661(.A(new_n1086), .B1(new_n531), .B2(new_n574), .C1(new_n572), .C2(new_n528), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1087), .A3(new_n581), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(KEYINPUT115), .A3(new_n1089), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1092), .B(new_n1093), .C1(new_n1089), .C2(G299), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1053), .A2(new_n776), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1084), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1094), .B1(new_n1084), .B2(new_n1095), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT116), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT61), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  OAI211_X1 g675(.A(KEYINPUT116), .B(new_n1100), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n984), .A2(G1348), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1028), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2067), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(KEYINPUT60), .A3(new_n612), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1108));
  OAI221_X1 g683(.A(KEYINPUT60), .B1(G2067), .B2(new_n1103), .C1(new_n984), .C2(G1348), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n613), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1099), .A2(new_n1101), .A3(new_n1106), .A4(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1024), .A2(G1996), .B1(new_n1028), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n564), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT59), .Z(new_n1115));
  NOR2_X1   g690(.A1(new_n1105), .A2(new_n612), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1097), .ZN(new_n1117));
  OAI22_X1  g692(.A1(new_n1111), .A2(new_n1115), .B1(new_n1096), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n993), .A2(new_n1004), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n944), .A2(new_n971), .A3(new_n1022), .A4(new_n1008), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1025), .A2(new_n1018), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT54), .B(new_n1122), .C1(new_n1026), .C2(G171), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1118), .A2(new_n1119), .A3(new_n1057), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1121), .A2(G171), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1125), .B(new_n1126), .C1(new_n1027), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1026), .B2(G171), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n1129), .B2(KEYINPUT54), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1078), .B(new_n1082), .C1(new_n1124), .C2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n963), .B1(new_n1063), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n957), .A2(new_n958), .B1(new_n950), .B2(new_n810), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n947), .A2(new_n948), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1135), .A2(G1986), .A3(G290), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT48), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1134), .A2(new_n1135), .B1(new_n961), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT46), .ZN(new_n1139));
  OR3_X1    g714(.A1(new_n1135), .A2(new_n1139), .A3(G1996), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n951), .A2(new_n798), .ZN(new_n1141));
  OR3_X1    g716(.A1(new_n1135), .A2(KEYINPUT125), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT125), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1139), .B1(new_n1135), .B2(G1996), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1146));
  XNOR2_X1  g721(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1138), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1133), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g724(.A1(new_n902), .A2(new_n904), .ZN(new_n1151));
  INV_X1    g725(.A(G227), .ZN(new_n1152));
  NOR2_X1   g726(.A1(G229), .A2(new_n460), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n653), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g728(.A(new_n1154), .B(KEYINPUT127), .ZN(new_n1155));
  AND4_X1   g729(.A1(new_n1151), .A2(new_n939), .A3(new_n940), .A4(new_n1155), .ZN(G308));
  NAND4_X1  g730(.A1(new_n1151), .A2(new_n939), .A3(new_n940), .A4(new_n1155), .ZN(G225));
endmodule


