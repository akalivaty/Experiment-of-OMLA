

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761;

  NAND2_X1 U372 ( .A1(n457), .A2(n455), .ZN(n759) );
  OR2_X1 U373 ( .A1(n611), .A2(n456), .ZN(n455) );
  XNOR2_X1 U374 ( .A(n464), .B(n735), .ZN(n646) );
  NAND2_X1 U375 ( .A1(G234), .A2(G237), .ZN(n527) );
  BUF_X1 U376 ( .A(n643), .Z(n732) );
  INV_X2 U377 ( .A(G128), .ZN(n494) );
  XNOR2_X2 U378 ( .A(n350), .B(KEYINPUT76), .ZN(n574) );
  NAND2_X1 U379 ( .A1(n533), .A2(n532), .ZN(n350) );
  XNOR2_X1 U380 ( .A(n417), .B(n542), .ZN(n467) );
  OR2_X2 U381 ( .A1(n438), .A2(KEYINPUT93), .ZN(n437) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n505) );
  BUF_X1 U383 ( .A(n582), .Z(n688) );
  NOR2_X1 U384 ( .A1(n611), .A2(n614), .ZN(n352) );
  AND2_X2 U385 ( .A1(n436), .A2(n437), .ZN(n401) );
  NAND2_X2 U386 ( .A1(n595), .A2(n655), .ZN(n432) );
  XNOR2_X2 U387 ( .A(n547), .B(n546), .ZN(n595) );
  XNOR2_X2 U388 ( .A(n438), .B(n375), .ZN(n683) );
  NOR2_X1 U389 ( .A1(n680), .A2(n562), .ZN(n563) );
  INV_X4 U390 ( .A(KEYINPUT4), .ZN(n371) );
  INV_X2 U391 ( .A(G953), .ZN(n753) );
  AND2_X1 U392 ( .A1(n459), .A2(n458), .ZN(n457) );
  XNOR2_X1 U393 ( .A(n477), .B(KEYINPUT33), .ZN(n717) );
  NOR2_X1 U394 ( .A1(n393), .A2(n562), .ZN(n532) );
  NAND2_X1 U395 ( .A1(n401), .A2(n434), .ZN(n393) );
  XNOR2_X1 U396 ( .A(n559), .B(n450), .ZN(n575) );
  XNOR2_X1 U397 ( .A(n370), .B(n473), .ZN(n650) );
  XNOR2_X1 U398 ( .A(n397), .B(n394), .ZN(n726) );
  NAND2_X1 U399 ( .A1(n498), .A2(n402), .ZN(n555) );
  XNOR2_X1 U400 ( .A(n504), .B(n462), .ZN(n538) );
  INV_X1 U401 ( .A(G143), .ZN(n495) );
  XNOR2_X1 U402 ( .A(G902), .B(KEYINPUT15), .ZN(n543) );
  INV_X1 U403 ( .A(n760), .ZN(n353) );
  INV_X1 U404 ( .A(n353), .ZN(n354) );
  NOR2_X2 U405 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X2 U406 ( .A(n520), .B(KEYINPUT70), .ZN(n374) );
  XNOR2_X2 U407 ( .A(n371), .B(G101), .ZN(n520) );
  AND2_X1 U408 ( .A1(n634), .A2(n411), .ZN(n581) );
  INV_X1 U409 ( .A(n538), .ZN(n474) );
  AND2_X1 U410 ( .A1(n713), .A2(n644), .ZN(n413) );
  INV_X1 U411 ( .A(n543), .ZN(n644) );
  INV_X1 U412 ( .A(KEYINPUT46), .ZN(n422) );
  XNOR2_X1 U413 ( .A(n577), .B(KEYINPUT103), .ZN(n634) );
  INV_X1 U414 ( .A(n628), .ZN(n381) );
  AND2_X1 U415 ( .A1(n627), .A2(KEYINPUT44), .ZN(n382) );
  XNOR2_X1 U416 ( .A(n421), .B(KEYINPUT20), .ZN(n513) );
  XNOR2_X1 U417 ( .A(n503), .B(n476), .ZN(n475) );
  XNOR2_X1 U418 ( .A(n506), .B(KEYINPUT5), .ZN(n476) );
  INV_X1 U419 ( .A(KEYINPUT3), .ZN(n462) );
  AND2_X1 U420 ( .A1(n445), .A2(G134), .ZN(n468) );
  XNOR2_X1 U421 ( .A(n510), .B(n511), .ZN(n558) );
  INV_X1 U422 ( .A(KEYINPUT17), .ZN(n418) );
  XNOR2_X1 U423 ( .A(G110), .B(KEYINPUT18), .ZN(n466) );
  AND2_X1 U424 ( .A1(n756), .A2(n372), .ZN(n446) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n441) );
  OR2_X1 U426 ( .A1(G237), .A2(G902), .ZN(n544) );
  INV_X1 U427 ( .A(n617), .ZN(n430) );
  XNOR2_X1 U428 ( .A(n551), .B(n550), .ZN(n572) );
  XNOR2_X1 U429 ( .A(n549), .B(G475), .ZN(n550) );
  OR2_X2 U430 ( .A1(n679), .A2(n680), .ZN(n684) );
  XNOR2_X1 U431 ( .A(n604), .B(KEYINPUT0), .ZN(n615) );
  INV_X1 U432 ( .A(G469), .ZN(n377) );
  XNOR2_X1 U433 ( .A(G128), .B(G119), .ZN(n512) );
  XNOR2_X1 U434 ( .A(KEYINPUT24), .B(G110), .ZN(n433) );
  INV_X1 U435 ( .A(KEYINPUT10), .ZN(n398) );
  XNOR2_X1 U436 ( .A(n523), .B(KEYINPUT23), .ZN(n395) );
  XOR2_X1 U437 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n553) );
  XNOR2_X1 U438 ( .A(KEYINPUT7), .B(G122), .ZN(n552) );
  XNOR2_X1 U439 ( .A(n555), .B(KEYINPUT97), .ZN(n453) );
  XNOR2_X1 U440 ( .A(n672), .B(n447), .ZN(n594) );
  INV_X1 U441 ( .A(KEYINPUT102), .ZN(n447) );
  XNOR2_X1 U442 ( .A(n683), .B(n388), .ZN(n607) );
  INV_X1 U443 ( .A(KEYINPUT87), .ZN(n388) );
  INV_X1 U444 ( .A(G478), .ZN(n450) );
  NOR2_X1 U445 ( .A1(G902), .A2(n721), .ZN(n559) );
  AND2_X1 U446 ( .A1(n413), .A2(G469), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n410), .B(KEYINPUT79), .ZN(n385) );
  INV_X1 U448 ( .A(G134), .ZN(n497) );
  AND2_X1 U449 ( .A1(n590), .A2(n444), .ZN(n443) );
  INV_X1 U450 ( .A(n666), .ZN(n444) );
  NOR2_X1 U451 ( .A1(n653), .A2(n358), .ZN(n378) );
  INV_X1 U452 ( .A(G140), .ZN(n488) );
  XNOR2_X1 U453 ( .A(n487), .B(n427), .ZN(n426) );
  XOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n487) );
  XOR2_X1 U455 ( .A(G143), .B(KEYINPUT95), .Z(n427) );
  XNOR2_X1 U456 ( .A(n523), .B(KEYINPUT90), .ZN(n742) );
  XNOR2_X1 U457 ( .A(n522), .B(n356), .ZN(n485) );
  XOR2_X1 U458 ( .A(G104), .B(KEYINPUT78), .Z(n522) );
  XNOR2_X1 U459 ( .A(G110), .B(G107), .ZN(n521) );
  XNOR2_X1 U460 ( .A(n642), .B(n597), .ZN(n711) );
  OR2_X1 U461 ( .A1(n607), .A2(n636), .ZN(n461) );
  XOR2_X1 U462 ( .A(KEYINPUT77), .B(KEYINPUT92), .Z(n515) );
  XNOR2_X1 U463 ( .A(n500), .B(n474), .ZN(n473) );
  XNOR2_X1 U464 ( .A(n392), .B(n475), .ZN(n370) );
  XNOR2_X1 U465 ( .A(n467), .B(n465), .ZN(n464) );
  XNOR2_X1 U466 ( .A(n374), .B(n466), .ZN(n465) );
  INV_X1 U467 ( .A(KEYINPUT105), .ZN(n478) );
  BUF_X1 U468 ( .A(n711), .Z(n750) );
  OR2_X1 U469 ( .A1(n643), .A2(n470), .ZN(n713) );
  NAND2_X1 U470 ( .A1(n471), .A2(KEYINPUT2), .ZN(n470) );
  AND2_X1 U471 ( .A1(n428), .A2(n655), .ZN(n584) );
  NOR2_X1 U472 ( .A1(n598), .A2(n429), .ZN(n428) );
  OR2_X1 U473 ( .A1(n695), .A2(n605), .ZN(n423) );
  NOR2_X1 U474 ( .A1(n591), .A2(n585), .ZN(n425) );
  XNOR2_X1 U475 ( .A(n618), .B(KEYINPUT81), .ZN(n619) );
  AND2_X1 U476 ( .A1(n386), .A2(n430), .ZN(n620) );
  NAND2_X1 U477 ( .A1(n355), .A2(KEYINPUT32), .ZN(n458) );
  OR2_X1 U478 ( .A1(n461), .A2(n614), .ZN(n355) );
  INV_X1 U479 ( .A(KEYINPUT19), .ZN(n578) );
  NOR2_X1 U480 ( .A1(n684), .A2(n439), .ZN(n435) );
  BUF_X1 U481 ( .A(n615), .Z(n630) );
  INV_X1 U482 ( .A(KEYINPUT1), .ZN(n375) );
  XNOR2_X1 U483 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U484 ( .A(n400), .B(n743), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n433), .B(n512), .ZN(n396) );
  XNOR2_X1 U486 ( .A(n452), .B(n451), .ZN(n721) );
  XNOR2_X1 U487 ( .A(n359), .B(n557), .ZN(n451) );
  XNOR2_X1 U488 ( .A(n556), .B(n453), .ZN(n452) );
  INV_X1 U489 ( .A(KEYINPUT101), .ZN(n448) );
  NAND2_X1 U490 ( .A1(n481), .A2(n480), .ZN(n479) );
  XNOR2_X1 U491 ( .A(n482), .B(n365), .ZN(n481) );
  XNOR2_X1 U492 ( .A(n383), .B(n367), .ZN(G75) );
  OR2_X1 U493 ( .A1(n385), .A2(n384), .ZN(n383) );
  OR2_X1 U494 ( .A1(n715), .A2(n362), .ZN(n384) );
  AND2_X1 U495 ( .A1(G227), .A2(n753), .ZN(n356) );
  INV_X1 U496 ( .A(KEYINPUT93), .ZN(n439) );
  AND2_X1 U497 ( .A1(G210), .A2(n544), .ZN(n357) );
  AND2_X1 U498 ( .A1(n635), .A2(n634), .ZN(n358) );
  INV_X2 U499 ( .A(G146), .ZN(n399) );
  AND2_X1 U500 ( .A1(G217), .A2(n558), .ZN(n359) );
  INV_X1 U501 ( .A(n372), .ZN(n677) );
  AND2_X1 U502 ( .A1(n598), .A2(n460), .ZN(n360) );
  XOR2_X1 U503 ( .A(KEYINPUT73), .B(KEYINPUT22), .Z(n361) );
  NAND2_X1 U504 ( .A1(n718), .A2(n753), .ZN(n362) );
  INV_X1 U505 ( .A(KEYINPUT32), .ZN(n460) );
  XNOR2_X1 U506 ( .A(n548), .B(KEYINPUT59), .ZN(n363) );
  XNOR2_X1 U507 ( .A(n651), .B(KEYINPUT110), .ZN(n364) );
  XOR2_X1 U508 ( .A(n719), .B(n720), .Z(n365) );
  XOR2_X1 U509 ( .A(n648), .B(n647), .Z(n366) );
  INV_X1 U510 ( .A(n728), .ZN(n480) );
  XOR2_X1 U511 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n367) );
  XOR2_X1 U512 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n368) );
  XOR2_X1 U513 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n369) );
  XNOR2_X1 U514 ( .A(n374), .B(n521), .ZN(n524) );
  INV_X1 U515 ( .A(n373), .ZN(n585) );
  NAND2_X1 U516 ( .A1(n373), .A2(n698), .ZN(n454) );
  XNOR2_X2 U517 ( .A(n545), .B(n357), .ZN(n373) );
  OR2_X1 U518 ( .A1(n593), .A2(n373), .ZN(n372) );
  INV_X1 U519 ( .A(n438), .ZN(n376) );
  XNOR2_X2 U520 ( .A(n526), .B(n377), .ZN(n438) );
  NOR2_X1 U521 ( .A1(n568), .A2(n376), .ZN(n579) );
  NAND2_X1 U522 ( .A1(n379), .A2(n378), .ZN(n639) );
  NAND2_X1 U523 ( .A1(n380), .A2(n625), .ZN(n379) );
  NAND2_X1 U524 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U525 ( .A(n387), .B(n616), .ZN(n386) );
  NAND2_X1 U526 ( .A1(n717), .A2(n630), .ZN(n387) );
  XNOR2_X2 U527 ( .A(G137), .B(G140), .ZN(n523) );
  INV_X1 U528 ( .A(n683), .ZN(n609) );
  AND2_X4 U529 ( .A1(n414), .A2(n413), .ZN(n390) );
  NAND2_X1 U530 ( .A1(n389), .A2(n414), .ZN(n482) );
  NAND2_X1 U531 ( .A1(n390), .A2(G475), .ZN(n645) );
  NAND2_X1 U532 ( .A1(n390), .A2(G210), .ZN(n649) );
  NAND2_X1 U533 ( .A1(n390), .A2(G472), .ZN(n652) );
  NAND2_X1 U534 ( .A1(n390), .A2(G478), .ZN(n722) );
  NAND2_X1 U535 ( .A1(n390), .A2(G217), .ZN(n725) );
  NAND2_X1 U536 ( .A1(n608), .A2(n698), .ZN(n508) );
  XNOR2_X2 U537 ( .A(n582), .B(KEYINPUT104), .ZN(n608) );
  XNOR2_X2 U538 ( .A(n391), .B(G472), .ZN(n582) );
  OR2_X2 U539 ( .A1(n650), .A2(G902), .ZN(n391) );
  XNOR2_X1 U540 ( .A(n392), .B(n399), .ZN(n525) );
  XNOR2_X1 U541 ( .A(n392), .B(KEYINPUT4), .ZN(n744) );
  XNOR2_X2 U542 ( .A(n555), .B(n499), .ZN(n392) );
  NOR2_X1 U543 ( .A1(n393), .A2(n688), .ZN(n629) );
  XNOR2_X2 U544 ( .A(n539), .B(n398), .ZN(n743) );
  XNOR2_X2 U545 ( .A(n399), .B(G125), .ZN(n539) );
  NAND2_X1 U546 ( .A1(n558), .A2(G221), .ZN(n400) );
  XNOR2_X1 U547 ( .A(n514), .B(n515), .ZN(n517) );
  NAND2_X1 U548 ( .A1(n543), .A2(G234), .ZN(n421) );
  NAND2_X1 U549 ( .A1(n496), .A2(n497), .ZN(n402) );
  NAND2_X1 U550 ( .A1(n435), .A2(n438), .ZN(n434) );
  XNOR2_X1 U551 ( .A(n403), .B(n368), .ZN(G60) );
  NAND2_X1 U552 ( .A1(n409), .A2(n480), .ZN(n403) );
  XNOR2_X1 U553 ( .A(n404), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U554 ( .A1(n408), .A2(n480), .ZN(n404) );
  NAND2_X2 U555 ( .A1(n405), .A2(n415), .ZN(n414) );
  OR2_X2 U556 ( .A1(n641), .A2(n643), .ZN(n405) );
  INV_X1 U557 ( .A(KEYINPUT2), .ZN(n415) );
  NAND2_X1 U558 ( .A1(n406), .A2(n443), .ZN(n442) );
  XNOR2_X1 U559 ( .A(n571), .B(n422), .ZN(n406) );
  XNOR2_X1 U560 ( .A(n407), .B(n369), .ZN(G51) );
  NAND2_X1 U561 ( .A1(n424), .A2(n480), .ZN(n407) );
  XNOR2_X1 U562 ( .A(n652), .B(n364), .ZN(n408) );
  XNOR2_X1 U563 ( .A(n645), .B(n363), .ZN(n409) );
  NAND2_X1 U564 ( .A1(n714), .A2(n713), .ZN(n410) );
  NOR2_X1 U565 ( .A1(n640), .A2(n639), .ZN(n472) );
  NOR2_X1 U566 ( .A1(G902), .A2(n548), .ZN(n551) );
  XNOR2_X1 U567 ( .A(n536), .B(n426), .ZN(n491) );
  INV_X1 U568 ( .A(n634), .ZN(n696) );
  INV_X1 U569 ( .A(n667), .ZN(n411) );
  NAND2_X1 U570 ( .A1(n575), .A2(n576), .ZN(n449) );
  XNOR2_X1 U571 ( .A(n649), .B(n366), .ZN(n424) );
  NAND2_X1 U572 ( .A1(n412), .A2(n415), .ZN(n714) );
  NAND2_X1 U573 ( .A1(n712), .A2(n750), .ZN(n412) );
  NAND2_X1 U574 ( .A1(n684), .A2(n439), .ZN(n436) );
  XNOR2_X1 U575 ( .A(n454), .B(n578), .ZN(n603) );
  XNOR2_X2 U576 ( .A(n416), .B(n361), .ZN(n611) );
  NAND2_X1 U577 ( .A1(n615), .A2(n606), .ZN(n416) );
  XNOR2_X1 U578 ( .A(n539), .B(n418), .ZN(n417) );
  NOR2_X1 U579 ( .A1(n719), .A2(G902), .ZN(n526) );
  XNOR2_X2 U580 ( .A(n620), .B(n619), .ZN(n627) );
  XNOR2_X2 U581 ( .A(n419), .B(KEYINPUT85), .ZN(n628) );
  NAND2_X1 U582 ( .A1(n759), .A2(n663), .ZN(n419) );
  NAND2_X1 U583 ( .A1(n420), .A2(n360), .ZN(n456) );
  INV_X1 U584 ( .A(n461), .ZN(n420) );
  XNOR2_X1 U585 ( .A(n537), .B(n536), .ZN(n463) );
  XNOR2_X2 U586 ( .A(n423), .B(KEYINPUT41), .ZN(n716) );
  NOR2_X2 U587 ( .A1(n574), .A2(n569), .ZN(n547) );
  XNOR2_X1 U588 ( .A(n442), .B(n441), .ZN(n440) );
  XNOR2_X1 U589 ( .A(n711), .B(KEYINPUT75), .ZN(n641) );
  INV_X1 U590 ( .A(n425), .ZN(n586) );
  INV_X1 U591 ( .A(n583), .ZN(n429) );
  NAND2_X1 U592 ( .A1(n431), .A2(n614), .ZN(n477) );
  XNOR2_X1 U593 ( .A(n631), .B(n478), .ZN(n431) );
  XNOR2_X1 U594 ( .A(n628), .B(n613), .ZN(n621) );
  NAND2_X1 U595 ( .A1(n760), .A2(n761), .ZN(n571) );
  XNOR2_X2 U596 ( .A(n432), .B(n561), .ZN(n760) );
  XNOR2_X2 U597 ( .A(n519), .B(n518), .ZN(n679) );
  NAND2_X1 U598 ( .A1(n440), .A2(n446), .ZN(n642) );
  NAND2_X1 U599 ( .A1(n445), .A2(n469), .ZN(n496) );
  NAND2_X1 U600 ( .A1(n495), .A2(G128), .ZN(n445) );
  XNOR2_X2 U601 ( .A(n449), .B(n448), .ZN(n672) );
  NOR2_X2 U602 ( .A1(n607), .A2(n588), .ZN(n675) );
  NAND2_X1 U603 ( .A1(n611), .A2(KEYINPUT32), .ZN(n459) );
  XNOR2_X2 U604 ( .A(n463), .B(n538), .ZN(n735) );
  INV_X1 U605 ( .A(n496), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n468), .A2(n469), .ZN(n498) );
  NAND2_X1 U607 ( .A1(n494), .A2(G143), .ZN(n469) );
  INV_X1 U608 ( .A(n642), .ZN(n471) );
  XNOR2_X1 U609 ( .A(n472), .B(KEYINPUT45), .ZN(n643) );
  XNOR2_X1 U610 ( .A(n479), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U611 ( .A(n483), .B(n525), .ZN(n719) );
  XNOR2_X1 U612 ( .A(n524), .B(n484), .ZN(n483) );
  XNOR2_X1 U613 ( .A(n485), .B(n742), .ZN(n484) );
  XNOR2_X2 U614 ( .A(n560), .B(KEYINPUT100), .ZN(n655) );
  NOR2_X2 U615 ( .A1(n576), .A2(n575), .ZN(n560) );
  XOR2_X2 U616 ( .A(G116), .B(G107), .Z(n554) );
  XNOR2_X1 U617 ( .A(n520), .B(G146), .ZN(n500) );
  XNOR2_X1 U618 ( .A(n489), .B(n488), .ZN(n490) );
  INV_X1 U619 ( .A(KEYINPUT80), .ZN(n597) );
  XNOR2_X1 U620 ( .A(n491), .B(n490), .ZN(n493) );
  INV_X1 U621 ( .A(KEYINPUT35), .ZN(n618) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n518) );
  NOR2_X1 U623 ( .A1(G952), .A2(n753), .ZN(n728) );
  XNOR2_X1 U624 ( .A(G113), .B(G122), .ZN(n486) );
  XNOR2_X1 U625 ( .A(n486), .B(G104), .ZN(n536) );
  NAND2_X1 U626 ( .A1(G214), .A2(n505), .ZN(n489) );
  XOR2_X1 U627 ( .A(KEYINPUT66), .B(G131), .Z(n499) );
  XNOR2_X1 U628 ( .A(n499), .B(n743), .ZN(n492) );
  XNOR2_X1 U629 ( .A(n493), .B(n492), .ZN(n548) );
  NAND2_X1 U630 ( .A1(G214), .A2(n544), .ZN(n698) );
  XOR2_X1 U631 ( .A(KEYINPUT94), .B(G113), .Z(n502) );
  XNOR2_X1 U632 ( .A(G137), .B(G116), .ZN(n501) );
  XNOR2_X1 U633 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U634 ( .A(G119), .B(KEYINPUT69), .ZN(n504) );
  NAND2_X1 U635 ( .A1(n505), .A2(G210), .ZN(n506) );
  INV_X1 U636 ( .A(KEYINPUT30), .ZN(n507) );
  XNOR2_X1 U637 ( .A(n508), .B(n507), .ZN(n533) );
  NAND2_X1 U638 ( .A1(n513), .A2(G221), .ZN(n509) );
  XNOR2_X1 U639 ( .A(n509), .B(KEYINPUT21), .ZN(n680) );
  NAND2_X1 U640 ( .A1(n753), .A2(G234), .ZN(n511) );
  XNOR2_X1 U641 ( .A(KEYINPUT65), .B(KEYINPUT8), .ZN(n510) );
  NOR2_X1 U642 ( .A1(n726), .A2(G902), .ZN(n519) );
  NAND2_X1 U643 ( .A1(n513), .A2(G217), .ZN(n514) );
  XNOR2_X1 U644 ( .A(KEYINPUT91), .B(KEYINPUT25), .ZN(n516) );
  XNOR2_X1 U645 ( .A(n527), .B(KEYINPUT88), .ZN(n528) );
  XNOR2_X1 U646 ( .A(KEYINPUT14), .B(n528), .ZN(n529) );
  NAND2_X1 U647 ( .A1(G952), .A2(n529), .ZN(n710) );
  NOR2_X1 U648 ( .A1(G953), .A2(n710), .ZN(n601) );
  NAND2_X1 U649 ( .A1(G902), .A2(n529), .ZN(n599) );
  OR2_X1 U650 ( .A1(n753), .A2(n599), .ZN(n530) );
  NOR2_X1 U651 ( .A1(G900), .A2(n530), .ZN(n531) );
  NOR2_X1 U652 ( .A1(n601), .A2(n531), .ZN(n562) );
  XOR2_X1 U653 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n535) );
  XNOR2_X1 U654 ( .A(n554), .B(n535), .ZN(n537) );
  NAND2_X1 U655 ( .A1(G224), .A2(n753), .ZN(n540) );
  XNOR2_X1 U656 ( .A(n541), .B(n540), .ZN(n542) );
  NAND2_X1 U657 ( .A1(n646), .A2(n543), .ZN(n545) );
  XOR2_X1 U658 ( .A(KEYINPUT38), .B(n585), .Z(n569) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n546) );
  XNOR2_X1 U660 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n549) );
  INV_X1 U661 ( .A(n572), .ZN(n576) );
  XNOR2_X1 U662 ( .A(n553), .B(n552), .ZN(n557) );
  XOR2_X1 U663 ( .A(n554), .B(KEYINPUT9), .Z(n556) );
  XOR2_X1 U664 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n561) );
  XOR2_X1 U665 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n567) );
  XNOR2_X1 U666 ( .A(KEYINPUT68), .B(n563), .ZN(n564) );
  NAND2_X1 U667 ( .A1(n564), .A2(n679), .ZN(n565) );
  XNOR2_X1 U668 ( .A(n565), .B(KEYINPUT67), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n608), .A2(n583), .ZN(n566) );
  XOR2_X1 U670 ( .A(n567), .B(n566), .Z(n568) );
  NOR2_X1 U671 ( .A1(n575), .A2(n572), .ZN(n701) );
  INV_X1 U672 ( .A(n701), .ZN(n605) );
  INV_X1 U673 ( .A(n569), .ZN(n699) );
  NAND2_X1 U674 ( .A1(n699), .A2(n698), .ZN(n695) );
  NAND2_X1 U675 ( .A1(n579), .A2(n716), .ZN(n570) );
  XNOR2_X1 U676 ( .A(n570), .B(KEYINPUT42), .ZN(n761) );
  NAND2_X1 U677 ( .A1(n575), .A2(n572), .ZN(n617) );
  OR2_X1 U678 ( .A1(n617), .A2(n585), .ZN(n573) );
  NOR2_X1 U679 ( .A1(n574), .A2(n573), .ZN(n666) );
  NOR2_X1 U680 ( .A1(n594), .A2(n655), .ZN(n577) );
  INV_X1 U681 ( .A(n603), .ZN(n580) );
  NAND2_X1 U682 ( .A1(n580), .A2(n579), .ZN(n667) );
  XOR2_X1 U683 ( .A(n581), .B(KEYINPUT47), .Z(n589) );
  XNOR2_X1 U684 ( .A(KEYINPUT6), .B(n688), .ZN(n598) );
  NAND2_X1 U685 ( .A1(n584), .A2(n698), .ZN(n591) );
  XNOR2_X1 U686 ( .A(n586), .B(KEYINPUT36), .ZN(n587) );
  XNOR2_X1 U687 ( .A(n587), .B(KEYINPUT108), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n589), .A2(n675), .ZN(n590) );
  NOR2_X1 U689 ( .A1(n609), .A2(n591), .ZN(n592) );
  XNOR2_X1 U690 ( .A(n592), .B(KEYINPUT43), .ZN(n593) );
  NAND2_X1 U691 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U692 ( .A(KEYINPUT109), .B(n596), .Z(n756) );
  INV_X1 U693 ( .A(KEYINPUT44), .ZN(n622) );
  NAND2_X1 U694 ( .A1(n622), .A2(KEYINPUT84), .ZN(n613) );
  INV_X1 U695 ( .A(n598), .ZN(n614) );
  XNOR2_X1 U696 ( .A(G898), .B(KEYINPUT89), .ZN(n731) );
  NAND2_X1 U697 ( .A1(G953), .A2(n731), .ZN(n738) );
  NOR2_X1 U698 ( .A1(n738), .A2(n599), .ZN(n600) );
  NOR2_X1 U699 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U700 ( .A1(n680), .A2(n605), .ZN(n606) );
  INV_X1 U701 ( .A(n679), .ZN(n636) );
  OR2_X1 U702 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U703 ( .A1(n611), .A2(n610), .ZN(n612) );
  NAND2_X1 U704 ( .A1(n612), .A2(n679), .ZN(n663) );
  XOR2_X1 U705 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n616) );
  NOR2_X1 U706 ( .A1(n683), .A2(n684), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n621), .A2(n627), .ZN(n624) );
  INV_X1 U708 ( .A(n627), .ZN(n757) );
  NAND2_X1 U709 ( .A1(n622), .A2(n757), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n626) );
  INV_X1 U711 ( .A(KEYINPUT64), .ZN(n625) );
  NOR2_X1 U712 ( .A1(n626), .A2(n625), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n629), .A2(n630), .ZN(n659) );
  INV_X1 U714 ( .A(n630), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n688), .A2(n631), .ZN(n692) );
  NOR2_X1 U716 ( .A1(n632), .A2(n692), .ZN(n633) );
  XNOR2_X1 U717 ( .A(n633), .B(KEYINPUT31), .ZN(n671) );
  NAND2_X1 U718 ( .A1(n659), .A2(n671), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n683), .ZN(n638) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(n352), .ZN(n637) );
  NOR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n653) );
  XNOR2_X1 U722 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n646), .B(KEYINPUT54), .ZN(n647) );
  XOR2_X1 U724 ( .A(n650), .B(KEYINPUT62), .Z(n651) );
  XNOR2_X1 U725 ( .A(G101), .B(n653), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(KEYINPUT111), .ZN(G3) );
  INV_X1 U727 ( .A(n655), .ZN(n669) );
  NOR2_X1 U728 ( .A1(n669), .A2(n659), .ZN(n656) );
  XOR2_X1 U729 ( .A(G104), .B(n656), .Z(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n658) );
  XNOR2_X1 U731 ( .A(G107), .B(KEYINPUT112), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n661) );
  NOR2_X1 U733 ( .A1(n672), .A2(n659), .ZN(n660) );
  XOR2_X1 U734 ( .A(n661), .B(n660), .Z(G9) );
  XOR2_X1 U735 ( .A(G110), .B(KEYINPUT113), .Z(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(G12) );
  NOR2_X1 U737 ( .A1(n672), .A2(n667), .ZN(n665) );
  XNOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(G30) );
  XOR2_X1 U740 ( .A(G143), .B(n666), .Z(G45) );
  NOR2_X1 U741 ( .A1(n669), .A2(n667), .ZN(n668) );
  XOR2_X1 U742 ( .A(G146), .B(n668), .Z(G48) );
  NOR2_X1 U743 ( .A1(n669), .A2(n671), .ZN(n670) );
  XOR2_X1 U744 ( .A(G113), .B(n670), .Z(G15) );
  NOR2_X1 U745 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U746 ( .A(KEYINPUT114), .B(n673), .Z(n674) );
  XNOR2_X1 U747 ( .A(G116), .B(n674), .ZN(G18) );
  XNOR2_X1 U748 ( .A(n675), .B(G125), .ZN(n676) );
  XNOR2_X1 U749 ( .A(n676), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U750 ( .A(G140), .B(n677), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n678), .B(KEYINPUT115), .ZN(G42) );
  XOR2_X1 U752 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n682) );
  NAND2_X1 U753 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n682), .B(n681), .ZN(n690) );
  NAND2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  XNOR2_X1 U757 ( .A(KEYINPUT117), .B(n686), .ZN(n687) );
  NOR2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U761 ( .A(KEYINPUT51), .B(n693), .Z(n694) );
  NAND2_X1 U762 ( .A1(n716), .A2(n694), .ZN(n707) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U764 ( .A(n697), .B(KEYINPUT119), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U766 ( .A(KEYINPUT118), .B(n700), .Z(n702) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U769 ( .A1(n717), .A2(n705), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U771 ( .A(KEYINPUT52), .B(n708), .Z(n709) );
  NOR2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n715) );
  INV_X1 U773 ( .A(n732), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n720) );
  XOR2_X1 U776 ( .A(n721), .B(KEYINPUT123), .Z(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n728), .A2(n724), .ZN(G63) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n728), .A2(n727), .ZN(G66) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n729) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(n729), .Z(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U784 ( .A1(G953), .A2(n732), .ZN(n733) );
  NOR2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n740) );
  XOR2_X1 U786 ( .A(G101), .B(n735), .Z(n736) );
  XNOR2_X1 U787 ( .A(G110), .B(n736), .ZN(n737) );
  NAND2_X1 U788 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(KEYINPUT124), .B(n741), .ZN(G69) );
  XNOR2_X1 U791 ( .A(n743), .B(n742), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n745), .B(n744), .ZN(n749) );
  XNOR2_X1 U793 ( .A(G227), .B(n749), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n747), .B(KEYINPUT126), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n755) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT125), .ZN(n751) );
  XNOR2_X1 U798 ( .A(n751), .B(n750), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U801 ( .A(G134), .B(n756), .ZN(G36) );
  XNOR2_X1 U802 ( .A(G122), .B(n757), .ZN(n758) );
  XNOR2_X1 U803 ( .A(n758), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U804 ( .A(n759), .B(G119), .ZN(G21) );
  XNOR2_X1 U805 ( .A(n354), .B(G131), .ZN(G33) );
  XNOR2_X1 U806 ( .A(n761), .B(G137), .ZN(G39) );
endmodule

