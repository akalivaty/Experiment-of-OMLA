//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT66), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n220));
  AND3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT65), .Z(new_n223));
  AOI21_X1  g0023(.A(new_n209), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n208), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n215), .B1(new_n216), .B2(new_n224), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n224), .A2(new_n216), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT67), .Z(new_n231));
  NOR2_X1   g0031(.A1(new_n229), .A2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n236), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G222), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G223), .A2(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n254), .B(new_n255), .C1(G77), .C2(new_n250), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G274), .ZN(new_n262));
  INV_X1    g0062(.A(G226), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n256), .B(new_n262), .C1(new_n263), .C2(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(G179), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n225), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n208), .A2(G1), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n201), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G50), .B2(new_n268), .ZN(new_n276));
  INV_X1    g0076(.A(new_n271), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT8), .B(G58), .Z(new_n278));
  NAND2_X1  g0078(.A1(new_n208), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT70), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT70), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(new_n208), .A3(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n278), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n277), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n266), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n267), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G238), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G232), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n250), .B(new_n292), .C1(new_n293), .C2(G1698), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n294), .B(new_n255), .C1(G107), .C2(new_n250), .ZN(new_n295));
  INV_X1    g0095(.A(new_n265), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G244), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n295), .A2(new_n262), .A3(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(G169), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n273), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n272), .A2(new_n301), .B1(new_n300), .B2(new_n269), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G20), .A2(G77), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(new_n279), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n284), .B2(new_n278), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n302), .B1(new_n306), .B2(new_n277), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n299), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n298), .B2(G190), .ZN(new_n311));
  INV_X1    g0111(.A(G200), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n298), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g0114(.A(new_n287), .B(KEYINPUT9), .Z(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n266), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(G200), .B2(new_n266), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n291), .B(new_n314), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT71), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n319), .B(KEYINPUT10), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT71), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n291), .A4(new_n314), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT75), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT73), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT12), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n331), .C1(new_n268), .C2(G68), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT74), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n268), .A2(KEYINPUT12), .A3(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(KEYINPUT74), .B2(new_n332), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n280), .A2(G77), .A3(new_n282), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n277), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n272), .B(G68), .C1(G1), .C2(new_n208), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n339), .B2(KEYINPUT11), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n327), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n333), .A2(new_n335), .B1(new_n339), .B2(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(new_n341), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT75), .A4(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n293), .A2(G1698), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n250), .B(new_n350), .C1(G226), .C2(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n255), .ZN(new_n354));
  INV_X1    g0154(.A(G238), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n262), .B1(new_n355), .B2(new_n265), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n261), .B1(new_n351), .B2(new_n352), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT13), .B1(new_n360), .B2(new_n356), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G190), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n362), .A2(KEYINPUT72), .A3(new_n312), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n359), .A2(new_n361), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(G200), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n349), .B(new_n363), .C1(new_n364), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n349), .B(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n289), .B1(new_n359), .B2(new_n361), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT14), .ZN(new_n372));
  AOI22_X1  g0172(.A1(G179), .A2(new_n362), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT76), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n366), .A2(new_n372), .A3(G169), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n359), .A2(G179), .A3(new_n361), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT76), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n379), .A2(new_n380), .A3(new_n374), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n370), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n323), .A2(new_n326), .A3(new_n368), .A4(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  OR2_X1    g0184(.A1(KEYINPUT3), .A2(G33), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n208), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n386), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n203), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n202), .A2(new_n203), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n284), .A2(G159), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n384), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g0197(.A1(KEYINPUT3), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(KEYINPUT3), .A2(G33), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n400), .B2(new_n208), .ZN(new_n401));
  NOR4_X1   g0201(.A1(new_n398), .A2(new_n399), .A3(new_n388), .A4(G20), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n396), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(KEYINPUT16), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n405), .A3(new_n271), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT8), .B(G58), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n273), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n272), .B1(new_n269), .B2(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n263), .A2(G1698), .ZN(new_n410));
  OAI221_X1 g0210(.A(new_n410), .B1(G223), .B2(G1698), .C1(new_n398), .C2(new_n399), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n255), .ZN(new_n414));
  INV_X1    g0214(.A(G274), .ZN(new_n415));
  INV_X1    g0215(.A(new_n225), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n415), .B1(new_n416), .B2(new_n260), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n296), .A2(G232), .B1(new_n259), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n316), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n261), .B1(new_n411), .B2(new_n412), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n262), .B1(new_n293), .B2(new_n265), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n312), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n406), .A2(new_n409), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT17), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n406), .A2(new_n423), .A3(new_n426), .A4(new_n409), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT78), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n414), .A2(new_n308), .A3(new_n418), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n289), .B1(new_n420), .B2(new_n421), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n406), .B2(new_n409), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n425), .A2(KEYINPUT78), .A3(new_n427), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n430), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n383), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n250), .A2(new_n208), .A3(G87), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G116), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G20), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n208), .B2(G107), .ZN(new_n444));
  INV_X1    g0244(.A(G107), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(KEYINPUT23), .A3(G20), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G87), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT24), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n250), .A2(new_n208), .A3(G87), .ZN(new_n453));
  INV_X1    g0253(.A(new_n449), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT24), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n440), .A3(new_n447), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n271), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n207), .A2(G33), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n268), .A2(new_n460), .A3(new_n225), .A4(new_n270), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n269), .A2(KEYINPUT25), .A3(new_n445), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT25), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n268), .B2(G107), .ZN(new_n465));
  AOI22_X1  g0265(.A1(G107), .A2(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT86), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n258), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n257), .A2(KEYINPUT5), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT5), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n473), .A2(new_n255), .A3(new_n415), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(G257), .A2(G1698), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n477), .B1(new_n250), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G250), .B(new_n251), .C1(new_n398), .C2(new_n399), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n261), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(G264), .A3(new_n261), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n478), .B1(new_n398), .B2(new_n399), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n255), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n308), .B(new_n474), .C1(new_n484), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n474), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n490), .A3(new_n482), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(G169), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n468), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n491), .A2(G190), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n481), .A2(new_n475), .A3(new_n483), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT87), .B1(new_n487), .B2(new_n482), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(new_n312), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT88), .B1(new_n499), .B2(new_n467), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n474), .B1(new_n484), .B2(new_n488), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(G200), .B1(new_n491), .B2(G190), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT88), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n459), .A4(new_n466), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n207), .B(G45), .C1(new_n257), .C2(KEYINPUT5), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n471), .A2(G41), .ZN(new_n508));
  OAI211_X1 g0308(.A(G270), .B(new_n261), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT84), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n473), .A2(new_n511), .A3(G270), .A4(new_n261), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G303), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n261), .B1(new_n400), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n251), .A2(G257), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G264), .A2(G1698), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n250), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n507), .A2(new_n508), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n515), .A2(new_n518), .B1(new_n417), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n289), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n269), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n461), .B2(new_n522), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n270), .A2(new_n225), .B1(G20), .B2(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G283), .ZN(new_n526));
  INV_X1    g0326(.A(G97), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n208), .C1(G33), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(KEYINPUT20), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n525), .A2(new_n528), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n524), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT21), .B1(new_n521), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n513), .A2(G179), .A3(new_n520), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n533), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n521), .A2(new_n534), .A3(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n513), .A2(new_n520), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G200), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n533), .C1(new_n316), .C2(new_n540), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(G244), .C1(new_n399), .C2(new_n398), .ZN(new_n546));
  INV_X1    g0346(.A(G244), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n385), .B2(new_n386), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n526), .C1(new_n548), .C2(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n250), .A2(G250), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n251), .B1(new_n550), .B2(KEYINPUT4), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n255), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(G257), .B(new_n261), .C1(new_n507), .C2(new_n508), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT79), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n473), .A2(KEYINPUT79), .A3(G257), .A4(new_n261), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n474), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n284), .A2(G77), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n561), .A2(new_n527), .A3(G107), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n562), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n208), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n445), .B1(new_n389), .B2(new_n390), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n271), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n268), .A2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n462), .B2(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n552), .A2(new_n557), .A3(G190), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n559), .A2(new_n567), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n558), .A2(new_n289), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n552), .A2(new_n557), .A3(new_n308), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n567), .A2(new_n569), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n258), .B2(G1), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n207), .A2(new_n415), .A3(G45), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n261), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G238), .A2(G1698), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n547), .B2(G1698), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n250), .B1(G33), .B2(G116), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n316), .B(new_n579), .C1(new_n582), .C2(new_n261), .ZN(new_n583));
  INV_X1    g0383(.A(new_n579), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n547), .A2(G1698), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G238), .B2(G1698), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n441), .B1(new_n586), .B2(new_n400), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n587), .B2(new_n255), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n583), .B1(new_n588), .B2(G200), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT83), .ZN(new_n590));
  NAND3_X1  g0390(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT82), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n591), .A2(new_n592), .A3(new_n208), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n592), .B1(new_n591), .B2(new_n208), .ZN(new_n594));
  NOR3_X1   g0394(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n208), .B(G68), .C1(new_n398), .C2(new_n399), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT19), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n279), .B2(new_n527), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n590), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n591), .A2(new_n208), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n591), .A2(new_n592), .A3(new_n208), .ZN(new_n604));
  INV_X1    g0404(.A(new_n595), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT83), .A3(new_n597), .A4(new_n599), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n601), .A2(new_n271), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n462), .A2(G87), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n304), .A2(new_n269), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n589), .A2(new_n608), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n571), .A2(new_n575), .A3(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n308), .B(new_n579), .C1(new_n582), .C2(new_n261), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT80), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n588), .A2(new_n615), .A3(new_n308), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n579), .B1(new_n582), .B2(new_n261), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n289), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT81), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT81), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n614), .A2(new_n616), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n608), .A2(new_n610), .ZN(new_n623));
  INV_X1    g0423(.A(new_n304), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n462), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n620), .A2(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n543), .A2(new_n612), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n438), .A2(new_n506), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n291), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT76), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n380), .B1(new_n379), .B2(new_n374), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n310), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n632), .A2(new_n370), .B1(new_n368), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n436), .B(new_n430), .C1(new_n634), .C2(KEYINPUT90), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(KEYINPUT90), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n435), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n629), .B1(new_n637), .B2(new_n324), .ZN(new_n638));
  INV_X1    g0438(.A(new_n438), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n608), .A2(new_n610), .A3(new_n625), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n618), .A2(new_n613), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n521), .A2(new_n534), .A3(KEYINPUT21), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n644), .A2(new_n535), .A3(new_n537), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n467), .B1(new_n489), .B2(new_n492), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n612), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n505), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n589), .B1(new_n640), .B2(new_n641), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n558), .A2(new_n289), .B1(new_n567), .B2(new_n569), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n653), .A2(KEYINPUT89), .A3(new_n573), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT89), .B1(new_n653), .B2(new_n573), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n650), .B(new_n652), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n653), .A2(new_n611), .A3(new_n573), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT26), .B1(new_n626), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n656), .A2(new_n658), .A3(new_n642), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n638), .B1(new_n639), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT91), .Z(G369));
  NAND3_X1  g0462(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT92), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT27), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(G213), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n494), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n670), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n468), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n506), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n645), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n534), .A3(new_n672), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n645), .B(new_n542), .C1(new_n533), .C2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT93), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT93), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n681), .A3(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G330), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n683), .B2(G330), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n675), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n646), .A2(new_n672), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n645), .A2(new_n672), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n506), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(G399));
  NOR2_X1   g0492(.A1(new_n211), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n605), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n228), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n642), .A2(new_n611), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n575), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n653), .A2(KEYINPUT89), .A3(new_n573), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n643), .B1(new_n703), .B2(new_n650), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n505), .A2(new_n647), .A3(new_n648), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n658), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n670), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(KEYINPUT29), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n494), .A2(new_n645), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n612), .B1(new_n500), .B2(new_n504), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n643), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n650), .B1(new_n626), .B2(new_n657), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT96), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n703), .A2(KEYINPUT26), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n650), .C1(new_n626), .C2(new_n657), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n709), .B1(new_n719), .B2(new_n670), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n558), .A2(new_n308), .A3(new_n540), .A4(new_n617), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n501), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n558), .A2(new_n617), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n484), .A2(new_n488), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n722), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n724), .A4(new_n723), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n670), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n627), .A2(new_n494), .A3(new_n505), .A4(new_n670), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n708), .B(new_n720), .C1(G330), .C2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n698), .B1(new_n737), .B2(G1), .ZN(G364));
  NOR2_X1   g0538(.A1(new_n686), .A2(new_n687), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n210), .A2(G20), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n694), .A2(G1), .A3(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n739), .B(new_n742), .C1(G330), .C2(new_n683), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n225), .B1(G20), .B2(new_n289), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n248), .A2(new_n258), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT98), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n211), .A2(new_n250), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n228), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n258), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n750), .B1(new_n751), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n751), .B2(new_n755), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n212), .A2(new_n250), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(KEYINPUT97), .B2(G355), .ZN(new_n759));
  OR2_X1    g0559(.A1(G355), .A2(KEYINPUT97), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n759), .A2(new_n760), .B1(new_n522), .B2(new_n211), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n749), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n747), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n208), .A2(new_n316), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n312), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G87), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n308), .A2(G200), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n208), .A2(G190), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n770), .B2(new_n300), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n765), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n400), .B(new_n771), .C1(G107), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G179), .A2(G200), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n208), .B1(new_n775), .B2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n527), .ZN(new_n777));
  NAND3_X1  g0577(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n316), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n201), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(G190), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n777), .B(new_n781), .C1(G68), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n769), .A2(new_n775), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n764), .A2(new_n768), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT99), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G58), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n774), .A2(new_n783), .A3(new_n787), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G322), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n400), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G326), .B2(new_n779), .ZN(new_n795));
  INV_X1    g0595(.A(new_n770), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G283), .A2(new_n773), .B1(new_n796), .B2(G311), .ZN(new_n797));
  INV_X1    g0597(.A(new_n766), .ZN(new_n798));
  INV_X1    g0598(.A(new_n784), .ZN(new_n799));
  AOI22_X1  g0599(.A1(G303), .A2(new_n798), .B1(new_n799), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(new_n776), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n801), .A2(G294), .B1(new_n782), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n795), .A2(new_n797), .A3(new_n800), .A4(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n763), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n762), .A2(new_n805), .A3(new_n742), .ZN(new_n806));
  INV_X1    g0606(.A(new_n746), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n683), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n743), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NOR2_X1   g0610(.A1(new_n747), .A2(new_n744), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n742), .B1(new_n300), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G87), .A2(new_n773), .B1(new_n799), .B2(G311), .ZN(new_n813));
  INV_X1    g0613(.A(G294), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n522), .B2(new_n770), .C1(new_n814), .C2(new_n788), .ZN(new_n815));
  INV_X1    g0615(.A(new_n782), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n816), .A2(new_n817), .B1(new_n780), .B2(new_n514), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n400), .B1(new_n766), .B2(new_n445), .ZN(new_n819));
  NOR4_X1   g0619(.A1(new_n815), .A2(new_n777), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n796), .A2(G159), .B1(G150), .B2(new_n782), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n780), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G143), .B2(new_n790), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G50), .A2(new_n798), .B1(new_n799), .B2(G132), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n400), .B1(new_n773), .B2(G68), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(new_n202), .C2(new_n776), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(new_n824), .B2(KEYINPUT34), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n820), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n672), .A2(new_n307), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n633), .B1(new_n313), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n633), .A2(new_n670), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n812), .B1(new_n763), .B2(new_n830), .C1(new_n836), .C2(new_n745), .ZN(new_n837));
  INV_X1    g0637(.A(new_n742), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n314), .A2(new_n670), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n660), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n840), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n706), .A2(KEYINPUT100), .A3(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n841), .A2(new_n843), .B1(new_n707), .B2(new_n835), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n736), .A2(G330), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(G384));
  INV_X1    g0650(.A(KEYINPUT35), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n564), .A2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n522), .B(new_n227), .C1(new_n564), .C2(new_n851), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n852), .B1(new_n854), .B2(KEYINPUT101), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(KEYINPUT101), .B2(new_n854), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g0657(.A(new_n754), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n201), .A2(G68), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n207), .B(G13), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n435), .A2(new_n669), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n370), .A2(new_n672), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n382), .A2(new_n368), .A3(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n368), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n370), .B(new_n672), .C1(new_n632), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n841), .A2(new_n843), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n869), .B2(new_n834), .ZN(new_n870));
  INV_X1    g0670(.A(new_n409), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n403), .A2(new_n404), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n277), .B1(new_n872), .B2(new_n384), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n405), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n874), .A2(new_n668), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n424), .B1(new_n874), .B2(new_n433), .ZN(new_n876));
  OAI21_X1  g0676(.A(KEYINPUT37), .B1(new_n876), .B2(new_n875), .ZN(new_n877));
  INV_X1    g0677(.A(new_n434), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n406), .A2(new_n409), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n669), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT37), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n424), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n437), .A2(new_n875), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n883), .A2(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n437), .A2(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n882), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n862), .B1(new_n870), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT104), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n883), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT18), .B1(new_n874), .B2(new_n433), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT18), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n434), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n428), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n875), .A2(new_n898), .B1(new_n877), .B2(new_n882), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n894), .B1(new_n899), .B2(KEYINPUT38), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n877), .A2(new_n882), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n880), .B1(new_n435), .B2(new_n428), .ZN(new_n903));
  OAI211_X1 g0703(.A(KEYINPUT102), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n892), .A2(new_n893), .A3(new_n900), .A4(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n382), .A2(new_n672), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n889), .A2(new_n890), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n890), .B1(new_n889), .B2(new_n910), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n438), .B1(new_n720), .B2(new_n708), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n638), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n914), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT31), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT105), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n918), .B1(new_n732), .B2(new_n919), .ZN(new_n920));
  AOI211_X1 g0720(.A(KEYINPUT105), .B(new_n670), .C1(new_n729), .C2(new_n731), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n734), .B(new_n735), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n835), .B1(new_n864), .B2(new_n866), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n905), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n883), .A2(KEYINPUT38), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n885), .A2(KEYINPUT38), .A3(new_n886), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n922), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT40), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n925), .A2(new_n930), .A3(new_n438), .A4(new_n922), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(G330), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n925), .A2(new_n930), .B1(new_n438), .B2(new_n922), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n917), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n207), .B2(new_n740), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n917), .A2(new_n934), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n861), .B1(new_n936), .B2(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n688), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n672), .A2(new_n574), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n940), .A2(new_n575), .A3(new_n571), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n672), .A2(new_n573), .A3(new_n653), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n691), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT45), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT44), .B1(new_n691), .B2(new_n943), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n939), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT45), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n944), .B(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n951), .A2(new_n688), .A3(new_n947), .A4(new_n946), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n506), .A2(new_n690), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n674), .B1(new_n645), .B2(new_n672), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n739), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n954), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n686), .B2(new_n687), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n737), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n693), .B(KEYINPUT41), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n741), .A2(G1), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT106), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n506), .A2(new_n690), .A3(new_n943), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(KEYINPUT42), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n575), .B1(new_n494), .B2(new_n941), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(KEYINPUT42), .B1(new_n670), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n652), .B1(new_n651), .B2(new_n670), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n642), .A2(new_n651), .A3(new_n670), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n969), .A2(new_n971), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n976), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n943), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n688), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n967), .A2(new_n982), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n772), .A2(new_n300), .B1(new_n784), .B2(new_n822), .ZN(new_n984));
  INV_X1    g0784(.A(G150), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n250), .B1(new_n776), .B2(new_n203), .C1(new_n985), .C2(new_n788), .ZN(new_n986));
  INV_X1    g0786(.A(G143), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n816), .A2(new_n785), .B1(new_n780), .B2(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n766), .A2(new_n202), .B1(new_n770), .B2(new_n201), .ZN(new_n989));
  OR4_X1    g0789(.A1(new_n984), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n772), .A2(new_n527), .B1(new_n784), .B2(new_n991), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n250), .B(new_n992), .C1(G283), .C2(new_n796), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n798), .A2(G116), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n994), .A2(new_n995), .B1(new_n779), .B2(G311), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n993), .B(new_n996), .C1(new_n514), .C2(new_n789), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n782), .A2(G294), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n445), .B2(new_n776), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n990), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT107), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n747), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n972), .A2(new_n746), .A3(new_n973), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n236), .A2(new_n753), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n749), .B1(new_n211), .B2(new_n624), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n742), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n983), .A2(new_n1008), .ZN(G387));
  NAND2_X1  g0809(.A1(new_n278), .A2(new_n201), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n695), .B(new_n258), .C1(new_n203), .C2(new_n300), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n752), .B1(new_n1011), .B2(new_n1012), .C1(new_n240), .C2(new_n258), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1013), .B1(G107), .B2(new_n212), .C1(new_n695), .C2(new_n758), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n742), .B1(new_n1014), .B2(new_n748), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n801), .A2(new_n624), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n780), .B2(new_n785), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n250), .B1(new_n772), .B2(new_n527), .C1(new_n816), .C2(new_n407), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n766), .A2(new_n300), .B1(new_n784), .B2(new_n985), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n788), .A2(new_n201), .B1(new_n770), .B2(new_n203), .ZN(new_n1020));
  NOR4_X1   g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n796), .A2(G303), .B1(G311), .B2(new_n782), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n793), .B2(new_n780), .C1(new_n789), .C2(new_n991), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT48), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n798), .A2(G294), .B1(new_n801), .B2(G283), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n250), .B1(new_n799), .B2(G326), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n522), .B2(new_n772), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n1029), .B2(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1021), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1015), .B1(new_n763), .B2(new_n1034), .C1(new_n675), .C2(new_n807), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n959), .A2(new_n737), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n693), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n959), .A2(new_n737), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1035), .B1(new_n960), .B2(new_n966), .C1(new_n1037), .C2(new_n1038), .ZN(G393));
  OR2_X1    g0839(.A1(new_n953), .A2(new_n1036), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n953), .A2(new_n1036), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n693), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT108), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n953), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n966), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT108), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT110), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n980), .A2(new_n746), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n245), .A2(new_n753), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n748), .B1(new_n527), .B2(new_n212), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n838), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n780), .A2(new_n985), .B1(new_n788), .B2(new_n785), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT51), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n776), .A2(new_n300), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n250), .B1(new_n772), .B2(new_n767), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(G50), .C2(new_n782), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n770), .A2(new_n407), .B1(new_n784), .B2(new_n987), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G68), .B2(new_n798), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n788), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1062), .A2(G311), .B1(G317), .B2(new_n779), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n770), .A2(new_n814), .B1(new_n784), .B2(new_n793), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G283), .B2(new_n798), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n400), .B1(new_n772), .B2(new_n445), .C1(new_n816), .C2(new_n514), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G116), .B2(new_n801), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1061), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1071), .B2(new_n747), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1049), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1047), .A2(new_n1048), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1048), .B1(new_n1047), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1042), .B1(new_n1075), .B2(new_n1076), .ZN(G390));
  NAND3_X1  g0877(.A1(new_n438), .A2(G330), .A3(new_n922), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n915), .A2(new_n638), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n922), .A2(G330), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n836), .B1(new_n1080), .B2(KEYINPUT113), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT113), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n922), .B2(G330), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n868), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n736), .A2(new_n867), .A3(G330), .A4(new_n836), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n834), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n672), .B(new_n832), .C1(new_n712), .C2(new_n718), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT112), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n923), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1091), .B1(new_n1080), .B2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT112), .A4(G330), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n868), .B1(new_n846), .B2(new_n835), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n656), .A2(new_n658), .A3(new_n642), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n839), .B(new_n840), .C1(new_n1097), .C2(new_n705), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT100), .B1(new_n706), .B2(new_n842), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n834), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1079), .B1(new_n1090), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n867), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n909), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n905), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1087), .B1(new_n841), .B2(new_n843), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1108), .B2(new_n868), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1109), .A2(KEYINPUT111), .B1(new_n907), .B2(new_n908), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n909), .B1(new_n1100), .B2(new_n867), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1107), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n900), .A2(new_n904), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT103), .B1(new_n883), .B2(KEYINPUT38), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n1119), .B2(new_n893), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n908), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1111), .A2(new_n1112), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n870), .A2(KEYINPUT111), .A3(new_n909), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1106), .B(new_n1085), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1103), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1124), .B(new_n1102), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n693), .A3(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1045), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n811), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(G116), .A2(new_n1062), .B1(new_n799), .B2(G294), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n203), .B2(new_n772), .C1(new_n527), .C2(new_n770), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n816), .A2(new_n445), .B1(new_n780), .B2(new_n817), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n400), .B1(new_n766), .B2(new_n767), .ZN(new_n1134));
  NOR4_X1   g0934(.A1(new_n1132), .A2(new_n1055), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT114), .Z(new_n1136));
  OAI21_X1  g0936(.A(new_n250), .B1(new_n772), .B2(new_n201), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G128), .B2(new_n779), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n801), .A2(G159), .B1(G137), .B2(new_n782), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n766), .A2(new_n985), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT53), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n796), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G132), .A2(new_n1062), .B1(new_n799), .B2(G125), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1140), .A2(new_n1142), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1136), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1149), .A2(KEYINPUT115), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n747), .B1(new_n1149), .B2(KEYINPUT115), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n838), .B1(new_n278), .B2(new_n1130), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n907), .A2(new_n908), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n744), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1128), .A2(new_n1129), .A3(new_n1155), .ZN(G378));
  OAI21_X1  g0956(.A(new_n838), .B1(G50), .B2(new_n1130), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n201), .B1(G33), .B2(G41), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n400), .B2(new_n257), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G41), .B(new_n250), .C1(new_n798), .C2(G77), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n202), .B2(new_n772), .C1(new_n817), .C2(new_n784), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT116), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n788), .A2(new_n445), .B1(new_n770), .B2(new_n304), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G68), .B2(new_n801), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G97), .A2(new_n782), .B1(new_n779), .B2(G116), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT58), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1159), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n801), .A2(G150), .B1(G125), .B2(new_n779), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT117), .Z(new_n1170));
  NAND2_X1  g0970(.A1(new_n782), .A2(G132), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n796), .A2(G137), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1144), .A2(new_n798), .B1(new_n1062), .B2(G128), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n773), .A2(G159), .ZN(new_n1177));
  AOI211_X1 g0977(.A(G33), .B(G41), .C1(new_n799), .C2(G124), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1157), .B1(new_n1180), .B2(new_n747), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT118), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n324), .A2(new_n291), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n668), .A2(new_n287), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1184), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n324), .A2(new_n291), .A3(new_n1187), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1186), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1182), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1186), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1185), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(KEYINPUT118), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1181), .B1(new_n1197), .B2(new_n745), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n925), .A2(new_n930), .A3(G330), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1197), .A2(new_n925), .A3(new_n930), .A4(G330), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n910), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1100), .A2(new_n888), .A3(new_n867), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n435), .B2(new_n669), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT104), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1205), .A2(new_n1209), .A3(new_n911), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n911), .B2(new_n1209), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1200), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1204), .B(new_n1203), .C1(new_n912), .C2(new_n913), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1205), .A2(new_n1209), .A3(new_n911), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(KEYINPUT119), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1212), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1199), .B1(new_n1216), .B2(new_n1045), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1079), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1127), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1127), .A2(new_n1218), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1216), .A2(new_n1219), .B1(new_n1222), .B2(KEYINPUT57), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1223), .B2(new_n694), .ZN(G375));
  NAND2_X1  g1024(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n868), .A2(new_n744), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n779), .A2(G132), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT121), .Z(new_n1228));
  AOI22_X1  g1028(.A1(G159), .A2(new_n798), .B1(new_n799), .B2(G128), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n1229), .B1(new_n985), .B2(new_n770), .C1(new_n789), .C2(new_n822), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n776), .A2(new_n201), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n250), .B1(new_n772), .B2(new_n202), .C1(new_n816), .C2(new_n1143), .ZN(new_n1232));
  OR4_X1    g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n400), .B1(new_n772), .B2(new_n300), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT120), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1016), .B1(new_n780), .B2(new_n814), .C1(new_n522), .C2(new_n816), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n788), .A2(new_n817), .B1(new_n770), .B2(new_n445), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n766), .A2(new_n527), .B1(new_n784), .B2(new_n514), .ZN(new_n1238));
  OR4_X1    g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n763), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n742), .B(new_n1240), .C1(new_n203), .C2(new_n811), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1225), .A2(new_n1045), .B1(new_n1226), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1103), .A2(new_n963), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1225), .A2(new_n1218), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(G381));
  OR2_X1    g1045(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1046), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT108), .B1(new_n949), .B2(new_n952), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1248), .A2(new_n1249), .A3(new_n966), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1073), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT110), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1074), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1008), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n967), .B2(new_n982), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1255), .A3(new_n1042), .ZN(new_n1256));
  OR3_X1    g1056(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1256), .A2(G378), .A3(G381), .A4(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1246), .A2(new_n1247), .A3(new_n1258), .ZN(G407));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G343), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1246), .A2(new_n1260), .A3(new_n1247), .A4(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(G213), .A3(G407), .ZN(G409));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  OAI211_X1 g1065(.A(KEYINPUT123), .B(new_n1103), .C1(new_n1244), .C2(KEYINPUT60), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT123), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1084), .A2(new_n1089), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT60), .B1(new_n1268), .B2(new_n1079), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1267), .B1(new_n1269), .B2(new_n1102), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n694), .B1(new_n1244), .B2(KEYINPUT60), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1266), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1242), .ZN(new_n1273));
  INV_X1    g1073(.A(G384), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1272), .A2(G384), .A3(new_n1242), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1217), .C1(new_n1223), .C2(new_n694), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n962), .B1(new_n1127), .B2(new_n1218), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1216), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1199), .B1(new_n1221), .B2(new_n1045), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1260), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1262), .B(new_n1277), .C1(new_n1278), .C2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT124), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1265), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1278), .A2(new_n1283), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1262), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1262), .A2(G2897), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1277), .B(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1289), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1277), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1287), .A2(new_n1288), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1286), .A2(new_n1292), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT125), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G390), .A2(G387), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(G396), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1298), .A2(new_n1256), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1299), .B1(new_n1298), .B2(new_n1256), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1297), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1299), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(G390), .A2(G387), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1255), .B1(new_n1253), .B2(new_n1042), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1298), .A2(new_n1256), .A3(new_n1299), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(KEYINPUT125), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1302), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1296), .A2(new_n1309), .ZN(new_n1310));
  OR2_X1    g1110(.A1(new_n1284), .A2(KEYINPUT63), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1284), .A2(KEYINPUT63), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .A4(new_n1292), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(G405));
  NOR2_X1   g1115(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1300), .A2(new_n1301), .A3(new_n1297), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1316), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1302), .A2(new_n1308), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1278), .A2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1260), .B2(G375), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(G375), .A2(KEYINPUT126), .A3(new_n1260), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1326), .B1(new_n1327), .B2(new_n1293), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1322), .B(new_n1329), .ZN(G402));
endmodule


