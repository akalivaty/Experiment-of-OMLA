//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1146, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G20), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR3_X1   g0016(.A1(new_n215), .A2(new_n216), .A3(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n211), .A2(new_n213), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  INV_X1    g0020(.A(G116), .ZN(new_n221));
  INV_X1    g0021(.A(G270), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G97), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n223), .B(new_n229), .C1(G58), .C2(G232), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(G1), .B2(G20), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n219), .B(new_n232), .C1(new_n214), .C2(new_n218), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT2), .ZN(new_n236));
  INV_X1    g0036(.A(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n222), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  INV_X1    g0043(.A(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  INV_X1    g0049(.A(G87), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(new_n227), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n209), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n254), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(G232), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n237), .A2(new_n263), .B1(new_n264), .B2(new_n262), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n254), .A2(new_n227), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n256), .A2(new_n268), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n267), .B(new_n270), .C1(new_n226), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT13), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G169), .ZN(new_n274));
  XOR2_X1   g0074(.A(new_n274), .B(KEYINPUT14), .Z(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n208), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n216), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(G77), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n281), .A2(new_n202), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n216), .A2(G68), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n279), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  XOR2_X1   g0087(.A(KEYINPUT70), .B(KEYINPUT11), .Z(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n288), .ZN(new_n290));
  INV_X1    g0090(.A(new_n279), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G1), .B2(new_n216), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G68), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT12), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n293), .A2(G68), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n289), .B(new_n299), .C1(KEYINPUT12), .C2(new_n295), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n277), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n261), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G107), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n261), .A2(G1698), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(new_n305), .B2(new_n226), .C1(G1698), .C2(new_n264), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n257), .ZN(new_n307));
  INV_X1    g0107(.A(G244), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n270), .C1(new_n308), .C2(new_n271), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G20), .A2(G77), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT15), .B(G87), .Z(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n312), .B1(new_n313), .B2(new_n281), .C1(new_n315), .C2(new_n282), .ZN(new_n316));
  INV_X1    g0116(.A(new_n294), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n316), .A2(new_n279), .B1(new_n283), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n283), .B2(new_n292), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n311), .B(new_n319), .C1(G169), .C2(new_n310), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n302), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(KEYINPUT3), .A2(G33), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT71), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT71), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n322), .B1(new_n325), .B2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT7), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n216), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT71), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n254), .ZN(new_n331));
  NAND2_X1  g0131(.A1(KEYINPUT71), .A2(G33), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT3), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(new_n216), .A3(new_n259), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT72), .A2(KEYINPUT7), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n327), .A2(new_n328), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n329), .A2(new_n337), .A3(G68), .ZN(new_n338));
  XNOR2_X1  g0138(.A(G58), .B(G68), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G20), .B1(G159), .B2(new_n280), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT16), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n258), .B1(new_n323), .B2(new_n324), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n343), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n260), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n328), .B1(new_n261), .B2(G20), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n225), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n340), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n341), .A2(new_n279), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n313), .A2(new_n294), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n293), .B2(new_n313), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT73), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n271), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G232), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n254), .A2(new_n250), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G223), .A2(G1698), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n333), .B2(new_n259), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n262), .A2(G226), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n355), .B(new_n270), .C1(new_n361), .C2(new_n256), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G169), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n359), .B(new_n357), .C1(new_n333), .C2(new_n259), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n257), .B1(new_n364), .B2(new_n356), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n365), .A2(G179), .A3(new_n355), .A4(new_n270), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n349), .A2(new_n353), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n365), .A2(new_n371), .A3(new_n355), .A4(new_n270), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n373), .A2(new_n353), .A3(new_n349), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n319), .B1(new_n310), .B2(G190), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n369), .B2(new_n310), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n380));
  INV_X1    g0180(.A(G222), .ZN(new_n381));
  OAI221_X1 g0181(.A(new_n380), .B1(new_n283), .B2(new_n261), .C1(new_n263), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n257), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n354), .A2(G226), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n270), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n317), .A2(new_n202), .ZN(new_n386));
  INV_X1    g0186(.A(G150), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n313), .A2(new_n282), .B1(new_n387), .B2(new_n281), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(G20), .B2(new_n203), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n386), .B1(new_n202), .B2(new_n292), .C1(new_n389), .C2(new_n291), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT9), .ZN(new_n391));
  AOI22_X1  g0191(.A1(G200), .A2(new_n385), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n392), .B1(new_n391), .B2(new_n390), .C1(new_n371), .C2(new_n385), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n385), .A2(G200), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(KEYINPUT69), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n393), .B(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n301), .B1(new_n273), .B2(G200), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n371), .B2(new_n273), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n385), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n276), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n390), .C1(G169), .C2(new_n402), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n398), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n321), .A2(new_n377), .A3(new_n379), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n333), .A2(new_n259), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(G257), .B2(G1698), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n262), .A2(G264), .ZN(new_n411));
  INV_X1    g0211(.A(G303), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n410), .A2(new_n411), .B1(new_n412), .B2(new_n261), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n257), .ZN(new_n414));
  INV_X1    g0214(.A(G45), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(G1), .ZN(new_n416));
  AND2_X1   g0216(.A1(KEYINPUT5), .A2(G41), .ZN(new_n417));
  NOR2_X1   g0217(.A1(KEYINPUT5), .A2(G41), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n419), .A2(new_n269), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n256), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G270), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G169), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n291), .B(new_n294), .C1(G1), .C2(new_n254), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(new_n221), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G283), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n216), .C1(G33), .C2(new_n227), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n430), .B(new_n279), .C1(new_n216), .C2(G116), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT20), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n432), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n428), .B1(G116), .B2(new_n294), .C1(new_n433), .C2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT21), .B1(new_n426), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(KEYINPUT21), .A3(G169), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n414), .A2(G179), .A3(new_n420), .A4(new_n422), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT75), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT75), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n442), .A3(new_n435), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n325), .A2(G116), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n216), .A2(G107), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n445), .A2(G20), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n409), .A2(new_n216), .A3(G87), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT76), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n409), .A2(KEYINPUT76), .A3(new_n216), .A4(G87), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(KEYINPUT22), .A3(new_n452), .ZN(new_n453));
  OR4_X1    g0253(.A1(KEYINPUT22), .A2(new_n303), .A3(G20), .A4(new_n250), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT24), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n446), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n456), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n279), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n427), .B(KEYINPUT74), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G107), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n294), .A2(G107), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n464), .B(KEYINPUT25), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n326), .A2(G1698), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n467), .A2(G250), .B1(G294), .B2(new_n325), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n326), .A2(new_n228), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT77), .B1(new_n469), .B2(G1698), .ZN(new_n470));
  AND4_X1   g0270(.A1(KEYINPUT77), .A2(new_n409), .A3(G257), .A4(G1698), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n468), .B(KEYINPUT78), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n257), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n420), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(G264), .B2(new_n421), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n276), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n425), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n466), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n444), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n227), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(new_n205), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(KEYINPUT6), .A3(G97), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n344), .A2(new_n345), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n491), .A2(G20), .B1(new_n492), .B2(G107), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n283), .B2(new_n281), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n279), .B1(G97), .B2(new_n462), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n326), .A2(new_n308), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT4), .B1(new_n496), .B2(new_n262), .ZN(new_n497));
  INV_X1    g0297(.A(G250), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT4), .A2(G244), .ZN(new_n499));
  OAI221_X1 g0299(.A(new_n429), .B1(new_n305), .B2(new_n498), .C1(new_n263), .C2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n257), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n421), .A2(G257), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n420), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n317), .A2(new_n227), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(G190), .A3(new_n420), .A4(new_n502), .ZN(new_n506));
  AND4_X1   g0306(.A1(new_n495), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(G169), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n501), .A2(G179), .A3(new_n420), .A4(new_n502), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n508), .A2(new_n509), .B1(new_n495), .B2(new_n505), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n409), .A2(G244), .A3(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n409), .A2(new_n262), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n445), .C1(new_n513), .C2(new_n226), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n257), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n256), .B(G250), .C1(G1), .C2(new_n415), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n416), .A2(G274), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n276), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n409), .A2(new_n216), .A3(G68), .ZN(new_n520));
  OAI221_X1 g0320(.A(KEYINPUT19), .B1(new_n206), .B2(G87), .C1(new_n266), .C2(G20), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n254), .A2(new_n227), .A3(G20), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n520), .B(new_n521), .C1(KEYINPUT19), .C2(new_n522), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n279), .B1(new_n317), .B2(new_n315), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n315), .B2(new_n461), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n519), .B(new_n525), .C1(G169), .C2(new_n518), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n462), .A2(G87), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n527), .A2(new_n524), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n528), .B(new_n530), .C1(new_n371), .C2(new_n529), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n476), .A2(G190), .A3(new_n478), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n460), .A2(new_n533), .A3(new_n463), .A4(new_n465), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n480), .A2(new_n369), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n511), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n435), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n423), .B2(new_n371), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G200), .B2(new_n423), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n484), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n408), .A2(new_n540), .ZN(G372));
  INV_X1    g0341(.A(new_n526), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n495), .A2(new_n505), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT79), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n508), .A2(new_n544), .A3(new_n509), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n508), .B2(new_n509), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n526), .A2(new_n531), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT26), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n542), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n510), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT26), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n436), .B1(new_n435), .B2(new_n439), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n483), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n551), .B(new_n553), .C1(new_n555), .C2(new_n536), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n408), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n400), .A2(new_n375), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n368), .B1(new_n321), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n405), .B1(new_n559), .B2(new_n397), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n557), .A2(new_n560), .ZN(G369));
  INV_X1    g0361(.A(G13), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n215), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n564), .A2(KEYINPUT27), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(KEYINPUT27), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(G213), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G343), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n483), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n466), .A2(new_n569), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT80), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n534), .A2(new_n535), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n570), .B1(new_n574), .B2(new_n483), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n444), .A2(new_n569), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n570), .ZN(new_n580));
  INV_X1    g0380(.A(new_n444), .ZN(new_n581));
  INV_X1    g0381(.A(new_n569), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n537), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n539), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n583), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n581), .A2(new_n584), .B1(new_n554), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G330), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n576), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n580), .A2(new_n589), .ZN(G399));
  INV_X1    g0390(.A(new_n217), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G41), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(G1), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n212), .B2(new_n593), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n596), .B(KEYINPUT28), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n511), .B(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n573), .A2(new_n548), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(new_n484), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n550), .B1(new_n548), .B2(new_n552), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(KEYINPUT85), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n549), .A2(KEYINPUT26), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(KEYINPUT85), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n601), .B(new_n526), .C1(new_n603), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n582), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT87), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n610), .A3(new_n582), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(KEYINPUT29), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n556), .A2(new_n582), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT29), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n540), .A2(new_n582), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n503), .A2(new_n529), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n424), .A2(G179), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n479), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n438), .A2(new_n529), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n501), .A2(new_n502), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n476), .A2(new_n620), .A3(new_n478), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(KEYINPUT30), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT30), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(KEYINPUT82), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n623), .A2(KEYINPUT30), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n619), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n569), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT83), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n619), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n619), .A2(new_n633), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n635), .B(new_n636), .C1(new_n625), .C2(new_n629), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n569), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT31), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n616), .A2(new_n632), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT84), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n644), .A3(G330), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n615), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n597), .B1(new_n647), .B2(G1), .ZN(G364));
  OR2_X1    g0448(.A1(new_n213), .A2(G45), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n409), .A2(new_n591), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n247), .C2(new_n415), .ZN(new_n651));
  INV_X1    g0451(.A(G355), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n261), .A2(new_n217), .ZN(new_n653));
  XOR2_X1   g0453(.A(new_n653), .B(KEYINPUT89), .Z(new_n654));
  OAI221_X1 g0454(.A(new_n651), .B1(G116), .B2(new_n217), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(G13), .A2(G33), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G20), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n208), .B1(G20), .B2(new_n425), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n563), .A2(G45), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n593), .A2(G1), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT88), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n216), .A2(G190), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n276), .A2(G200), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G311), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n216), .A2(new_n371), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n369), .A2(G179), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n665), .A2(new_n671), .ZN(new_n673));
  INV_X1    g0473(.A(G283), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n672), .A2(new_n412), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(G179), .A2(G200), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n665), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AOI211_X1 g0478(.A(new_n669), .B(new_n675), .C1(G329), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n371), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n261), .B1(new_n681), .B2(G326), .ZN(new_n682));
  INV_X1    g0482(.A(G322), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n670), .A2(new_n666), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(G190), .ZN(new_n686));
  XNOR2_X1  g0486(.A(KEYINPUT33), .B(G317), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(G294), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n216), .B1(new_n676), .B2(G190), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n679), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT90), .ZN(new_n692));
  INV_X1    g0492(.A(new_n672), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G87), .ZN(new_n694));
  INV_X1    g0494(.A(new_n681), .ZN(new_n695));
  OAI221_X1 g0495(.A(new_n694), .B1(new_n227), .B2(new_n690), .C1(new_n695), .C2(new_n202), .ZN(new_n696));
  AOI211_X1 g0496(.A(new_n303), .B(new_n696), .C1(G68), .C2(new_n686), .ZN(new_n697));
  INV_X1    g0497(.A(new_n667), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G77), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n678), .A2(G159), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT32), .Z(new_n701));
  INV_X1    g0501(.A(new_n684), .ZN(new_n702));
  INV_X1    g0502(.A(new_n673), .ZN(new_n703));
  AOI22_X1  g0503(.A1(G58), .A2(new_n702), .B1(new_n703), .B2(G107), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n697), .A2(new_n699), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n692), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n664), .B1(new_n706), .B2(new_n659), .ZN(new_n707));
  INV_X1    g0507(.A(new_n658), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n661), .B(new_n707), .C1(new_n586), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n587), .A2(new_n663), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n586), .A2(G330), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(G396));
  NAND2_X1  g0512(.A1(new_n319), .A2(new_n569), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n379), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n320), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n320), .A2(new_n569), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n646), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(new_n613), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n663), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n303), .B1(new_n672), .B2(new_n486), .ZN(new_n721));
  INV_X1    g0521(.A(new_n686), .ZN(new_n722));
  OAI22_X1  g0522(.A1(new_n722), .A2(new_n674), .B1(new_n695), .B2(new_n412), .ZN(new_n723));
  INV_X1    g0523(.A(new_n690), .ZN(new_n724));
  AOI211_X1 g0524(.A(new_n721), .B(new_n723), .C1(G97), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n678), .A2(G311), .ZN(new_n726));
  AOI22_X1  g0526(.A1(G294), .A2(new_n702), .B1(new_n698), .B2(G116), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n703), .A2(G87), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(new_n726), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n409), .B1(new_n244), .B2(new_n690), .ZN(new_n731));
  INV_X1    g0531(.A(G132), .ZN(new_n732));
  OAI22_X1  g0532(.A1(new_n672), .A2(new_n202), .B1(new_n677), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n698), .A2(G159), .B1(G137), .B2(new_n681), .ZN(new_n734));
  XOR2_X1   g0534(.A(KEYINPUT92), .B(G143), .Z(new_n735));
  OAI221_X1 g0535(.A(new_n734), .B1(new_n387), .B2(new_n722), .C1(new_n684), .C2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT34), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n731), .B(new_n733), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n738), .B1(new_n737), .B2(new_n736), .C1(new_n225), .C2(new_n673), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n664), .B1(new_n740), .B2(new_n659), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n659), .A2(new_n656), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n717), .ZN(new_n744));
  OAI221_X1 g0544(.A(new_n741), .B1(G77), .B2(new_n743), .C1(new_n744), .C2(new_n657), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n720), .A2(new_n745), .ZN(G384));
  INV_X1    g0546(.A(KEYINPUT40), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n349), .A2(new_n353), .ZN(new_n748));
  INV_X1    g0548(.A(new_n567), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n748), .A2(KEYINPUT94), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT94), .B1(new_n748), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n373), .A2(new_n353), .A3(new_n349), .ZN(new_n753));
  NOR4_X1   g0553(.A1(new_n752), .A2(KEYINPUT37), .A3(new_n367), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT37), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n341), .A2(new_n279), .ZN(new_n757));
  AOI21_X1  g0557(.A(KEYINPUT16), .B1(new_n338), .B2(new_n340), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n353), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n363), .A2(new_n366), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n760), .B2(new_n749), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n761), .A2(new_n374), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n755), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n376), .A2(new_n749), .A3(new_n759), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT38), .Z(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n638), .A2(KEYINPUT31), .ZN(new_n768));
  OR3_X1    g0568(.A1(new_n622), .A2(new_n627), .A3(new_n628), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n634), .B1(new_n769), .B2(new_n624), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n582), .B1(new_n770), .B2(new_n636), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n540), .B2(new_n582), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n768), .B1(new_n772), .B2(new_n631), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n301), .A2(new_n569), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n302), .A2(new_n400), .A3(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n301), .B(new_n569), .C1(new_n277), .C2(new_n401), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n773), .A2(new_n744), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n747), .B1(new_n767), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT100), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT96), .B1(new_n753), .B2(new_n367), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n748), .A2(new_n760), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT96), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n784), .A2(new_n785), .A3(new_n374), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(new_n751), .C2(new_n750), .ZN(new_n787));
  AND3_X1   g0587(.A1(new_n787), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n788));
  AOI21_X1  g0588(.A(KEYINPUT97), .B1(new_n787), .B2(KEYINPUT37), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n788), .A2(new_n789), .A3(new_n754), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n376), .A2(new_n752), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n782), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT98), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n763), .A2(KEYINPUT38), .A3(new_n764), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n787), .A2(KEYINPUT37), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT97), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n787), .A2(KEYINPUT97), .A3(KEYINPUT37), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n799), .A2(new_n755), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n791), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(KEYINPUT98), .A3(new_n782), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n795), .A2(new_n796), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT99), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT99), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n795), .A2(new_n803), .A3(new_n806), .A4(new_n796), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n773), .A2(KEYINPUT40), .A3(new_n744), .A4(new_n777), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n780), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AOI211_X1 g0611(.A(KEYINPUT100), .B(new_n809), .C1(new_n805), .C2(new_n807), .ZN(new_n812));
  OAI211_X1 g0612(.A(G330), .B(new_n779), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n408), .A2(new_n773), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT101), .ZN(new_n817));
  INV_X1    g0617(.A(new_n779), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT98), .B1(new_n802), .B2(new_n782), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n794), .B(new_n781), .C1(new_n801), .C2(new_n791), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n806), .B1(new_n821), .B2(new_n796), .ZN(new_n822));
  INV_X1    g0622(.A(new_n807), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n810), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n808), .A2(new_n780), .A3(new_n810), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n814), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n804), .A2(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n766), .A2(KEYINPUT39), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n302), .A2(new_n569), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n716), .A2(KEYINPUT93), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n613), .C2(new_n717), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n766), .A2(new_n777), .A3(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n368), .A2(new_n749), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n615), .A2(new_n408), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n841), .A2(new_n560), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n840), .B(new_n842), .Z(new_n843));
  OR2_X1    g0643(.A1(new_n829), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(G1), .B1(new_n562), .B2(G20), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n829), .A2(new_n843), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT103), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n844), .A2(KEYINPUT102), .A3(new_n845), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n849), .A2(KEYINPUT103), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n848), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n221), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n854));
  INV_X1    g0654(.A(new_n211), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(KEYINPUT35), .C2(new_n491), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT36), .ZN(new_n857));
  OAI21_X1  g0657(.A(G77), .B1(new_n244), .B2(new_n225), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n858), .A2(new_n212), .B1(G50), .B2(new_n225), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(G1), .A3(new_n562), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n853), .A2(new_n857), .A3(new_n860), .ZN(G367));
  INV_X1    g0661(.A(new_n580), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n543), .A2(new_n569), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n599), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n547), .A2(new_n582), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT42), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n862), .B(new_n866), .C1(new_n867), .C2(new_n570), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n579), .A2(new_n866), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n869), .A2(KEYINPUT42), .B1(new_n510), .B2(new_n582), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n588), .A2(new_n866), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n528), .A2(new_n582), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n542), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n548), .B2(new_n873), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT43), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n871), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n872), .B1(new_n871), .B2(new_n876), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n875), .A2(KEYINPUT43), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OR3_X1    g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n877), .B2(new_n878), .ZN(new_n882));
  XOR2_X1   g0682(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n883));
  XOR2_X1   g0683(.A(new_n592), .B(new_n883), .Z(new_n884));
  INV_X1    g0684(.A(KEYINPUT45), .ZN(new_n885));
  INV_X1    g0685(.A(new_n866), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n862), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT45), .B1(new_n580), .B2(new_n866), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(KEYINPUT44), .C1(new_n580), .C2(new_n866), .ZN(new_n891));
  XNOR2_X1  g0691(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n862), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n889), .A2(new_n589), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n579), .A2(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n576), .A2(new_n578), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n579), .A2(KEYINPUT106), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(new_n587), .ZN(new_n899));
  INV_X1    g0699(.A(new_n647), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n891), .B(new_n893), .C1(new_n887), .C2(new_n888), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n588), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n894), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n884), .B1(new_n904), .B2(new_n647), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n662), .A2(G1), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n881), .B(new_n882), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n650), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n660), .B1(new_n217), .B2(new_n315), .C1(new_n241), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n673), .A2(new_n283), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n672), .A2(new_n244), .B1(new_n667), .B2(new_n202), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n910), .B(new_n911), .C1(G137), .C2(new_n678), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n724), .A2(G68), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n686), .A2(G159), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n695), .B2(new_n735), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(G150), .B2(new_n702), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n912), .A2(new_n261), .A3(new_n913), .A4(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n684), .A2(new_n412), .B1(new_n673), .B2(new_n227), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n326), .B1(new_n695), .B2(new_n668), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n918), .B(new_n919), .C1(G283), .C2(new_n698), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT46), .B1(new_n693), .B2(G116), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n722), .A2(new_n689), .B1(new_n690), .B2(new_n486), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n693), .A2(KEYINPUT46), .A3(G116), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT107), .Z(new_n925));
  NAND3_X1  g0725(.A1(new_n920), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(G317), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n677), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n917), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT47), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n664), .B1(new_n930), .B2(new_n659), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n909), .B(new_n931), .C1(new_n875), .C2(new_n708), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n907), .A2(new_n932), .ZN(G387));
  INV_X1    g0733(.A(new_n594), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n313), .A2(G50), .ZN(new_n935));
  XOR2_X1   g0735(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g0738(.A1(G68), .A2(G77), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n937), .A2(new_n415), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n650), .B(new_n940), .C1(new_n238), .C2(new_n415), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n941), .B1(G107), .B2(new_n217), .C1(new_n594), .C2(new_n654), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n660), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n698), .A2(G303), .B1(G322), .B2(new_n681), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n668), .B2(new_n722), .C1(new_n927), .C2(new_n684), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT48), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n674), .B2(new_n690), .C1(new_n689), .C2(new_n672), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT49), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n678), .A2(G326), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n409), .B1(G116), .B2(new_n703), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G97), .A2(new_n703), .B1(new_n678), .B2(G150), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n202), .B2(new_n684), .C1(new_n283), .C2(new_n672), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G159), .B2(new_n681), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n315), .A2(new_n690), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n722), .A2(new_n313), .B1(new_n667), .B2(new_n225), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT109), .Z(new_n960));
  NAND4_X1  g0760(.A1(new_n956), .A2(new_n409), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT110), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n953), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n664), .B1(new_n963), .B2(new_n659), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n943), .B(new_n964), .C1(new_n575), .C2(new_n708), .ZN(new_n965));
  INV_X1    g0765(.A(new_n906), .ZN(new_n966));
  INV_X1    g0766(.A(new_n899), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n592), .B1(new_n967), .B2(new_n647), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n965), .B1(new_n966), .B2(new_n899), .C1(new_n968), .C2(new_n901), .ZN(G393));
  NAND3_X1  g0769(.A1(new_n894), .A2(new_n906), .A3(new_n903), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n660), .B1(new_n227), .B2(new_n217), .C1(new_n252), .C2(new_n908), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n690), .A2(new_n283), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n728), .B1(new_n313), .B2(new_n667), .C1(new_n677), .C2(new_n735), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n972), .B(new_n973), .C1(G68), .C2(new_n693), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n326), .B1(G50), .B2(new_n686), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n702), .A2(G159), .B1(G150), .B2(new_n681), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT51), .Z(new_n977));
  NAND3_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n672), .A2(new_n674), .B1(new_n677), .B2(new_n683), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT111), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n695), .A2(new_n927), .B1(new_n684), .B2(new_n668), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT52), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n261), .B1(new_n698), .B2(G294), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n722), .A2(new_n412), .B1(new_n690), .B2(new_n221), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G107), .B2(new_n703), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n978), .B1(new_n980), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n664), .B1(new_n987), .B2(new_n659), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n971), .B(new_n988), .C1(new_n866), .C2(new_n708), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n970), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n901), .B1(new_n903), .B2(new_n894), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n991), .A2(new_n593), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n990), .B1(new_n992), .B2(new_n904), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(G390));
  AND3_X1   g0794(.A1(new_n841), .A2(new_n560), .A3(new_n815), .ZN(new_n995));
  INV_X1    g0795(.A(new_n837), .ZN(new_n996));
  INV_X1    g0796(.A(new_n645), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n644), .B1(new_n641), .B2(G330), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n744), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n777), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G330), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n778), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n996), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n646), .A2(new_n744), .A3(new_n777), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n609), .A2(new_n611), .A3(new_n716), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n715), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n773), .A2(G330), .A3(new_n744), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n1000), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n995), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n833), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n808), .B(new_n1013), .C1(new_n1008), .C2(new_n1000), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n999), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n996), .B2(new_n1000), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n830), .A2(new_n831), .A3(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n777), .A4(new_n1017), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1012), .B(new_n1018), .C1(new_n1019), .C2(new_n1003), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n841), .A2(new_n560), .A3(new_n815), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n777), .B1(new_n646), .B2(new_n744), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n837), .B1(new_n1022), .B2(new_n1003), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1006), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND4_X1   g0825(.A1(new_n1015), .A2(new_n1014), .A3(new_n777), .A4(new_n1017), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1003), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1020), .A2(new_n1028), .A3(new_n592), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G68), .A2(new_n703), .B1(new_n678), .B2(G294), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n227), .B2(new_n667), .C1(new_n221), .C2(new_n684), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n694), .B1(new_n722), .B2(new_n486), .C1(new_n674), .C2(new_n695), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1031), .A2(new_n972), .A3(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(KEYINPUT54), .B(G143), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n698), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G50), .A2(new_n703), .B1(new_n678), .B2(G125), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n732), .B2(new_n684), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n672), .A2(KEYINPUT53), .A3(new_n387), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n681), .A2(G128), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n724), .A2(G159), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT53), .B1(new_n672), .B2(new_n387), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(G137), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n261), .B1(new_n722), .B2(new_n1043), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1037), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1033), .A2(new_n303), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n664), .B1(new_n1047), .B2(new_n659), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n832), .B2(new_n657), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n313), .B2(new_n742), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1018), .B1(new_n1019), .B2(new_n1003), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n906), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1029), .A2(new_n1052), .ZN(G378));
  INV_X1    g0853(.A(KEYINPUT116), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n397), .A2(new_n404), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT114), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n390), .A2(new_n749), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1058));
  XOR2_X1   g0858(.A(new_n1057), .B(new_n1058), .Z(new_n1059));
  XNOR2_X1  g0859(.A(new_n1056), .B(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT115), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n827), .B2(G330), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n813), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n840), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n813), .A2(new_n1063), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n825), .A2(new_n826), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(G330), .A3(new_n779), .A4(new_n1061), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n840), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n966), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1060), .A2(new_n656), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n742), .A2(new_n202), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n315), .A2(new_n667), .B1(new_n674), .B2(new_n677), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G58), .B2(new_n703), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n283), .B2(new_n672), .C1(new_n486), .C2(new_n684), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n913), .B1(new_n722), .B2(new_n227), .C1(new_n221), .C2(new_n695), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1076), .A2(G41), .A3(new_n409), .A4(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT58), .Z(new_n1079));
  AOI22_X1  g0879(.A1(new_n724), .A2(G150), .B1(G125), .B2(new_n681), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT113), .Z(new_n1081));
  NAND2_X1  g0881(.A1(new_n702), .A2(G128), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n686), .A2(G132), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n693), .A2(new_n1034), .B1(new_n698), .B2(G137), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1081), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT59), .Z(new_n1086));
  AOI21_X1  g0886(.A(G41), .B1(new_n703), .B2(G159), .ZN(new_n1087));
  AOI21_X1  g0887(.A(G33), .B1(new_n678), .B2(G124), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n333), .ZN(new_n1090));
  AOI21_X1  g0890(.A(G41), .B1(new_n1090), .B2(G33), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1079), .B(new_n1089), .C1(G50), .C2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n663), .B1(new_n1092), .B2(new_n659), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1072), .A2(new_n1073), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1054), .B1(new_n1071), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1069), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n906), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n1094), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1065), .A2(KEYINPUT117), .A3(new_n1070), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT57), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n1028), .B2(new_n995), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1066), .A2(new_n1068), .A3(new_n1105), .A4(new_n1069), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1028), .A2(new_n995), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1103), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1110), .A3(new_n592), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1101), .A2(new_n1111), .ZN(G375));
  OAI21_X1  g0912(.A(new_n906), .B1(new_n1011), .B2(new_n1005), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n672), .A2(new_n227), .B1(new_n677), .B2(new_n412), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT119), .Z(new_n1115));
  AOI22_X1  g0915(.A1(new_n686), .A2(G116), .B1(new_n681), .B2(G294), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n486), .B2(new_n667), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n958), .A3(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n261), .B(new_n910), .C1(G283), .C2(new_n702), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n1117), .B2(KEYINPUT118), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n724), .A2(G50), .B1(new_n1034), .B2(new_n686), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n244), .B2(new_n673), .C1(new_n732), .C2(new_n695), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G150), .A2(new_n698), .B1(new_n678), .B2(G128), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n693), .A2(G159), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n702), .A2(G137), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1124), .A2(new_n409), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1119), .A2(new_n1121), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n664), .B1(new_n1128), .B2(new_n659), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(G68), .B2(new_n743), .C1(new_n777), .C2(new_n657), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1113), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n884), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1012), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT121), .ZN(G381));
  NOR4_X1   g0938(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1139));
  INV_X1    g0939(.A(G378), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n593), .B1(new_n1109), .B2(new_n1103), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1096), .A2(new_n1100), .B1(new_n1141), .B2(new_n1107), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n907), .A2(new_n993), .A3(new_n932), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .A4(new_n1144), .ZN(G407));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1140), .ZN(new_n1146));
  OAI211_X1 g0946(.A(G407), .B(G213), .C1(G343), .C2(new_n1146), .ZN(G409));
  INV_X1    g0947(.A(KEYINPUT125), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT61), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1102), .A2(new_n906), .A3(new_n1106), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1029), .A2(new_n1052), .A3(new_n1094), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1108), .B(new_n1134), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n568), .A2(G213), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(KEYINPUT124), .C1(new_n1140), .C2(new_n1142), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT124), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1140), .B1(new_n1101), .B2(new_n1111), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT60), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n593), .B1(new_n1135), .B2(new_n1161), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1162), .B(new_n1012), .C1(new_n1161), .C2(new_n1135), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1133), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(G384), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1133), .A2(new_n1163), .A3(G384), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n568), .A2(G213), .A3(G2897), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1156), .A2(new_n1160), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1168), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT62), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1149), .B(new_n1171), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1168), .ZN(new_n1176));
  AOI21_X1  g0976(.A(KEYINPUT122), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n1158), .A2(new_n1159), .A3(new_n1168), .A4(new_n1178), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1179), .A3(KEYINPUT62), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1148), .B1(new_n1174), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n993), .B1(new_n907), .B2(new_n932), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(G393), .B(G396), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1183), .A2(new_n1143), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1144), .B2(new_n1182), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1187), .A3(KEYINPUT126), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT126), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(G375), .A2(G378), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT124), .B1(new_n1192), .B2(new_n1155), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1158), .A2(new_n1159), .A3(new_n1157), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1176), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT62), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1171), .A2(new_n1149), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1192), .A2(new_n1155), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1178), .B1(new_n1198), .B2(new_n1168), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1175), .A2(KEYINPUT122), .A3(new_n1176), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1173), .A3(new_n1200), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1196), .A2(new_n1197), .A3(KEYINPUT125), .A4(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1181), .A2(new_n1191), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT123), .B(KEYINPUT63), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1185), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1187), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT63), .B(new_n1176), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT61), .B1(new_n1198), .B2(new_n1170), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1203), .A2(new_n1211), .ZN(G405));
  NAND2_X1  g1012(.A1(new_n1192), .A2(new_n1146), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(new_n1176), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1190), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT127), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1215), .A2(new_n1216), .A3(new_n1188), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT127), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1214), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1214), .B2(new_n1218), .ZN(G402));
endmodule


