

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U548 ( .A(n710), .ZN(n748) );
  BUF_X1 U549 ( .A(n674), .Z(n598) );
  NOR2_X1 U550 ( .A1(n623), .A2(G651), .ZN(n644) );
  NOR2_X2 U551 ( .A1(n537), .A2(n536), .ZN(G160) );
  XNOR2_X1 U552 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n526) );
  NOR2_X1 U553 ( .A1(G543), .A2(G651), .ZN(n640) );
  NAND2_X1 U554 ( .A1(n640), .A2(G89), .ZN(n513) );
  XNOR2_X1 U555 ( .A(n513), .B(KEYINPUT4), .ZN(n515) );
  XOR2_X1 U556 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  INV_X1 U557 ( .A(G651), .ZN(n517) );
  NOR2_X1 U558 ( .A1(n623), .A2(n517), .ZN(n634) );
  NAND2_X1 U559 ( .A1(G76), .A2(n634), .ZN(n514) );
  NAND2_X1 U560 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U561 ( .A(n516), .B(KEYINPUT5), .ZN(n524) );
  XNOR2_X1 U562 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n522) );
  NOR2_X1 U563 ( .A1(G543), .A2(n517), .ZN(n518) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n518), .Z(n636) );
  NAND2_X1 U565 ( .A1(G63), .A2(n636), .ZN(n520) );
  NAND2_X1 U566 ( .A1(G51), .A2(n644), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n522), .B(n521), .ZN(n523) );
  NAND2_X1 U569 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U570 ( .A(n526), .B(n525), .ZN(G168) );
  XOR2_X1 U571 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U572 ( .A(G2105), .ZN(n533) );
  AND2_X4 U573 ( .A1(n533), .A2(G2104), .ZN(n884) );
  NAND2_X1 U574 ( .A1(G101), .A2(n884), .ZN(n527) );
  XNOR2_X1 U575 ( .A(n527), .B(KEYINPUT65), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT23), .ZN(n532) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT17), .B(n529), .Z(n530) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(n530), .ZN(n674) );
  NAND2_X1 U580 ( .A1(G137), .A2(n674), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n537) );
  NOR2_X1 U582 ( .A1(G2104), .A2(n533), .ZN(n879) );
  NAND2_X1 U583 ( .A1(G125), .A2(n879), .ZN(n535) );
  AND2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NAND2_X1 U585 ( .A1(G113), .A2(n880), .ZN(n534) );
  NAND2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT103), .B(G2435), .Z(n539) );
  XNOR2_X1 U588 ( .A(G2430), .B(G2438), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n539), .B(n538), .ZN(n546) );
  XOR2_X1 U590 ( .A(G2446), .B(G2454), .Z(n541) );
  XNOR2_X1 U591 ( .A(G2451), .B(G2443), .ZN(n540) );
  XNOR2_X1 U592 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U593 ( .A(n542), .B(G2427), .Z(n544) );
  XNOR2_X1 U594 ( .A(G1341), .B(G1348), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n546), .B(n545), .ZN(n547) );
  AND2_X1 U597 ( .A1(n547), .A2(G14), .ZN(G401) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G120), .ZN(G236) );
  INV_X1 U602 ( .A(G69), .ZN(G235) );
  INV_X1 U603 ( .A(G108), .ZN(G238) );
  NAND2_X1 U604 ( .A1(G52), .A2(n644), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(n548), .Z(n555) );
  NAND2_X1 U606 ( .A1(G90), .A2(n640), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G77), .A2(n634), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n551), .B(KEYINPUT9), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G64), .A2(n636), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U612 ( .A1(n555), .A2(n554), .ZN(G171) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n560) );
  XOR2_X1 U614 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n557) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT70), .B(n558), .Z(n829) );
  NAND2_X1 U618 ( .A1(n829), .A2(G567), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n560), .B(n559), .ZN(G234) );
  NAND2_X1 U620 ( .A1(G56), .A2(n636), .ZN(n561) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n561), .Z(n567) );
  NAND2_X1 U622 ( .A1(n640), .A2(G81), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G68), .A2(n634), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  NOR2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U628 ( .A1(n644), .A2(G43), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n937) );
  INV_X1 U630 ( .A(G860), .ZN(n605) );
  OR2_X1 U631 ( .A1(n937), .A2(n605), .ZN(G153) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G79), .A2(n634), .ZN(n576) );
  NAND2_X1 U634 ( .A1(G92), .A2(n640), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G66), .A2(n636), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G54), .A2(n644), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT73), .B(n572), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT15), .ZN(n936) );
  OR2_X1 U642 ( .A1(n936), .A2(G868), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT74), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G868), .A2(G286), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G78), .A2(n634), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G53), .A2(n644), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G91), .A2(n640), .ZN(n584) );
  NAND2_X1 U651 ( .A1(G65), .A2(n636), .ZN(n583) );
  NAND2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(n587), .B(KEYINPUT69), .Z(n946) );
  OR2_X1 U655 ( .A1(n946), .A2(G868), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G297) );
  INV_X1 U657 ( .A(n946), .ZN(G299) );
  NAND2_X1 U658 ( .A1(n605), .A2(G559), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n590), .A2(n936), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U661 ( .A1(G868), .A2(n937), .ZN(n594) );
  NAND2_X1 U662 ( .A1(G868), .A2(n936), .ZN(n592) );
  NOR2_X1 U663 ( .A1(G559), .A2(n592), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G282) );
  NAND2_X1 U665 ( .A1(n879), .A2(G123), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT18), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G111), .A2(n880), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n884), .A2(G99), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G135), .A2(n598), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n922) );
  XNOR2_X1 U673 ( .A(n922), .B(G2096), .ZN(n603) );
  INV_X1 U674 ( .A(G2100), .ZN(n835) );
  NAND2_X1 U675 ( .A1(n603), .A2(n835), .ZN(G156) );
  NAND2_X1 U676 ( .A1(G559), .A2(n936), .ZN(n604) );
  XOR2_X1 U677 ( .A(n937), .B(n604), .Z(n652) );
  NAND2_X1 U678 ( .A1(n605), .A2(n652), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G67), .A2(n636), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G55), .A2(n644), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G93), .A2(n640), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G80), .A2(n634), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n655) );
  XOR2_X1 U686 ( .A(n612), .B(n655), .Z(G145) );
  NAND2_X1 U687 ( .A1(G60), .A2(n636), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G47), .A2(n644), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G85), .A2(n640), .ZN(n615) );
  XNOR2_X1 U691 ( .A(KEYINPUT67), .B(n615), .ZN(n616) );
  NOR2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n634), .A2(G72), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G290) );
  NAND2_X1 U695 ( .A1(G49), .A2(n644), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U698 ( .A1(n636), .A2(n622), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G87), .A2(n623), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT77), .B(n624), .Z(n625) );
  NAND2_X1 U701 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U702 ( .A1(G88), .A2(n640), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G75), .A2(n634), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U705 ( .A(KEYINPUT80), .B(n629), .ZN(n633) );
  NAND2_X1 U706 ( .A1(G62), .A2(n636), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G50), .A2(n644), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(G166) );
  NAND2_X1 U710 ( .A1(G73), .A2(n634), .ZN(n635) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n635), .Z(n639) );
  NAND2_X1 U712 ( .A1(n636), .A2(G61), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT78), .B(n637), .Z(n638) );
  NOR2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U715 ( .A1(n640), .A2(G86), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT79), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G48), .A2(n644), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(G305) );
  XNOR2_X1 U720 ( .A(G288), .B(KEYINPUT19), .ZN(n648) );
  XOR2_X1 U721 ( .A(G299), .B(G166), .Z(n647) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U723 ( .A(n655), .B(n649), .Z(n650) );
  XNOR2_X1 U724 ( .A(G290), .B(n650), .ZN(n651) );
  XNOR2_X1 U725 ( .A(n651), .B(G305), .ZN(n895) );
  XNOR2_X1 U726 ( .A(n895), .B(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n653), .A2(G868), .ZN(n654) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n654), .Z(n657) );
  OR2_X1 U729 ( .A1(n655), .A2(G868), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n659) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U738 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U739 ( .A1(G235), .A2(G236), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n663), .B(KEYINPUT83), .ZN(n664) );
  NOR2_X1 U741 ( .A1(G238), .A2(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G57), .A2(n665), .ZN(n907) );
  NAND2_X1 U743 ( .A1(n907), .A2(G567), .ZN(n670) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U746 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G96), .A2(n668), .ZN(n908) );
  NAND2_X1 U748 ( .A1(n908), .A2(G2106), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n909) );
  NOR2_X1 U750 ( .A1(n671), .A2(n909), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n672), .B(KEYINPUT84), .ZN(n832) );
  NAND2_X1 U752 ( .A1(n832), .A2(G36), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT85), .B(n673), .Z(G176) );
  NAND2_X1 U754 ( .A1(n884), .A2(G102), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G138), .A2(n674), .ZN(n675) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U757 ( .A1(G126), .A2(n879), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G114), .A2(n880), .ZN(n677) );
  NAND2_X1 U759 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U760 ( .A1(n680), .A2(n679), .ZN(G164) );
  XOR2_X1 U761 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  XNOR2_X1 U762 ( .A(G1986), .B(G290), .ZN(n956) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n683) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n683), .A2(n681), .ZN(n824) );
  NAND2_X1 U766 ( .A1(n956), .A2(n824), .ZN(n814) );
  INV_X1 U767 ( .A(KEYINPUT90), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n682), .B(n681), .ZN(n684) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n686) );
  INV_X1 U770 ( .A(KEYINPUT64), .ZN(n685) );
  XNOR2_X2 U771 ( .A(n686), .B(n685), .ZN(n710) );
  NAND2_X1 U772 ( .A1(n748), .A2(G8), .ZN(n775) );
  NOR2_X1 U773 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U774 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NOR2_X1 U775 ( .A1(n775), .A2(n688), .ZN(n764) );
  NOR2_X1 U776 ( .A1(n748), .A2(G2084), .ZN(n690) );
  INV_X1 U777 ( .A(KEYINPUT91), .ZN(n689) );
  XNOR2_X1 U778 ( .A(n690), .B(n689), .ZN(n730) );
  NAND2_X1 U779 ( .A1(G8), .A2(n730), .ZN(n746) );
  XNOR2_X1 U780 ( .A(G2078), .B(KEYINPUT93), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n691), .B(KEYINPUT25), .ZN(n996) );
  NAND2_X1 U782 ( .A1(n996), .A2(n710), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n748), .A2(G1961), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U785 ( .A(n694), .B(KEYINPUT94), .Z(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(G171), .ZN(n726) );
  INV_X1 U787 ( .A(n748), .ZN(n695) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n695), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n748), .A2(G1348), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U791 ( .A(n698), .B(KEYINPUT96), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n748), .A2(G1341), .ZN(n700) );
  INV_X1 U793 ( .A(n937), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n704) );
  XNOR2_X1 U795 ( .A(G1996), .B(KEYINPUT95), .ZN(n997) );
  INV_X1 U796 ( .A(n997), .ZN(n701) );
  AND2_X1 U797 ( .A1(n710), .A2(n701), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n702), .B(KEYINPUT26), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n708), .A2(n936), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U802 ( .A(KEYINPUT97), .B(n707), .ZN(n717) );
  OR2_X1 U803 ( .A1(n708), .A2(n936), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G2072), .A2(n710), .ZN(n709) );
  XNOR2_X1 U805 ( .A(n709), .B(KEYINPUT27), .ZN(n712) );
  INV_X1 U806 ( .A(G1956), .ZN(n844) );
  NOR2_X1 U807 ( .A1(n710), .A2(n844), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n719) );
  NOR2_X1 U809 ( .A1(n946), .A2(n719), .ZN(n714) );
  INV_X1 U810 ( .A(KEYINPUT28), .ZN(n713) );
  XNOR2_X1 U811 ( .A(n714), .B(n713), .ZN(n718) );
  NAND2_X1 U812 ( .A1(n715), .A2(n718), .ZN(n716) );
  NOR2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n723) );
  INV_X1 U814 ( .A(n718), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n946), .A2(n719), .ZN(n720) );
  NOR2_X1 U816 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U817 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U818 ( .A(n724), .B(KEYINPUT29), .Z(n725) );
  NAND2_X1 U819 ( .A1(n726), .A2(n725), .ZN(n742) );
  INV_X1 U820 ( .A(G1966), .ZN(n727) );
  AND2_X1 U821 ( .A1(G8), .A2(n727), .ZN(n728) );
  AND2_X1 U822 ( .A1(n748), .A2(n728), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT92), .ZN(n743) );
  INV_X1 U824 ( .A(n730), .ZN(n731) );
  NAND2_X1 U825 ( .A1(G8), .A2(n731), .ZN(n732) );
  NOR2_X1 U826 ( .A1(n743), .A2(n732), .ZN(n733) );
  XOR2_X1 U827 ( .A(KEYINPUT30), .B(n733), .Z(n734) );
  NOR2_X1 U828 ( .A1(G168), .A2(n734), .ZN(n738) );
  OR2_X1 U829 ( .A1(n735), .A2(G171), .ZN(n736) );
  XOR2_X1 U830 ( .A(KEYINPUT98), .B(n736), .Z(n737) );
  NOR2_X1 U831 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U832 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n740), .B(n739), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n747) );
  INV_X1 U835 ( .A(n747), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n746), .A2(n745), .ZN(n765) );
  XOR2_X1 U838 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n757) );
  NAND2_X1 U839 ( .A1(n747), .A2(G286), .ZN(n754) );
  NOR2_X1 U840 ( .A1(n748), .A2(G2090), .ZN(n749) );
  XNOR2_X1 U841 ( .A(n749), .B(KEYINPUT100), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n775), .A2(G1971), .ZN(n750) );
  NOR2_X1 U843 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U844 ( .A1(n752), .A2(G303), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U846 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U847 ( .A(n757), .B(n756), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n765), .A2(n767), .ZN(n760) );
  NOR2_X1 U849 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U850 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U852 ( .A(n761), .B(KEYINPUT102), .ZN(n762) );
  AND2_X1 U853 ( .A1(n762), .A2(n775), .ZN(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n782) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n950) );
  AND2_X1 U856 ( .A1(n765), .A2(n950), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n771) );
  INV_X1 U858 ( .A(n950), .ZN(n769) );
  NOR2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G303), .A2(G1971), .ZN(n768) );
  NOR2_X1 U861 ( .A1(n774), .A2(n768), .ZN(n951) );
  OR2_X1 U862 ( .A1(n769), .A2(n951), .ZN(n770) );
  AND2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n775), .A2(n772), .ZN(n773) );
  OR2_X1 U865 ( .A1(KEYINPUT33), .A2(n773), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n774), .A2(KEYINPUT33), .ZN(n776) );
  NOR2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n778) );
  XOR2_X1 U868 ( .A(G1981), .B(G305), .Z(n943) );
  INV_X1 U869 ( .A(n943), .ZN(n777) );
  NOR2_X1 U870 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U872 ( .A1(n782), .A2(n781), .ZN(n812) );
  NAND2_X1 U873 ( .A1(n884), .A2(G104), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G140), .A2(n598), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n785), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G128), .A2(n879), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G116), .A2(n880), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n788), .Z(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n791), .ZN(n892) );
  XNOR2_X1 U883 ( .A(KEYINPUT37), .B(G2067), .ZN(n822) );
  NOR2_X1 U884 ( .A1(n892), .A2(n822), .ZN(n918) );
  NAND2_X1 U885 ( .A1(n824), .A2(n918), .ZN(n820) );
  NAND2_X1 U886 ( .A1(n879), .A2(G119), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G131), .A2(n598), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U889 ( .A1(G107), .A2(n880), .ZN(n794) );
  XNOR2_X1 U890 ( .A(KEYINPUT87), .B(n794), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n884), .A2(G95), .ZN(n797) );
  NAND2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n876) );
  AND2_X1 U894 ( .A1(n876), .A2(G1991), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n879), .A2(G129), .ZN(n800) );
  NAND2_X1 U896 ( .A1(G141), .A2(n598), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n884), .A2(G105), .ZN(n801) );
  XOR2_X1 U899 ( .A(KEYINPUT38), .B(n801), .Z(n802) );
  NOR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n880), .A2(G117), .ZN(n804) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n871) );
  NAND2_X1 U903 ( .A1(G1996), .A2(n871), .ZN(n806) );
  XOR2_X1 U904 ( .A(KEYINPUT88), .B(n806), .Z(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n926) );
  XNOR2_X1 U906 ( .A(KEYINPUT89), .B(n824), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n926), .A2(n809), .ZN(n817) );
  INV_X1 U908 ( .A(n817), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n820), .A2(n810), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n827) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n871), .ZN(n920) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n876), .ZN(n923) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n815) );
  NOR2_X1 U915 ( .A1(n923), .A2(n815), .ZN(n816) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U917 ( .A1(n920), .A2(n818), .ZN(n819) );
  XNOR2_X1 U918 ( .A(n819), .B(KEYINPUT39), .ZN(n821) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n892), .A2(n822), .ZN(n915) );
  NAND2_X1 U921 ( .A1(n823), .A2(n915), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n828), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U926 ( .A(n829), .ZN(G223) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT104), .B(n830), .Z(n831) );
  NAND2_X1 U929 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U932 ( .A(KEYINPUT105), .B(n834), .Z(G188) );
  XOR2_X1 U933 ( .A(G96), .B(KEYINPUT106), .Z(G221) );
  XNOR2_X1 U934 ( .A(n835), .B(G2096), .ZN(n837) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U940 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1976), .B(G1971), .Z(n846) );
  XOR2_X1 U944 ( .A(G1986), .B(n844), .Z(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT41), .B(G1981), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U953 ( .A1(n879), .A2(G124), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G112), .A2(n880), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U957 ( .A1(n884), .A2(G100), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G136), .A2(n598), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U961 ( .A(n922), .B(G162), .Z(n870) );
  NAND2_X1 U962 ( .A1(G127), .A2(n879), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G115), .A2(n880), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT47), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G139), .A2(n598), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n884), .A2(G103), .ZN(n866) );
  XOR2_X1 U969 ( .A(KEYINPUT108), .B(n866), .Z(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(n911) );
  XNOR2_X1 U971 ( .A(G160), .B(n911), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n870), .B(n869), .ZN(n875) );
  XNOR2_X1 U973 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n871), .B(KEYINPUT46), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U976 ( .A(n875), .B(n874), .Z(n878) );
  XOR2_X1 U977 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n891) );
  NAND2_X1 U979 ( .A1(G130), .A2(n879), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G118), .A2(n880), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(KEYINPUT107), .B(n883), .Z(n889) );
  NAND2_X1 U983 ( .A1(n884), .A2(G106), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G142), .A2(n598), .ZN(n885) );
  NAND2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U986 ( .A(n887), .B(KEYINPUT45), .Z(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U988 ( .A(n891), .B(n890), .Z(n893) );
  XOR2_X1 U989 ( .A(n893), .B(n892), .Z(n894) );
  NOR2_X1 U990 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n937), .B(n895), .ZN(n897) );
  XOR2_X1 U992 ( .A(G301), .B(n936), .Z(n896) );
  XNOR2_X1 U993 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n898), .B(G286), .ZN(n899) );
  NOR2_X1 U995 ( .A1(G37), .A2(n899), .ZN(G397) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT49), .B(n900), .Z(n903) );
  NOR2_X1 U998 ( .A1(G401), .A2(n909), .ZN(n901) );
  XNOR2_X1 U999 ( .A(KEYINPUT110), .B(n901), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(KEYINPUT111), .B(n904), .ZN(n906) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(G225) );
  XOR2_X1 U1004 ( .A(KEYINPUT112), .B(G225), .Z(G308) );
  NOR2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(G325) );
  INV_X1 U1007 ( .A(G325), .ZN(G261) );
  INV_X1 U1008 ( .A(n909), .ZN(G319) );
  INV_X1 U1009 ( .A(G57), .ZN(G237) );
  INV_X1 U1010 ( .A(KEYINPUT55), .ZN(n1009) );
  XNOR2_X1 U1011 ( .A(G164), .B(G2078), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n910), .B(KEYINPUT113), .ZN(n913) );
  XOR2_X1 U1013 ( .A(G2072), .B(n911), .Z(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(n914), .B(KEYINPUT50), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n931) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n921), .Z(n925) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n929) );
  XNOR2_X1 U1023 ( .A(G160), .B(G2084), .ZN(n927) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(KEYINPUT52), .B(n932), .ZN(n933) );
  XOR2_X1 U1028 ( .A(KEYINPUT114), .B(n933), .Z(n934) );
  NAND2_X1 U1029 ( .A1(n1009), .A2(n934), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(G29), .ZN(n1018) );
  XOR2_X1 U1031 ( .A(KEYINPUT56), .B(G16), .Z(n964) );
  XNOR2_X1 U1032 ( .A(n936), .B(G1348), .ZN(n941) );
  XOR2_X1 U1033 ( .A(G171), .B(G1961), .Z(n939) );
  XNOR2_X1 U1034 ( .A(n937), .B(G1341), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n961) );
  XNOR2_X1 U1037 ( .A(G1966), .B(KEYINPUT118), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n942), .B(G168), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT57), .ZN(n959) );
  XOR2_X1 U1041 ( .A(n946), .B(G1956), .Z(n947) );
  XNOR2_X1 U1042 ( .A(n947), .B(KEYINPUT119), .ZN(n949) );
  NAND2_X1 U1043 ( .A1(G303), .A2(G1971), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1047 ( .A(KEYINPUT120), .B(n954), .Z(n955) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1049 ( .A(KEYINPUT121), .B(n957), .Z(n958) );
  NAND2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n962), .ZN(n963) );
  NOR2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n1015) );
  XOR2_X1 U1054 ( .A(G20), .B(G1956), .Z(n968) );
  XNOR2_X1 U1055 ( .A(G1341), .B(G19), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1981), .B(G6), .ZN(n965) );
  NOR2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1059 ( .A(KEYINPUT59), .B(G1348), .Z(n969) );
  XNOR2_X1 U1060 ( .A(G4), .B(n969), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(KEYINPUT60), .B(n972), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G21), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1961), .B(G5), .ZN(n973) );
  NOR2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n984) );
  XNOR2_X1 U1067 ( .A(G1986), .B(G24), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(G22), .B(G1971), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1976), .B(KEYINPUT123), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(G23), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT58), .B(n982), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1075 ( .A(n985), .B(KEYINPUT124), .Z(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(G16), .A2(n987), .ZN(n1012) );
  XNOR2_X1 U1078 ( .A(G2084), .B(G34), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n988), .B(KEYINPUT54), .ZN(n1007) );
  XNOR2_X1 U1080 ( .A(G2090), .B(G35), .ZN(n1004) );
  XNOR2_X1 U1081 ( .A(KEYINPUT115), .B(G2067), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(G26), .ZN(n995) );
  XOR2_X1 U1083 ( .A(G25), .B(G1991), .Z(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(G28), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(KEYINPUT116), .B(G2072), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(G33), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(n996), .B(G27), .Z(n999) );
  XNOR2_X1 U1090 ( .A(n997), .B(G32), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT53), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT117), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(G29), .A2(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(G11), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT125), .B(n1016), .Z(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  XOR2_X1 U1105 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

