//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT95), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G71gat), .B(G78gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT21), .ZN(new_n207));
  NAND2_X1  g006(.A1(G231gat), .A2(G233gat), .ZN(new_n208));
  XOR2_X1   g007(.A(new_n207), .B(new_n208), .Z(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n205), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n204), .B(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n212), .A2(KEYINPUT96), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(KEYINPUT96), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT21), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216));
  INV_X1    g015(.A(G1gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(KEYINPUT16), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G1gat), .B2(new_n216), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(G8gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n215), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n210), .B(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT97), .B(G183gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G155gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n226), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G190gat), .B(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G43gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(G50gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(G50gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT15), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT90), .B(G50gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT91), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n241), .A3(new_n233), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n234), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT15), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n237), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G29gat), .ZN(new_n246));
  INV_X1    g045(.A(G36gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT14), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT14), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G29gat), .B2(G36gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n248), .B(new_n250), .C1(new_n246), .C2(new_n247), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n236), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256));
  INV_X1    g055(.A(G85gat), .ZN(new_n257));
  INV_X1    g056(.A(G92gat), .ZN(new_n258));
  AOI22_X1  g057(.A1(KEYINPUT8), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n257), .B2(new_n258), .ZN(new_n261));
  NAND4_X1  g060(.A1(KEYINPUT99), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G99gat), .B(G106gat), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n263), .B(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n255), .A2(new_n266), .B1(KEYINPUT41), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT17), .B1(new_n252), .B2(new_n254), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT17), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n270), .B(new_n253), .C1(new_n245), .C2(new_n251), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n266), .B(KEYINPUT100), .Z(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G134gat), .ZN(new_n275));
  INV_X1    g074(.A(G134gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n268), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n232), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n267), .A2(KEYINPUT41), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT98), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G162gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n275), .A2(new_n232), .A3(new_n277), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n279), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n279), .B2(new_n283), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n230), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(G211gat), .A2(G218gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(G211gat), .A2(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(G197gat), .A2(G204gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G183gat), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT24), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT25), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OR3_X1    g115(.A1(new_n304), .A2(new_n302), .A3(KEYINPUT24), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n306), .A2(new_n310), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n306), .A2(new_n321), .A3(new_n316), .A4(new_n317), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n304), .A2(new_n302), .A3(KEYINPUT24), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n304), .A2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n302), .A2(G183gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(KEYINPUT24), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(KEYINPUT65), .A3(new_n316), .A4(new_n310), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT66), .A2(KEYINPUT27), .A3(G183gat), .ZN(new_n334));
  AND2_X1   g133(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n302), .B(new_n334), .C1(new_n335), .C2(KEYINPUT27), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n333), .B1(new_n336), .B2(new_n326), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n321), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n312), .A2(new_n313), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT26), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n337), .A2(new_n340), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n331), .A2(new_n332), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n331), .A2(new_n344), .B1(new_n346), .B2(new_n332), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n301), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n346), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n332), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n300), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n353), .A3(KEYINPUT71), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n351), .A2(new_n355), .A3(new_n352), .A4(new_n300), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AND4_X1   g162(.A1(KEYINPUT75), .A2(new_n357), .A3(KEYINPUT30), .A4(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n354), .B2(new_n356), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT75), .B1(new_n365), .B2(KEYINPUT30), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n363), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n357), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n354), .A2(KEYINPUT72), .A3(new_n356), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n362), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n367), .A2(KEYINPUT84), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n363), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n365), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n374), .A2(new_n378), .A3(new_n370), .A4(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT76), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G155gat), .ZN(new_n386));
  INV_X1    g185(.A(G162gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G148gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G141gat), .ZN(new_n393));
  INV_X1    g192(.A(G141gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G148gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n390), .A2(KEYINPUT2), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n385), .A2(new_n391), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G141gat), .B(G148gat), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n390), .B(new_n388), .C1(new_n399), .C2(KEYINPUT2), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n402));
  XNOR2_X1  g201(.A(G113gat), .B(G120gat), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(KEYINPUT1), .ZN(new_n404));
  INV_X1    g203(.A(G127gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT1), .ZN(new_n406));
  INV_X1    g205(.A(G113gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(G120gat), .ZN(new_n408));
  INV_X1    g207(.A(G120gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(G113gat), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n406), .B(new_n276), .C1(new_n408), .C2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n404), .A2(new_n405), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n404), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n401), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n411), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G127gat), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n404), .A2(new_n405), .A3(new_n411), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n400), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT85), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT85), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT78), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n398), .A2(new_n427), .A3(new_n400), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n398), .B2(new_n400), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n412), .A2(new_n413), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n398), .A2(new_n433), .A3(new_n400), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT77), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT77), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n398), .A2(new_n400), .A3(new_n436), .A4(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n418), .A2(KEYINPUT3), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n431), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n416), .A2(new_n417), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n425), .B1(new_n443), .B2(new_n422), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT39), .B(new_n424), .C1(new_n444), .C2(new_n423), .ZN(new_n445));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G85gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT0), .B(G57gat), .ZN(new_n448));
  XOR2_X1   g247(.A(new_n447), .B(new_n448), .Z(new_n449));
  AND3_X1   g248(.A1(new_n432), .A2(new_n440), .A3(new_n442), .ZN(new_n450));
  OR3_X1    g249(.A1(new_n450), .A2(KEYINPUT39), .A3(new_n421), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n422), .B1(new_n414), .B2(new_n426), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n441), .B(KEYINPUT4), .C1(new_n429), .C2(new_n428), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n420), .B2(new_n422), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n450), .A2(new_n455), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT86), .B1(new_n461), .B2(new_n449), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n460), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n432), .A2(new_n440), .A3(new_n455), .A4(new_n442), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  INV_X1    g265(.A(new_n449), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n445), .A2(KEYINPUT40), .A3(new_n449), .A4(new_n451), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n454), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n375), .A2(new_n382), .A3(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT83), .B(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT29), .B1(new_n295), .B2(new_n299), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n418), .B1(new_n481), .B2(KEYINPUT3), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n300), .B1(new_n438), .B2(new_n346), .ZN(new_n485));
  NAND2_X1  g284(.A1(G228gat), .A2(G233gat), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n438), .A2(new_n346), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT80), .A3(new_n301), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n430), .B1(KEYINPUT3), .B2(new_n481), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT29), .B1(new_n435), .B2(new_n437), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n300), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n487), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n475), .A2(new_n476), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n480), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n486), .ZN(new_n498));
  INV_X1    g297(.A(new_n487), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n480), .A2(new_n498), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n478), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n499), .A3(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(new_n479), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n480), .A3(new_n496), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n504), .A3(new_n477), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n372), .A2(KEYINPUT37), .A3(new_n373), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT37), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n357), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n362), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT38), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT38), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n348), .A2(new_n353), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n363), .B1(new_n514), .B2(KEYINPUT37), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n516), .A2(KEYINPUT87), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n365), .B1(new_n516), .B2(KEYINPUT87), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n467), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n463), .A2(new_n464), .A3(new_n449), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT79), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n463), .A2(KEYINPUT79), .A3(new_n464), .A4(new_n449), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n520), .B1(new_n526), .B2(new_n469), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n512), .A2(new_n517), .A3(new_n518), .A4(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n472), .A2(new_n507), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n465), .A2(new_n467), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(new_n530), .A3(new_n524), .A4(new_n525), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(new_n519), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n367), .A2(new_n532), .A3(new_n370), .A4(new_n374), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n349), .A2(new_n441), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n331), .A2(new_n431), .A3(new_n344), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT34), .ZN(new_n538));
  INV_X1    g337(.A(G227gat), .ZN(new_n539));
  INV_X1    g338(.A(G233gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n537), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n538), .B1(new_n537), .B2(new_n542), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G43gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(G71gat), .B(G99gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n541), .A3(new_n536), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n535), .A2(KEYINPUT69), .A3(new_n541), .A4(new_n536), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT33), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n550), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT70), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n559), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n560), .A2(KEYINPUT33), .A3(new_n561), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n556), .B(new_n562), .C1(new_n553), .C2(new_n554), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n547), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n562), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(KEYINPUT32), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n553), .A2(new_n554), .B1(new_n556), .B2(KEYINPUT33), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n566), .B(new_n546), .C1(new_n567), .C2(new_n550), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n529), .A2(new_n534), .A3(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n501), .A2(new_n505), .A3(new_n568), .A4(new_n564), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT35), .B1(new_n533), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT88), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n375), .A2(new_n382), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n506), .A2(new_n527), .A3(new_n569), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT35), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT88), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n580), .B(KEYINPUT35), .C1(new_n533), .C2(new_n573), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n287), .B1(new_n572), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n584));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT12), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n221), .B(new_n253), .C1(new_n245), .C2(new_n251), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT92), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n269), .A2(new_n222), .A3(new_n271), .ZN(new_n592));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT93), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT18), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n591), .A2(new_n592), .A3(new_n597), .A4(new_n593), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n589), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n591), .B1(new_n255), .B2(new_n221), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n593), .B(KEYINPUT13), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n594), .A2(new_n596), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n601), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G230gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n540), .ZN(new_n610));
  INV_X1    g409(.A(new_n266), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n265), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n613), .B2(new_n212), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n206), .B(new_n266), .C1(new_n612), .C2(new_n265), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT10), .B(new_n266), .C1(new_n213), .C2(new_n214), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n610), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI211_X1 g418(.A(new_n609), .B(new_n540), .C1(new_n614), .C2(new_n616), .ZN(new_n620));
  OAI21_X1  g419(.A(KEYINPUT102), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n583), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n532), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT103), .B(G1gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(G1324gat));
  INV_X1    g430(.A(new_n576), .ZN(new_n632));
  NAND2_X1  g431(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n583), .A2(new_n627), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(KEYINPUT104), .B(new_n637), .C1(new_n634), .C2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n636), .A2(new_n637), .ZN(new_n644));
  OAI21_X1  g443(.A(G8gat), .B1(new_n628), .B2(new_n576), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT104), .B1(new_n636), .B2(new_n637), .ZN(new_n647));
  INV_X1    g446(.A(new_n641), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n644), .B(new_n645), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT105), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n628), .A2(new_n652), .A3(new_n571), .ZN(new_n653));
  INV_X1    g452(.A(new_n569), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n583), .A2(new_n627), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT106), .Z(G1326gat));
  NAND3_X1  g456(.A1(new_n583), .A2(new_n627), .A3(new_n506), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  AOI21_X1  g460(.A(new_n286), .B1(new_n572), .B2(new_n582), .ZN(new_n662));
  INV_X1    g461(.A(new_n230), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n662), .A2(new_n627), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n532), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n246), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT45), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n572), .A2(new_n582), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n284), .A2(new_n285), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n230), .B(KEYINPUT108), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n672), .A2(new_n627), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n532), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n667), .A2(new_n676), .ZN(G1328gat));
  NAND3_X1  g476(.A1(new_n664), .A2(new_n247), .A3(new_n632), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT46), .ZN(new_n679));
  OAI21_X1  g478(.A(G36gat), .B1(new_n675), .B2(new_n576), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(KEYINPUT46), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1329gat));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n685));
  OAI21_X1  g484(.A(G43gat), .B1(new_n675), .B2(new_n571), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n664), .A2(new_n233), .A3(new_n654), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1330gat));
  OAI21_X1  g489(.A(new_n238), .B1(new_n675), .B2(new_n507), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n507), .A2(new_n238), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT111), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n664), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g495(.A1(new_n583), .A2(new_n626), .A3(new_n608), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n665), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n576), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(G1333gat));
  INV_X1    g504(.A(new_n571), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n698), .A2(G71gat), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(G71gat), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n697), .B2(new_n569), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT50), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT112), .B(KEYINPUT113), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n714), .B(new_n716), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n506), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g518(.A1(new_n607), .A2(new_n230), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n672), .A2(new_n626), .A3(new_n674), .A4(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(new_n257), .A3(new_n532), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n668), .A2(new_n669), .A3(new_n720), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n662), .A2(KEYINPUT51), .A3(new_n720), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(KEYINPUT114), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n662), .A2(new_n728), .A3(KEYINPUT51), .A4(new_n720), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n727), .A2(new_n665), .A3(new_n626), .A4(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n722), .B1(new_n257), .B2(new_n730), .ZN(G1336gat));
  NOR2_X1   g530(.A1(new_n576), .A2(G92gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n727), .A2(new_n626), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G92gat), .B1(new_n721), .B2(new_n576), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n726), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n626), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n735), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT115), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n662), .B(new_n671), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n745), .A2(new_n626), .A3(new_n632), .A4(new_n720), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(G92gat), .B1(new_n737), .B2(new_n739), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n743), .B(new_n744), .C1(new_n747), .C2(new_n735), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n748), .ZN(G1337gat));
  NOR2_X1   g548(.A1(new_n569), .A2(G99gat), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n727), .A2(new_n626), .A3(new_n729), .A4(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G99gat), .B1(new_n721), .B2(new_n571), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1338gat));
  OR2_X1    g552(.A1(new_n721), .A2(new_n507), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G106gat), .ZN(new_n755));
  INV_X1    g554(.A(new_n626), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n507), .A2(G106gat), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n727), .A2(new_n729), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n754), .A2(G106gat), .B1(new_n737), .B2(new_n757), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(new_n759), .ZN(G1339gat));
  OR3_X1    g561(.A1(new_n619), .A2(new_n620), .A3(new_n624), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n625), .B1(new_n619), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n617), .A2(new_n618), .A3(new_n610), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT54), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n619), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT116), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n763), .B(new_n772), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n769), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n768), .A2(KEYINPUT117), .A3(new_n769), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n771), .A2(new_n773), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n601), .A2(new_n606), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n601), .A2(new_n606), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n591), .A2(new_n592), .ZN(new_n783));
  INV_X1    g582(.A(new_n593), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT118), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT118), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n788), .C1(new_n602), .C2(new_n603), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n588), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n599), .A2(new_n589), .A3(new_n604), .A4(new_n605), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n626), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n669), .B1(new_n782), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n669), .A2(new_n794), .A3(new_n778), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n673), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n287), .A2(new_n626), .A3(new_n607), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n632), .A2(new_n532), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n573), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n608), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(new_n407), .ZN(G1340gat));
  OAI21_X1  g605(.A(G120gat), .B1(new_n804), .B2(new_n756), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n626), .A2(new_n409), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT119), .Z(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n804), .B2(new_n809), .ZN(G1341gat));
  XNOR2_X1  g609(.A(KEYINPUT68), .B(G127gat), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n804), .A2(new_n673), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n804), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n230), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n811), .B2(new_n814), .ZN(G1342gat));
  NAND2_X1  g614(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n813), .A2(new_n669), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n817), .B(new_n818), .Z(G1343gat));
  AOI21_X1  g618(.A(new_n507), .B1(new_n797), .B2(new_n799), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT120), .B1(new_n820), .B2(KEYINPUT57), .ZN(new_n821));
  INV_X1    g620(.A(new_n770), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n607), .A2(new_n822), .A3(new_n774), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n792), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n796), .B1(new_n824), .B2(new_n286), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n799), .B1(new_n825), .B2(new_n230), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(KEYINPUT57), .A3(new_n506), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT57), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n607), .A2(new_n778), .B1(new_n794), .B2(new_n626), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n795), .B1(new_n830), .B2(new_n669), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n798), .B1(new_n831), .B2(new_n673), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n828), .B(new_n829), .C1(new_n832), .C2(new_n507), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n821), .A2(new_n827), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n706), .A2(new_n632), .A3(new_n532), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n607), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G141gat), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n571), .A2(new_n506), .ZN(new_n839));
  XOR2_X1   g638(.A(new_n839), .B(KEYINPUT121), .Z(new_n840));
  NAND3_X1  g639(.A1(new_n800), .A2(new_n801), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n608), .A2(G141gat), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n838), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT58), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n847), .B(new_n844), .C1(new_n836), .C2(G141gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(G1344gat));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n850), .B(G148gat), .C1(new_n851), .C2(new_n756), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n826), .B2(new_n506), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n832), .A2(new_n829), .A3(new_n507), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n626), .B(new_n835), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(G148gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n856), .B2(new_n850), .ZN(new_n857));
  INV_X1    g656(.A(new_n841), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n392), .A3(new_n626), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1345gat));
  NOR3_X1   g659(.A1(new_n851), .A2(new_n386), .A3(new_n673), .ZN(new_n861));
  AOI21_X1  g660(.A(G155gat), .B1(new_n858), .B2(new_n230), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(G1346gat));
  OAI21_X1  g662(.A(new_n387), .B1(new_n841), .B2(new_n286), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n669), .A2(G162gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n851), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT123), .ZN(G1347gat));
  NAND2_X1  g666(.A1(new_n632), .A2(new_n532), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n573), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n800), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT124), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT124), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n312), .A3(new_n607), .ZN(new_n874));
  OAI21_X1  g673(.A(G169gat), .B1(new_n870), .B2(new_n608), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1348gat));
  NOR3_X1   g675(.A1(new_n870), .A2(new_n313), .A3(new_n756), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n873), .A2(new_n626), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n313), .ZN(G1349gat));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n870), .A2(new_n880), .A3(new_n673), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n870), .B2(new_n673), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(G183gat), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n800), .A2(new_n230), .A3(new_n338), .A4(new_n869), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n870), .B2(new_n286), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT61), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n871), .A2(new_n302), .A3(new_n669), .A4(new_n872), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(G1351gat));
  NOR2_X1   g692(.A1(new_n868), .A2(new_n706), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT127), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n853), .B2(new_n854), .ZN(new_n896));
  OAI21_X1  g695(.A(G197gat), .B1(new_n896), .B2(new_n608), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n820), .A2(new_n894), .ZN(new_n898));
  INV_X1    g697(.A(G197gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n607), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1352gat));
  INV_X1    g700(.A(G204gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n626), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT62), .Z(new_n904));
  OAI211_X1 g703(.A(new_n626), .B(new_n895), .C1(new_n853), .C2(new_n854), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G204gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1353gat));
  INV_X1    g706(.A(G211gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n898), .A2(new_n908), .A3(new_n230), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n230), .B(new_n895), .C1(new_n853), .C2(new_n854), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n910), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT63), .B1(new_n910), .B2(G211gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(G1354gat));
  OAI21_X1  g712(.A(G218gat), .B1(new_n896), .B2(new_n286), .ZN(new_n914));
  INV_X1    g713(.A(G218gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n915), .A3(new_n669), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1355gat));
endmodule


