

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(n527), .A2(n567), .ZN(n758) );
  BUF_X2 U556 ( .A(n758), .Z(n787) );
  INV_X1 U557 ( .A(n895), .ZN(n1001) );
  NAND2_X1 U558 ( .A1(n552), .A2(KEYINPUT29), .ZN(n553) );
  AND2_X1 U559 ( .A1(n555), .A2(n556), .ZN(n554) );
  NOR2_X1 U560 ( .A1(n557), .A2(n524), .ZN(n556) );
  XNOR2_X1 U561 ( .A(n756), .B(KEYINPUT97), .ZN(n766) );
  NOR2_X1 U562 ( .A1(n787), .A2(n1026), .ZN(n760) );
  AND2_X1 U563 ( .A1(n564), .A2(n563), .ZN(n562) );
  XNOR2_X1 U564 ( .A(n648), .B(n647), .ZN(n895) );
  NOR2_X2 U565 ( .A1(n602), .A2(n601), .ZN(G160) );
  AND2_X2 U566 ( .A1(n538), .A2(G2104), .ZN(n743) );
  NOR2_X2 U567 ( .A1(n691), .A2(n582), .ZN(n705) );
  INV_X1 U568 ( .A(G2105), .ZN(n538) );
  NAND2_X1 U569 ( .A1(n832), .A2(n575), .ZN(n547) );
  NAND2_X1 U570 ( .A1(n565), .A2(n572), .ZN(n564) );
  NOR2_X1 U571 ( .A1(n749), .A2(n751), .ZN(n565) );
  NOR2_X1 U572 ( .A1(n763), .A2(n996), .ZN(n764) );
  AND2_X1 U573 ( .A1(n545), .A2(n542), .ZN(n541) );
  NOR2_X1 U574 ( .A1(n544), .A2(n543), .ZN(n542) );
  INV_X1 U575 ( .A(n1013), .ZN(n543) );
  AND2_X1 U576 ( .A1(n566), .A2(n569), .ZN(n568) );
  NAND2_X1 U577 ( .A1(KEYINPUT64), .A2(G1384), .ZN(n569) );
  NOR2_X1 U578 ( .A1(n573), .A2(n576), .ZN(n645) );
  NAND2_X1 U579 ( .A1(n536), .A2(KEYINPUT88), .ZN(n535) );
  NAND2_X1 U580 ( .A1(G102), .A2(G2104), .ZN(n536) );
  NOR2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n530) );
  INV_X1 U582 ( .A(G102), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n533), .A2(G2104), .ZN(n532) );
  NAND2_X1 U584 ( .A1(n596), .A2(n598), .ZN(n597) );
  INV_X1 U585 ( .A(G2104), .ZN(n596) );
  INV_X1 U586 ( .A(KEYINPUT98), .ZN(n769) );
  NOR2_X1 U587 ( .A1(n779), .A2(n781), .ZN(n557) );
  NOR2_X1 U588 ( .A1(n827), .A2(n828), .ZN(n544) );
  INV_X1 U589 ( .A(n857), .ZN(n567) );
  INV_X1 U590 ( .A(G1384), .ZN(n571) );
  NAND2_X1 U591 ( .A1(n541), .A2(n539), .ZN(n836) );
  NAND2_X1 U592 ( .A1(n540), .A2(KEYINPUT106), .ZN(n539) );
  INV_X1 U593 ( .A(KEYINPUT88), .ZN(n533) );
  AND2_X1 U594 ( .A1(n646), .A2(n645), .ZN(n648) );
  INV_X1 U595 ( .A(KEYINPUT1), .ZN(n583) );
  AND2_X1 U596 ( .A1(n537), .A2(n535), .ZN(n534) );
  INV_X1 U597 ( .A(KEYINPUT23), .ZN(n592) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  OR2_X1 U599 ( .A1(G171), .A2(n793), .ZN(n522) );
  OR2_X1 U600 ( .A1(G168), .A2(n792), .ZN(n523) );
  AND2_X1 U601 ( .A1(G171), .A2(n793), .ZN(n524) );
  OR2_X1 U602 ( .A1(n840), .A2(n839), .ZN(n525) );
  NOR2_X1 U603 ( .A1(n821), .A2(n840), .ZN(n526) );
  AND2_X1 U604 ( .A1(n562), .A2(n568), .ZN(n527) );
  AND2_X1 U605 ( .A1(n872), .A2(n871), .ZN(n528) );
  NAND2_X1 U606 ( .A1(n534), .A2(n529), .ZN(n746) );
  NAND2_X1 U607 ( .A1(n530), .A2(n538), .ZN(n529) );
  NAND2_X1 U608 ( .A1(G2105), .A2(KEYINPUT88), .ZN(n537) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n545) );
  INV_X1 U610 ( .A(n547), .ZN(n540) );
  AND2_X1 U611 ( .A1(n827), .A2(n828), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n874) );
  INV_X1 U613 ( .A(KEYINPUT110), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n550), .A2(n528), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n551), .A2(n525), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n837), .B(KEYINPUT109), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n523), .A2(n522), .ZN(n560) );
  AND2_X1 U618 ( .A1(n779), .A2(n781), .ZN(n558) );
  INV_X1 U619 ( .A(n780), .ZN(n552) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n558), .A2(n780), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n561), .A2(n559), .ZN(n796) );
  XNOR2_X1 U623 ( .A(n560), .B(n794), .ZN(n559) );
  INV_X1 U624 ( .A(n750), .ZN(n572) );
  NAND2_X1 U625 ( .A1(n750), .A2(n570), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n749), .A2(n570), .ZN(n566) );
  NOR2_X1 U627 ( .A1(n750), .A2(n749), .ZN(G164) );
  AND2_X1 U628 ( .A1(n751), .A2(n571), .ZN(n570) );
  AND2_X1 U629 ( .A1(G2104), .A2(G2105), .ZN(n925) );
  XNOR2_X1 U630 ( .A(n796), .B(n795), .ZN(n814) );
  XOR2_X1 U631 ( .A(KEYINPUT70), .B(n644), .Z(n573) );
  NAND2_X1 U632 ( .A1(n1011), .A2(n819), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n574), .A2(n820), .ZN(n575) );
  AND2_X1 U634 ( .A1(G54), .A2(n710), .ZN(n576) );
  INV_X2 U635 ( .A(G2105), .ZN(n598) );
  INV_X1 U636 ( .A(KEYINPUT26), .ZN(n759) );
  NAND2_X1 U637 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U638 ( .A(KEYINPUT30), .B(KEYINPUT99), .ZN(n790) );
  INV_X1 U639 ( .A(KEYINPUT29), .ZN(n781) );
  INV_X1 U640 ( .A(KEYINPUT101), .ZN(n795) );
  INV_X1 U641 ( .A(KEYINPUT106), .ZN(n828) );
  NAND2_X1 U642 ( .A1(n702), .A2(G66), .ZN(n641) );
  XNOR2_X1 U643 ( .A(KEYINPUT15), .B(KEYINPUT71), .ZN(n647) );
  NOR2_X1 U644 ( .A1(G543), .A2(G651), .ZN(n701) );
  NAND2_X1 U645 ( .A1(G89), .A2(n701), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT72), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  XOR2_X1 U648 ( .A(G543), .B(KEYINPUT0), .Z(n691) );
  INV_X1 U649 ( .A(G651), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G76), .A2(n705), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U652 ( .A(n581), .B(KEYINPUT5), .ZN(n590) );
  NOR2_X1 U653 ( .A1(G543), .A2(n582), .ZN(n584) );
  XNOR2_X2 U654 ( .A(n584), .B(n583), .ZN(n702) );
  NAND2_X1 U655 ( .A1(n702), .A2(G63), .ZN(n585) );
  XOR2_X1 U656 ( .A(KEYINPUT73), .B(n585), .Z(n587) );
  NOR2_X2 U657 ( .A1(G651), .A2(n691), .ZN(n710) );
  NAND2_X1 U658 ( .A1(n710), .A2(G51), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U660 ( .A(KEYINPUT6), .B(n588), .Z(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n591), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U663 ( .A1(G101), .A2(n743), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(n592), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n925), .A2(G113), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n602) );
  XNOR2_X2 U667 ( .A(n597), .B(KEYINPUT17), .ZN(n744) );
  NAND2_X1 U668 ( .A1(n744), .A2(G137), .ZN(n600) );
  NOR2_X4 U669 ( .A1(n598), .A2(G2104), .ZN(n926) );
  NAND2_X1 U670 ( .A1(G125), .A2(n926), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT111), .B(G2435), .Z(n604) );
  XNOR2_X1 U673 ( .A(G2430), .B(G2438), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(n611) );
  XOR2_X1 U675 ( .A(G2446), .B(G2454), .Z(n606) );
  XNOR2_X1 U676 ( .A(G2451), .B(G2443), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n607) );
  XOR2_X1 U678 ( .A(n607), .B(G2427), .Z(n609) );
  XNOR2_X1 U679 ( .A(G1341), .B(G1348), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n612) );
  AND2_X1 U682 ( .A1(n612), .A2(G14), .ZN(G401) );
  NAND2_X1 U683 ( .A1(G77), .A2(n705), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G90), .A2(n701), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U686 ( .A(KEYINPUT9), .B(n615), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n710), .A2(G52), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G64), .A2(n702), .ZN(n616) );
  AND2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(G301) );
  INV_X1 U691 ( .A(G301), .ZN(G171) );
  AND2_X1 U692 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U693 ( .A(G57), .ZN(G237) );
  INV_X1 U694 ( .A(G132), .ZN(G219) );
  INV_X1 U695 ( .A(G82), .ZN(G220) );
  NAND2_X1 U696 ( .A1(G75), .A2(n705), .ZN(n621) );
  NAND2_X1 U697 ( .A1(G88), .A2(n701), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G62), .A2(n702), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT81), .B(n622), .Z(n624) );
  NAND2_X1 U701 ( .A1(n710), .A2(G50), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n626), .A2(n625), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G7), .A2(G661), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT66), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT10), .B(n628), .ZN(G223) );
  INV_X1 U707 ( .A(G223), .ZN(n889) );
  NAND2_X1 U708 ( .A1(n889), .A2(G567), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT11), .B(n629), .Z(G234) );
  NAND2_X1 U710 ( .A1(n701), .A2(G81), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT12), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G68), .A2(n705), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT13), .B(n633), .Z(n637) );
  NAND2_X1 U715 ( .A1(G56), .A2(n702), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT67), .ZN(n635) );
  XNOR2_X1 U717 ( .A(n635), .B(KEYINPUT14), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U719 ( .A1(n710), .A2(G43), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n996) );
  INV_X1 U721 ( .A(G860), .ZN(n659) );
  OR2_X1 U722 ( .A1(n996), .A2(n659), .ZN(G153) );
  NAND2_X1 U723 ( .A1(G301), .A2(G868), .ZN(n640) );
  XNOR2_X1 U724 ( .A(n640), .B(KEYINPUT68), .ZN(n650) );
  INV_X1 U725 ( .A(G868), .ZN(n713) );
  NAND2_X1 U726 ( .A1(G92), .A2(n701), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n643), .B(KEYINPUT69), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n705), .A2(G79), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n713), .A2(n1001), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G284) );
  NAND2_X1 U732 ( .A1(G53), .A2(n710), .ZN(n652) );
  NAND2_X1 U733 ( .A1(G65), .A2(n702), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G78), .A2(n705), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G91), .A2(n701), .ZN(n653) );
  NAND2_X1 U737 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U738 ( .A1(n656), .A2(n655), .ZN(n1004) );
  INV_X1 U739 ( .A(n1004), .ZN(G299) );
  NOR2_X1 U740 ( .A1(G286), .A2(n713), .ZN(n658) );
  NOR2_X1 U741 ( .A1(G868), .A2(G299), .ZN(n657) );
  NOR2_X1 U742 ( .A1(n658), .A2(n657), .ZN(G297) );
  NAND2_X1 U743 ( .A1(n659), .A2(G559), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n660), .A2(n895), .ZN(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(KEYINPUT16), .ZN(n662) );
  XNOR2_X1 U746 ( .A(KEYINPUT74), .B(n662), .ZN(G148) );
  NOR2_X1 U747 ( .A1(G868), .A2(n996), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n895), .A2(G868), .ZN(n663) );
  NOR2_X1 U749 ( .A1(G559), .A2(n663), .ZN(n664) );
  NOR2_X1 U750 ( .A1(n665), .A2(n664), .ZN(G282) );
  NAND2_X1 U751 ( .A1(G99), .A2(n743), .ZN(n667) );
  NAND2_X1 U752 ( .A1(G111), .A2(n925), .ZN(n666) );
  NAND2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n674) );
  BUF_X1 U754 ( .A(n744), .Z(n929) );
  NAND2_X1 U755 ( .A1(n929), .A2(G135), .ZN(n668) );
  XNOR2_X1 U756 ( .A(KEYINPUT75), .B(n668), .ZN(n671) );
  NAND2_X1 U757 ( .A1(n926), .A2(G123), .ZN(n669) );
  XOR2_X1 U758 ( .A(KEYINPUT18), .B(n669), .Z(n670) );
  NOR2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U760 ( .A(KEYINPUT76), .B(n672), .Z(n673) );
  NOR2_X1 U761 ( .A1(n674), .A2(n673), .ZN(n976) );
  XNOR2_X1 U762 ( .A(n976), .B(G2096), .ZN(n676) );
  INV_X1 U763 ( .A(G2100), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n676), .A2(n675), .ZN(G156) );
  NAND2_X1 U765 ( .A1(G93), .A2(n701), .ZN(n678) );
  NAND2_X1 U766 ( .A1(G67), .A2(n702), .ZN(n677) );
  NAND2_X1 U767 ( .A1(n678), .A2(n677), .ZN(n681) );
  NAND2_X1 U768 ( .A1(G80), .A2(n705), .ZN(n679) );
  XNOR2_X1 U769 ( .A(KEYINPUT79), .B(n679), .ZN(n680) );
  NOR2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U771 ( .A1(n710), .A2(G55), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n683), .A2(n682), .ZN(n721) );
  XNOR2_X1 U773 ( .A(KEYINPUT78), .B(n996), .ZN(n685) );
  NAND2_X1 U774 ( .A1(G559), .A2(n895), .ZN(n684) );
  XOR2_X1 U775 ( .A(KEYINPUT77), .B(n684), .Z(n724) );
  XNOR2_X1 U776 ( .A(n685), .B(n724), .ZN(n686) );
  NOR2_X1 U777 ( .A1(G860), .A2(n686), .ZN(n687) );
  XOR2_X1 U778 ( .A(n721), .B(n687), .Z(G145) );
  NAND2_X1 U779 ( .A1(G49), .A2(n710), .ZN(n689) );
  NAND2_X1 U780 ( .A1(G74), .A2(G651), .ZN(n688) );
  NAND2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U782 ( .A1(n702), .A2(n690), .ZN(n693) );
  NAND2_X1 U783 ( .A1(n691), .A2(G87), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n693), .A2(n692), .ZN(G288) );
  NAND2_X1 U785 ( .A1(G72), .A2(n705), .ZN(n695) );
  NAND2_X1 U786 ( .A1(G85), .A2(n701), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n698) );
  NAND2_X1 U788 ( .A1(G60), .A2(n702), .ZN(n696) );
  XNOR2_X1 U789 ( .A(KEYINPUT65), .B(n696), .ZN(n697) );
  NOR2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n710), .A2(G47), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(G290) );
  NAND2_X1 U793 ( .A1(G86), .A2(n701), .ZN(n704) );
  NAND2_X1 U794 ( .A1(G61), .A2(n702), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U796 ( .A1(n705), .A2(G73), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT2), .B(n706), .Z(n707) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U799 ( .A(n709), .B(KEYINPUT80), .ZN(n712) );
  NAND2_X1 U800 ( .A1(G48), .A2(n710), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n712), .A2(n711), .ZN(G305) );
  AND2_X1 U802 ( .A1(n713), .A2(n721), .ZN(n714) );
  XNOR2_X1 U803 ( .A(n714), .B(KEYINPUT85), .ZN(n728) );
  XNOR2_X1 U804 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n716) );
  XNOR2_X1 U805 ( .A(n996), .B(KEYINPUT83), .ZN(n715) );
  XNOR2_X1 U806 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n1004), .B(n717), .ZN(n719) );
  XNOR2_X1 U808 ( .A(G288), .B(G166), .ZN(n718) );
  XNOR2_X1 U809 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n720), .B(G290), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U812 ( .A(n723), .B(G305), .ZN(n894) );
  XNOR2_X1 U813 ( .A(n894), .B(KEYINPUT84), .ZN(n725) );
  XNOR2_X1 U814 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U815 ( .A1(G868), .A2(n726), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(G295) );
  NAND2_X1 U817 ( .A1(G2084), .A2(G2078), .ZN(n729) );
  XOR2_X1 U818 ( .A(KEYINPUT20), .B(n729), .Z(n730) );
  NAND2_X1 U819 ( .A1(G2090), .A2(n730), .ZN(n731) );
  XNOR2_X1 U820 ( .A(KEYINPUT21), .B(n731), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(G2072), .ZN(n733) );
  XNOR2_X1 U822 ( .A(KEYINPUT86), .B(n733), .ZN(G158) );
  XNOR2_X1 U823 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U824 ( .A1(G220), .A2(G219), .ZN(n734) );
  XOR2_X1 U825 ( .A(KEYINPUT22), .B(n734), .Z(n735) );
  NOR2_X1 U826 ( .A1(G218), .A2(n735), .ZN(n736) );
  NAND2_X1 U827 ( .A1(G96), .A2(n736), .ZN(n942) );
  NAND2_X1 U828 ( .A1(n942), .A2(G2106), .ZN(n740) );
  NAND2_X1 U829 ( .A1(G69), .A2(G120), .ZN(n737) );
  NOR2_X1 U830 ( .A1(G237), .A2(n737), .ZN(n738) );
  NAND2_X1 U831 ( .A1(G108), .A2(n738), .ZN(n943) );
  NAND2_X1 U832 ( .A1(n943), .A2(G567), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n944) );
  NAND2_X1 U834 ( .A1(G661), .A2(G483), .ZN(n741) );
  NOR2_X1 U835 ( .A1(n944), .A2(n741), .ZN(n742) );
  XOR2_X1 U836 ( .A(KEYINPUT87), .B(n742), .Z(n893) );
  NAND2_X1 U837 ( .A1(n893), .A2(G36), .ZN(G176) );
  INV_X1 U838 ( .A(G166), .ZN(G303) );
  NAND2_X1 U839 ( .A1(n744), .A2(G138), .ZN(n745) );
  NAND2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U841 ( .A1(G114), .A2(n925), .ZN(n748) );
  NAND2_X1 U842 ( .A1(n926), .A2(G126), .ZN(n747) );
  NAND2_X1 U843 ( .A1(n748), .A2(n747), .ZN(n749) );
  INV_X1 U844 ( .A(KEYINPUT64), .ZN(n751) );
  NAND2_X1 U845 ( .A1(G160), .A2(G40), .ZN(n857) );
  NAND2_X1 U846 ( .A1(n758), .A2(G1348), .ZN(n753) );
  XNOR2_X1 U847 ( .A(n753), .B(KEYINPUT96), .ZN(n755) );
  INV_X1 U848 ( .A(n758), .ZN(n807) );
  NAND2_X1 U849 ( .A1(n807), .A2(G2067), .ZN(n754) );
  INV_X1 U850 ( .A(n766), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n757), .A2(n1001), .ZN(n765) );
  INV_X1 U852 ( .A(G1996), .ZN(n1026) );
  XNOR2_X1 U853 ( .A(n760), .B(n759), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n787), .A2(G1341), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U857 ( .A1(n766), .A2(n895), .ZN(n767) );
  NAND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n770) );
  XNOR2_X1 U859 ( .A(n770), .B(n769), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n807), .A2(G2072), .ZN(n771) );
  XNOR2_X1 U861 ( .A(n771), .B(KEYINPUT27), .ZN(n773) );
  AND2_X1 U862 ( .A1(G1956), .A2(n787), .ZN(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n776), .A2(n1004), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n780) );
  NOR2_X1 U866 ( .A1(n776), .A2(n1004), .ZN(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U869 ( .A(G2078), .B(KEYINPUT25), .ZN(n1025) );
  NOR2_X1 U870 ( .A1(n787), .A2(n1025), .ZN(n783) );
  AND2_X1 U871 ( .A1(n787), .A2(G1961), .ZN(n782) );
  NOR2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n793) );
  NOR2_X1 U873 ( .A1(n787), .A2(G2084), .ZN(n785) );
  INV_X1 U874 ( .A(KEYINPUT94), .ZN(n784) );
  XNOR2_X1 U875 ( .A(n785), .B(n784), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n786), .A2(G8), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G8), .A2(n787), .ZN(n840) );
  NOR2_X1 U878 ( .A1(G1966), .A2(n840), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n791) );
  XNOR2_X1 U880 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U881 ( .A(KEYINPUT100), .B(KEYINPUT31), .ZN(n794) );
  NAND2_X1 U882 ( .A1(n814), .A2(G286), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n797), .B(KEYINPUT102), .ZN(n803) );
  NOR2_X1 U884 ( .A1(G2090), .A2(n758), .ZN(n799) );
  NOR2_X1 U885 ( .A1(G1971), .A2(n840), .ZN(n798) );
  NOR2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n800), .A2(G303), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT103), .B(n801), .Z(n802) );
  NAND2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n804), .A2(G8), .ZN(n805) );
  XNOR2_X1 U891 ( .A(n805), .B(KEYINPUT32), .ZN(n817) );
  NAND2_X1 U892 ( .A1(KEYINPUT94), .A2(G1966), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n806), .A2(n758), .ZN(n812) );
  INV_X1 U894 ( .A(G2084), .ZN(n1037) );
  NAND2_X1 U895 ( .A1(KEYINPUT94), .A2(n807), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n1037), .A2(n808), .ZN(n810) );
  NAND2_X1 U897 ( .A1(KEYINPUT94), .A2(G2084), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n813), .A2(G8), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n817), .A2(n816), .ZN(n832) );
  NOR2_X1 U903 ( .A1(G288), .A2(G1976), .ZN(n818) );
  XNOR2_X1 U904 ( .A(n818), .B(KEYINPUT104), .ZN(n822) );
  INV_X1 U905 ( .A(n822), .ZN(n1011) );
  INV_X1 U906 ( .A(KEYINPUT33), .ZN(n819) );
  NOR2_X1 U907 ( .A1(G1971), .A2(G303), .ZN(n820) );
  NAND2_X1 U908 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  INV_X1 U909 ( .A(n1005), .ZN(n821) );
  NOR2_X1 U910 ( .A1(KEYINPUT33), .A2(n526), .ZN(n826) );
  NAND2_X1 U911 ( .A1(KEYINPUT33), .A2(n822), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NOR2_X1 U913 ( .A1(n840), .A2(n824), .ZN(n825) );
  NOR2_X1 U914 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U915 ( .A(G1981), .B(G305), .Z(n1013) );
  NOR2_X1 U916 ( .A1(G2090), .A2(G303), .ZN(n829) );
  XOR2_X1 U917 ( .A(KEYINPUT107), .B(n829), .Z(n830) );
  NAND2_X1 U918 ( .A1(G8), .A2(n830), .ZN(n831) );
  NAND2_X1 U919 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U920 ( .A(n833), .B(KEYINPUT108), .ZN(n834) );
  NAND2_X1 U921 ( .A1(n834), .A2(n840), .ZN(n835) );
  NAND2_X1 U922 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U923 ( .A1(G1981), .A2(G305), .ZN(n838) );
  XOR2_X1 U924 ( .A(n838), .B(KEYINPUT24), .Z(n839) );
  NAND2_X1 U925 ( .A1(G107), .A2(n925), .ZN(n842) );
  NAND2_X1 U926 ( .A1(G119), .A2(n926), .ZN(n841) );
  NAND2_X1 U927 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U928 ( .A(KEYINPUT92), .B(n843), .Z(n847) );
  NAND2_X1 U929 ( .A1(G95), .A2(n743), .ZN(n845) );
  NAND2_X1 U930 ( .A1(G131), .A2(n929), .ZN(n844) );
  AND2_X1 U931 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U932 ( .A1(n847), .A2(n846), .ZN(n918) );
  AND2_X1 U933 ( .A1(n918), .A2(G1991), .ZN(n856) );
  NAND2_X1 U934 ( .A1(G117), .A2(n925), .ZN(n849) );
  NAND2_X1 U935 ( .A1(G141), .A2(n929), .ZN(n848) );
  NAND2_X1 U936 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U937 ( .A1(n743), .A2(G105), .ZN(n850) );
  XOR2_X1 U938 ( .A(KEYINPUT38), .B(n850), .Z(n851) );
  NOR2_X1 U939 ( .A1(n852), .A2(n851), .ZN(n854) );
  NAND2_X1 U940 ( .A1(n926), .A2(G129), .ZN(n853) );
  NAND2_X1 U941 ( .A1(n854), .A2(n853), .ZN(n922) );
  AND2_X1 U942 ( .A1(n922), .A2(G1996), .ZN(n855) );
  NOR2_X1 U943 ( .A1(n856), .A2(n855), .ZN(n975) );
  NOR2_X1 U944 ( .A1(n857), .A2(n527), .ZN(n884) );
  XNOR2_X1 U945 ( .A(KEYINPUT93), .B(n884), .ZN(n858) );
  NOR2_X1 U946 ( .A1(n975), .A2(n858), .ZN(n877) );
  INV_X1 U947 ( .A(n877), .ZN(n872) );
  NAND2_X1 U948 ( .A1(n925), .A2(G116), .ZN(n859) );
  XNOR2_X1 U949 ( .A(n859), .B(KEYINPUT90), .ZN(n861) );
  NAND2_X1 U950 ( .A1(G128), .A2(n926), .ZN(n860) );
  NAND2_X1 U951 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U952 ( .A(n862), .B(KEYINPUT35), .ZN(n867) );
  NAND2_X1 U953 ( .A1(G104), .A2(n743), .ZN(n864) );
  NAND2_X1 U954 ( .A1(G140), .A2(n929), .ZN(n863) );
  NAND2_X1 U955 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U956 ( .A(KEYINPUT34), .B(n865), .Z(n866) );
  NAND2_X1 U957 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U958 ( .A(n868), .B(KEYINPUT36), .Z(n938) );
  XNOR2_X1 U959 ( .A(G2067), .B(KEYINPUT37), .ZN(n869) );
  XOR2_X1 U960 ( .A(n869), .B(KEYINPUT89), .Z(n882) );
  OR2_X1 U961 ( .A1(n938), .A2(n882), .ZN(n870) );
  XOR2_X1 U962 ( .A(KEYINPUT91), .B(n870), .Z(n880) );
  INV_X1 U963 ( .A(n880), .ZN(n981) );
  NAND2_X1 U964 ( .A1(n884), .A2(n981), .ZN(n871) );
  XNOR2_X1 U965 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U966 ( .A1(n998), .A2(n884), .ZN(n873) );
  NAND2_X1 U967 ( .A1(n874), .A2(n873), .ZN(n887) );
  NOR2_X1 U968 ( .A1(G1996), .A2(n922), .ZN(n988) );
  NOR2_X1 U969 ( .A1(G1991), .A2(n918), .ZN(n977) );
  NOR2_X1 U970 ( .A1(G1986), .A2(G290), .ZN(n875) );
  NOR2_X1 U971 ( .A1(n977), .A2(n875), .ZN(n876) );
  NOR2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U973 ( .A1(n988), .A2(n878), .ZN(n879) );
  XNOR2_X1 U974 ( .A(n879), .B(KEYINPUT39), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n881), .A2(n880), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n882), .A2(n938), .ZN(n974) );
  NAND2_X1 U977 ( .A1(n883), .A2(n974), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U979 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U980 ( .A(n888), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U981 ( .A1(G2106), .A2(n889), .ZN(G217) );
  NAND2_X1 U982 ( .A1(G15), .A2(G2), .ZN(n890) );
  XOR2_X1 U983 ( .A(KEYINPUT112), .B(n890), .Z(n891) );
  NAND2_X1 U984 ( .A1(G661), .A2(n891), .ZN(G259) );
  NAND2_X1 U985 ( .A1(G3), .A2(G1), .ZN(n892) );
  NAND2_X1 U986 ( .A1(n893), .A2(n892), .ZN(G188) );
  XOR2_X1 U987 ( .A(n894), .B(G286), .Z(n897) );
  XNOR2_X1 U988 ( .A(G171), .B(n895), .ZN(n896) );
  XNOR2_X1 U989 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U990 ( .A1(G37), .A2(n898), .ZN(G397) );
  NAND2_X1 U991 ( .A1(G124), .A2(n926), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(KEYINPUT44), .ZN(n906) );
  NAND2_X1 U993 ( .A1(G112), .A2(n925), .ZN(n901) );
  NAND2_X1 U994 ( .A1(G136), .A2(n929), .ZN(n900) );
  NAND2_X1 U995 ( .A1(n901), .A2(n900), .ZN(n904) );
  NAND2_X1 U996 ( .A1(G100), .A2(n743), .ZN(n902) );
  XNOR2_X1 U997 ( .A(KEYINPUT115), .B(n902), .ZN(n903) );
  NOR2_X1 U998 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1000 ( .A(KEYINPUT116), .B(n907), .Z(G162) );
  XOR2_X1 U1001 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n909) );
  XNOR2_X1 U1002 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n917) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n743), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n929), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n916) );
  NAND2_X1 U1007 ( .A1(G115), .A2(n925), .ZN(n913) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n926), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n914), .Z(n915) );
  NOR2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(n970) );
  XOR2_X1 U1012 ( .A(n917), .B(n970), .Z(n920) );
  XOR2_X1 U1013 ( .A(G160), .B(n918), .Z(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G162), .B(n921), .ZN(n924) );
  XOR2_X1 U1016 ( .A(G164), .B(n922), .Z(n923) );
  XNOR2_X1 U1017 ( .A(n924), .B(n923), .ZN(n937) );
  NAND2_X1 U1018 ( .A1(G118), .A2(n925), .ZN(n928) );
  NAND2_X1 U1019 ( .A1(G130), .A2(n926), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n935) );
  NAND2_X1 U1021 ( .A1(n929), .A2(G142), .ZN(n930) );
  XOR2_X1 U1022 ( .A(KEYINPUT117), .B(n930), .Z(n932) );
  NAND2_X1 U1023 ( .A1(n743), .A2(G106), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1025 ( .A(n933), .B(KEYINPUT45), .Z(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1027 ( .A(n937), .B(n936), .Z(n940) );
  XNOR2_X1 U1028 ( .A(n976), .B(n938), .ZN(n939) );
  XNOR2_X1 U1029 ( .A(n940), .B(n939), .ZN(n941) );
  NOR2_X1 U1030 ( .A1(G37), .A2(n941), .ZN(G395) );
  INV_X1 U1032 ( .A(G120), .ZN(G236) );
  INV_X1 U1033 ( .A(G96), .ZN(G221) );
  INV_X1 U1034 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(G325) );
  INV_X1 U1036 ( .A(G325), .ZN(G261) );
  INV_X1 U1037 ( .A(n944), .ZN(G319) );
  XOR2_X1 U1038 ( .A(G2100), .B(G2096), .Z(n946) );
  XNOR2_X1 U1039 ( .A(KEYINPUT42), .B(G2678), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n946), .B(n945), .ZN(n950) );
  XOR2_X1 U1041 ( .A(KEYINPUT43), .B(G2090), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n949) );
  XOR2_X1 U1044 ( .A(n950), .B(n949), .Z(n952) );
  XNOR2_X1 U1045 ( .A(G2084), .B(G2078), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(n952), .B(n951), .ZN(G227) );
  XOR2_X1 U1047 ( .A(G2474), .B(G1961), .Z(n954) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G1976), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n954), .B(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(n955), .B(KEYINPUT113), .Z(n957) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G1991), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n957), .B(n956), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G1956), .B(G1966), .Z(n959) );
  XNOR2_X1 U1054 ( .A(G1981), .B(G1971), .ZN(n958) );
  XNOR2_X1 U1055 ( .A(n959), .B(n958), .ZN(n960) );
  XOR2_X1 U1056 ( .A(n961), .B(n960), .Z(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT41), .B(KEYINPUT114), .ZN(n962) );
  XNOR2_X1 U1058 ( .A(n963), .B(n962), .ZN(G229) );
  NOR2_X1 U1059 ( .A1(G397), .A2(G395), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n964), .B(KEYINPUT120), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(G319), .A2(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(G401), .A2(n966), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(G227), .A2(G229), .ZN(n967) );
  XOR2_X1 U1064 ( .A(KEYINPUT49), .B(n967), .Z(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(G225) );
  INV_X1 U1066 ( .A(G225), .ZN(G308) );
  INV_X1 U1067 ( .A(G108), .ZN(G238) );
  INV_X1 U1068 ( .A(KEYINPUT55), .ZN(n1042) );
  XOR2_X1 U1069 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1071 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1072 ( .A(KEYINPUT50), .B(n973), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G160), .B(G2084), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT121), .B(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT51), .B(n989), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT122), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(n993), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n1042), .A2(n994), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n995), .A2(G29), .ZN(n1049) );
  XOR2_X1 U1089 ( .A(G16), .B(KEYINPUT56), .Z(n1021) );
  XNOR2_X1 U1090 ( .A(G166), .B(G1971), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1341), .B(n996), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1018) );
  XNOR2_X1 U1096 ( .A(G1956), .B(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(G1961), .B(G171), .Z(n1007) );
  XNOR2_X1 U1099 ( .A(KEYINPUT124), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G168), .B(G1966), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT57), .B(n1014), .Z(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(KEYINPUT125), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1047) );
  XNOR2_X1 U1109 ( .A(G2090), .B(G35), .ZN(n1036) );
  XOR2_X1 U1110 ( .A(G25), .B(G1991), .Z(n1022) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(G28), .ZN(n1032) );
  XNOR2_X1 U1112 ( .A(G2067), .B(G26), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(G33), .B(G2072), .ZN(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1030) );
  XOR2_X1 U1115 ( .A(n1025), .B(G27), .Z(n1028) );
  XOR2_X1 U1116 ( .A(n1026), .B(G32), .Z(n1027) );
  NOR2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1120 ( .A(KEYINPUT53), .B(n1033), .Z(n1034) );
  XNOR2_X1 U1121 ( .A(n1034), .B(KEYINPUT123), .ZN(n1035) );
  NOR2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1040) );
  XNOR2_X1 U1123 ( .A(G34), .B(KEYINPUT54), .ZN(n1038) );
  XNOR2_X1 U1124 ( .A(n1038), .B(n1037), .ZN(n1039) );
  NAND2_X1 U1125 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XNOR2_X1 U1126 ( .A(n1042), .B(n1041), .ZN(n1044) );
  INV_X1 U1127 ( .A(G29), .ZN(n1043) );
  NAND2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(G11), .A2(n1045), .ZN(n1046) );
  NOR2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1131 ( .A1(n1049), .A2(n1048), .ZN(n1074) );
  XNOR2_X1 U1132 ( .A(G1961), .B(G5), .ZN(n1050) );
  XNOR2_X1 U1133 ( .A(n1050), .B(KEYINPUT126), .ZN(n1057) );
  XNOR2_X1 U1134 ( .A(G1976), .B(G23), .ZN(n1052) );
  XNOR2_X1 U1135 ( .A(G1971), .B(G22), .ZN(n1051) );
  NOR2_X1 U1136 ( .A1(n1052), .A2(n1051), .ZN(n1054) );
  XOR2_X1 U1137 ( .A(G1986), .B(G24), .Z(n1053) );
  NAND2_X1 U1138 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  XNOR2_X1 U1139 ( .A(KEYINPUT58), .B(n1055), .ZN(n1056) );
  NOR2_X1 U1140 ( .A1(n1057), .A2(n1056), .ZN(n1068) );
  XNOR2_X1 U1141 ( .A(KEYINPUT59), .B(G1348), .ZN(n1058) );
  XNOR2_X1 U1142 ( .A(n1058), .B(G4), .ZN(n1065) );
  XNOR2_X1 U1143 ( .A(G1956), .B(G20), .ZN(n1063) );
  XNOR2_X1 U1144 ( .A(G1981), .B(G6), .ZN(n1060) );
  XNOR2_X1 U1145 ( .A(G1341), .B(G19), .ZN(n1059) );
  NOR2_X1 U1146 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
  XNOR2_X1 U1147 ( .A(KEYINPUT127), .B(n1061), .ZN(n1062) );
  NOR2_X1 U1148 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  NAND2_X1 U1149 ( .A1(n1065), .A2(n1064), .ZN(n1066) );
  XOR2_X1 U1150 ( .A(KEYINPUT60), .B(n1066), .Z(n1067) );
  NAND2_X1 U1151 ( .A1(n1068), .A2(n1067), .ZN(n1070) );
  XNOR2_X1 U1152 ( .A(G21), .B(G1966), .ZN(n1069) );
  NOR2_X1 U1153 ( .A1(n1070), .A2(n1069), .ZN(n1071) );
  XOR2_X1 U1154 ( .A(KEYINPUT61), .B(n1071), .Z(n1072) );
  NOR2_X1 U1155 ( .A1(G16), .A2(n1072), .ZN(n1073) );
  NOR2_X1 U1156 ( .A1(n1074), .A2(n1073), .ZN(n1075) );
  XNOR2_X1 U1157 ( .A(n1075), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1158 ( .A(G311), .ZN(G150) );
endmodule

