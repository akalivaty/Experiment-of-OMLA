

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596;

  NOR2_X1 U328 ( .A1(n479), .A2(n504), .ZN(n369) );
  XNOR2_X1 U329 ( .A(n432), .B(n431), .ZN(n440) );
  XNOR2_X1 U330 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U331 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  XOR2_X1 U332 ( .A(G120GAT), .B(G204GAT), .Z(n296) );
  AND2_X1 U333 ( .A1(n540), .A2(n580), .ZN(n371) );
  XNOR2_X1 U334 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n475) );
  XNOR2_X1 U335 ( .A(n476), .B(n475), .ZN(n541) );
  XNOR2_X1 U336 ( .A(n430), .B(n296), .ZN(n431) );
  XNOR2_X1 U337 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U338 ( .A(n382), .B(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U339 ( .A(n440), .B(n439), .ZN(n463) );
  XOR2_X1 U340 ( .A(KEYINPUT95), .B(n370), .Z(n580) );
  XNOR2_X1 U341 ( .A(n484), .B(KEYINPUT122), .ZN(n576) );
  XOR2_X1 U342 ( .A(n333), .B(n332), .Z(n548) );
  XNOR2_X1 U343 ( .A(n487), .B(G190GAT), .ZN(n488) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n461) );
  XNOR2_X1 U345 ( .A(n489), .B(n488), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n298) );
  XNOR2_X1 U348 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n312) );
  XOR2_X1 U350 ( .A(G155GAT), .B(G162GAT), .Z(n300) );
  XNOR2_X1 U351 ( .A(G127GAT), .B(G148GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U353 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n302) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n304), .B(n303), .Z(n310) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n305) );
  XNOR2_X1 U358 ( .A(n305), .B(KEYINPUT2), .ZN(n354) );
  XOR2_X1 U359 ( .A(G85GAT), .B(n354), .Z(n307) );
  NAND2_X1 U360 ( .A1(G225GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(G29GAT), .B(n308), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U365 ( .A(KEYINPUT0), .B(G134GAT), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT81), .B(G120GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(n315), .ZN(n332) );
  XOR2_X1 U369 ( .A(n316), .B(n332), .Z(n531) );
  INV_X1 U370 ( .A(n531), .ZN(n544) );
  XOR2_X1 U371 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n318) );
  XNOR2_X1 U372 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(G169GAT), .B(n319), .Z(n347) );
  XOR2_X1 U375 ( .A(KEYINPUT85), .B(G190GAT), .Z(n321) );
  XNOR2_X1 U376 ( .A(G43GAT), .B(G99GAT), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U378 ( .A(G183GAT), .B(KEYINPUT83), .Z(n323) );
  XNOR2_X1 U379 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U381 ( .A(n325), .B(n324), .Z(n330) );
  XOR2_X1 U382 ( .A(G15GAT), .B(G127GAT), .Z(n406) );
  XOR2_X1 U383 ( .A(G176GAT), .B(G71GAT), .Z(n327) );
  NAND2_X1 U384 ( .A1(G227GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n406), .B(n328), .ZN(n329) );
  XNOR2_X1 U387 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n347), .B(n331), .ZN(n333) );
  INV_X1 U389 ( .A(n548), .ZN(n504) );
  XNOR2_X1 U390 ( .A(KEYINPUT27), .B(KEYINPUT93), .ZN(n348) );
  XOR2_X1 U391 ( .A(KEYINPUT76), .B(G211GAT), .Z(n335) );
  XNOR2_X1 U392 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n409) );
  XOR2_X1 U394 ( .A(n409), .B(G92GAT), .Z(n337) );
  NAND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U397 ( .A(G36GAT), .B(G190GAT), .Z(n396) );
  XOR2_X1 U398 ( .A(n338), .B(n396), .Z(n345) );
  XOR2_X1 U399 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n340) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U402 ( .A(G218GAT), .B(KEYINPUT88), .Z(n341) );
  XOR2_X1 U403 ( .A(n342), .B(n341), .Z(n363) );
  INV_X1 U404 ( .A(n363), .ZN(n343) );
  XOR2_X1 U405 ( .A(G176GAT), .B(G64GAT), .Z(n430) );
  XOR2_X1 U406 ( .A(n343), .B(n430), .Z(n344) );
  XNOR2_X1 U407 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U408 ( .A(n347), .B(n346), .Z(n514) );
  XOR2_X1 U409 ( .A(n348), .B(n514), .Z(n540) );
  XOR2_X1 U410 ( .A(KEYINPUT86), .B(G211GAT), .Z(n350) );
  NAND2_X1 U411 ( .A1(G228GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U413 ( .A(n351), .B(KEYINPUT22), .Z(n356) );
  XOR2_X1 U414 ( .A(G78GAT), .B(G148GAT), .Z(n353) );
  XNOR2_X1 U415 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n434) );
  XNOR2_X1 U417 ( .A(n434), .B(n354), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U419 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n358) );
  XNOR2_X1 U420 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n360), .B(n359), .Z(n362) );
  XOR2_X1 U423 ( .A(G50GAT), .B(G162GAT), .Z(n397) );
  XOR2_X1 U424 ( .A(G22GAT), .B(G155GAT), .Z(n405) );
  XNOR2_X1 U425 ( .A(n397), .B(n405), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U427 ( .A(n364), .B(n363), .Z(n479) );
  XOR2_X1 U428 ( .A(n479), .B(KEYINPUT28), .Z(n517) );
  INV_X1 U429 ( .A(n517), .ZN(n546) );
  NAND2_X1 U430 ( .A1(n540), .A2(n546), .ZN(n365) );
  NOR2_X1 U431 ( .A1(n504), .A2(n365), .ZN(n366) );
  NAND2_X1 U432 ( .A1(n544), .A2(n366), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n367), .B(KEYINPUT94), .ZN(n381) );
  XNOR2_X1 U434 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U436 ( .A(KEYINPUT97), .B(n371), .ZN(n378) );
  INV_X1 U437 ( .A(n514), .ZN(n533) );
  NOR2_X1 U438 ( .A1(n548), .A2(n533), .ZN(n372) );
  XOR2_X1 U439 ( .A(KEYINPUT98), .B(n372), .Z(n373) );
  NAND2_X1 U440 ( .A1(n373), .A2(n479), .ZN(n376) );
  XNOR2_X1 U441 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n374), .B(KEYINPUT25), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  NAND2_X1 U444 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U445 ( .A1(n379), .A2(n531), .ZN(n380) );
  NAND2_X1 U446 ( .A1(n381), .A2(n380), .ZN(n382) );
  INV_X1 U447 ( .A(n497), .ZN(n420) );
  XOR2_X1 U448 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n384) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U451 ( .A(n385), .B(KEYINPUT75), .Z(n391) );
  XOR2_X1 U452 ( .A(G29GAT), .B(G43GAT), .Z(n387) );
  XNOR2_X1 U453 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n441) );
  XOR2_X1 U455 ( .A(G92GAT), .B(KEYINPUT73), .Z(n389) );
  XNOR2_X1 U456 ( .A(G99GAT), .B(G85GAT), .ZN(n388) );
  XNOR2_X1 U457 ( .A(n389), .B(n388), .ZN(n425) );
  XNOR2_X1 U458 ( .A(n441), .B(n425), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U460 ( .A(KEYINPUT9), .B(G106GAT), .Z(n393) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(G218GAT), .ZN(n392) );
  XNOR2_X1 U462 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U463 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U464 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U465 ( .A(n399), .B(n398), .Z(n573) );
  XNOR2_X1 U466 ( .A(KEYINPUT36), .B(n573), .ZN(n594) );
  XOR2_X1 U467 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n401) );
  XNOR2_X1 U468 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n418) );
  XOR2_X1 U470 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n403) );
  NAND2_X1 U471 ( .A1(G231GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U473 ( .A(G64GAT), .B(n404), .ZN(n416) );
  XOR2_X1 U474 ( .A(KEYINPUT77), .B(n405), .Z(n408) );
  XNOR2_X1 U475 ( .A(n406), .B(G78GAT), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U477 ( .A(n410), .B(n409), .Z(n414) );
  XOR2_X1 U478 ( .A(KEYINPUT69), .B(G1GAT), .Z(n453) );
  XOR2_X1 U479 ( .A(KEYINPUT70), .B(KEYINPUT13), .Z(n412) );
  XNOR2_X1 U480 ( .A(G71GAT), .B(G57GAT), .ZN(n411) );
  XNOR2_X1 U481 ( .A(n412), .B(n411), .ZN(n433) );
  XNOR2_X1 U482 ( .A(n453), .B(n433), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U484 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U485 ( .A(n418), .B(n417), .Z(n589) );
  NOR2_X1 U486 ( .A1(n594), .A2(n589), .ZN(n419) );
  NAND2_X1 U487 ( .A1(n420), .A2(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(KEYINPUT108), .B(n421), .ZN(n422) );
  XNOR2_X1 U489 ( .A(KEYINPUT37), .B(n422), .ZN(n530) );
  INV_X1 U490 ( .A(n425), .ZN(n424) );
  INV_X1 U491 ( .A(KEYINPUT71), .ZN(n423) );
  NAND2_X1 U492 ( .A1(n424), .A2(n423), .ZN(n427) );
  NAND2_X1 U493 ( .A1(n425), .A2(KEYINPUT71), .ZN(n426) );
  NAND2_X1 U494 ( .A1(n427), .A2(n426), .ZN(n429) );
  AND2_X1 U495 ( .A1(G230GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U498 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n436) );
  XNOR2_X1 U499 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n435) );
  XOR2_X1 U500 ( .A(n436), .B(n435), .Z(n437) );
  XOR2_X1 U501 ( .A(n441), .B(KEYINPUT65), .Z(n443) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U503 ( .A(n443), .B(n442), .ZN(n459) );
  XOR2_X1 U504 ( .A(KEYINPUT68), .B(G8GAT), .Z(n445) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(G113GAT), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U507 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n447) );
  XNOR2_X1 U508 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n457) );
  XOR2_X1 U511 ( .A(G22GAT), .B(G197GAT), .Z(n451) );
  XNOR2_X1 U512 ( .A(G36GAT), .B(G50GAT), .ZN(n450) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U514 ( .A(n452), .B(G141GAT), .Z(n455) );
  XNOR2_X1 U515 ( .A(G169GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U518 ( .A(n459), .B(n458), .Z(n549) );
  INV_X1 U519 ( .A(n549), .ZN(n582) );
  NOR2_X1 U520 ( .A1(n463), .A2(n582), .ZN(n498) );
  NAND2_X1 U521 ( .A1(n530), .A2(n498), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT38), .B(n460), .Z(n516) );
  NAND2_X1 U523 ( .A1(n516), .A2(n504), .ZN(n462) );
  XOR2_X1 U524 ( .A(n463), .B(KEYINPUT64), .Z(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT41), .B(n464), .Z(n575) );
  INV_X1 U526 ( .A(n575), .ZN(n551) );
  NAND2_X1 U527 ( .A1(n551), .A2(n549), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT46), .ZN(n467) );
  INV_X1 U529 ( .A(n589), .ZN(n570) );
  XOR2_X1 U530 ( .A(n570), .B(KEYINPUT113), .Z(n555) );
  INV_X1 U531 ( .A(n573), .ZN(n558) );
  AND2_X1 U532 ( .A1(n555), .A2(n573), .ZN(n466) );
  AND2_X1 U533 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U534 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n468) );
  XNOR2_X1 U535 ( .A(n469), .B(n468), .ZN(n474) );
  NOR2_X1 U536 ( .A1(n594), .A2(n570), .ZN(n470) );
  XOR2_X1 U537 ( .A(KEYINPUT45), .B(n470), .Z(n471) );
  NOR2_X1 U538 ( .A1(n463), .A2(n471), .ZN(n472) );
  NAND2_X1 U539 ( .A1(n582), .A2(n472), .ZN(n473) );
  NAND2_X1 U540 ( .A1(n474), .A2(n473), .ZN(n476) );
  NOR2_X1 U541 ( .A1(n541), .A2(n533), .ZN(n477) );
  XOR2_X1 U542 ( .A(KEYINPUT54), .B(n477), .Z(n478) );
  NOR2_X2 U543 ( .A1(n544), .A2(n478), .ZN(n581) );
  NAND2_X1 U544 ( .A1(n581), .A2(n479), .ZN(n482) );
  XOR2_X1 U545 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n480) );
  NAND2_X1 U546 ( .A1(n483), .A2(n504), .ZN(n484) );
  NOR2_X1 U547 ( .A1(n576), .A2(n582), .ZN(n486) );
  XNOR2_X1 U548 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(G1348GAT) );
  NOR2_X1 U550 ( .A1(n576), .A2(n573), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n487) );
  NOR2_X1 U552 ( .A1(n576), .A2(n555), .ZN(n492) );
  INV_X1 U553 ( .A(G183GAT), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n490), .B(KEYINPUT124), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1350GAT) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT104), .ZN(n494) );
  XOR2_X1 U558 ( .A(KEYINPUT103), .B(n494), .Z(n501) );
  NAND2_X1 U559 ( .A1(n573), .A2(n589), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n495), .B(KEYINPUT16), .ZN(n496) );
  NOR2_X1 U561 ( .A1(n497), .A2(n496), .ZN(n520) );
  NAND2_X1 U562 ( .A1(n498), .A2(n520), .ZN(n499) );
  XOR2_X1 U563 ( .A(KEYINPUT102), .B(n499), .Z(n508) );
  NAND2_X1 U564 ( .A1(n508), .A2(n544), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1324GAT) );
  XOR2_X1 U566 ( .A(G8GAT), .B(KEYINPUT105), .Z(n503) );
  NAND2_X1 U567 ( .A1(n514), .A2(n508), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(KEYINPUT35), .Z(n506) );
  NAND2_X1 U570 ( .A1(n508), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G15GAT), .B(n507), .ZN(G1326GAT) );
  XOR2_X1 U573 ( .A(G22GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U574 ( .A1(n517), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1327GAT) );
  NAND2_X1 U576 ( .A1(n516), .A2(n544), .ZN(n513) );
  XNOR2_X1 U577 ( .A(G29GAT), .B(KEYINPUT109), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT39), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(G1328GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n516), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G36GAT), .B(n515), .ZN(G1329GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G50GAT), .B(n518), .ZN(G1331GAT) );
  NOR2_X1 U584 ( .A1(n575), .A2(n549), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT110), .ZN(n529) );
  NAND2_X1 U586 ( .A1(n520), .A2(n529), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n531), .A2(n525), .ZN(n521) );
  XOR2_X1 U588 ( .A(G57GAT), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT42), .B(n522), .ZN(G1332GAT) );
  NOR2_X1 U590 ( .A1(n533), .A2(n525), .ZN(n523) );
  XOR2_X1 U591 ( .A(G64GAT), .B(n523), .Z(G1333GAT) );
  NOR2_X1 U592 ( .A1(n548), .A2(n525), .ZN(n524) );
  XOR2_X1 U593 ( .A(G71GAT), .B(n524), .Z(G1334GAT) );
  NOR2_X1 U594 ( .A1(n546), .A2(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U597 ( .A(G78GAT), .B(n528), .Z(G1335GAT) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U599 ( .A1(n531), .A2(n537), .ZN(n532) );
  XOR2_X1 U600 ( .A(G85GAT), .B(n532), .Z(G1336GAT) );
  NOR2_X1 U601 ( .A1(n533), .A2(n537), .ZN(n534) );
  XOR2_X1 U602 ( .A(KEYINPUT112), .B(n534), .Z(n535) );
  XNOR2_X1 U603 ( .A(G92GAT), .B(n535), .ZN(G1337GAT) );
  NOR2_X1 U604 ( .A1(n548), .A2(n537), .ZN(n536) );
  XOR2_X1 U605 ( .A(G99GAT), .B(n536), .Z(G1338GAT) );
  NOR2_X1 U606 ( .A1(n546), .A2(n537), .ZN(n538) );
  XOR2_X1 U607 ( .A(KEYINPUT44), .B(n538), .Z(n539) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n539), .ZN(G1339GAT) );
  INV_X1 U609 ( .A(n540), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(n545), .Z(n563) );
  NAND2_X1 U613 ( .A1(n546), .A2(n563), .ZN(n547) );
  NOR2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n559), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(G120GAT), .B(KEYINPUT49), .Z(n553) );
  NAND2_X1 U618 ( .A1(n559), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1341GAT) );
  INV_X1 U620 ( .A(n559), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT50), .B(n556), .Z(n557) );
  XNOR2_X1 U623 ( .A(G127GAT), .B(n557), .ZN(G1342GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n561) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(G134GAT), .B(n562), .Z(G1343GAT) );
  NAND2_X1 U628 ( .A1(n580), .A2(n563), .ZN(n572) );
  NOR2_X1 U629 ( .A1(n582), .A2(n572), .ZN(n564) );
  XOR2_X1 U630 ( .A(G141GAT), .B(n564), .Z(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT118), .B(n565), .ZN(G1344GAT) );
  NOR2_X1 U632 ( .A1(n572), .A2(n575), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n567) );
  XNOR2_X1 U634 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1345GAT) );
  NOR2_X1 U637 ( .A1(n570), .A2(n572), .ZN(n571) );
  XOR2_X1 U638 ( .A(G155GAT), .B(n571), .Z(G1346GAT) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G162GAT), .B(n574), .Z(G1347GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n593) );
  NOR2_X1 U646 ( .A1(n582), .A2(n593), .ZN(n586) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT60), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT126), .B(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT61), .Z(n588) );
  INV_X1 U652 ( .A(n593), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n590), .A2(n463), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U655 ( .A(G211GAT), .B(KEYINPUT127), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1354GAT) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(n595), .Z(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

