//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n190), .B2(G116), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n188), .A3(G119), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  XOR2_X1   g008(.A(KEYINPUT2), .B(G113), .Z(new_n195));
  AND2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G134), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n201), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(G131), .B1(new_n201), .B2(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n217), .A2(new_n226), .A3(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(G128), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n223), .B1(new_n228), .B2(new_n220), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT0), .A4(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n206), .A2(G137), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n207), .B2(new_n209), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n202), .B1(new_n204), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n213), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n199), .B1(new_n230), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n220), .ZN(new_n243));
  INV_X1    g057(.A(G128), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n221), .B1(G143), .B2(new_n216), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n226), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n246), .B2(new_n225), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n214), .B(new_n213), .C1(new_n247), .C2(new_n223), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n233), .A2(new_n234), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n237), .A2(new_n239), .A3(G131), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n212), .B1(new_n205), .B2(new_n211), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n252), .A3(new_n198), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n187), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n253), .A2(new_n187), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT28), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT28), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(KEYINPUT27), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n258), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n256), .A2(new_n270), .A3(new_n258), .A4(new_n266), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT30), .B1(new_n230), .B2(new_n241), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n248), .A2(new_n252), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n198), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n248), .A2(new_n252), .A3(new_n198), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n275), .A2(new_n276), .A3(new_n263), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n198), .B1(new_n248), .B2(new_n252), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT28), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n264), .B1(new_n279), .B2(new_n258), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n265), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n268), .A2(new_n269), .A3(new_n271), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G472), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n257), .B1(new_n242), .B2(new_n253), .ZN(new_n285));
  INV_X1    g099(.A(new_n258), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n264), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n253), .A2(new_n263), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT31), .B1(new_n275), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n272), .A2(new_n274), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n290), .B2(new_n199), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT67), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n275), .A2(new_n294), .A3(new_n288), .A4(KEYINPUT31), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n287), .B(new_n289), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n284), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n248), .A2(new_n252), .A3(new_n273), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n273), .B1(new_n248), .B2(new_n252), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n199), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n288), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n292), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n294), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n291), .A2(KEYINPUT67), .A3(new_n292), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n287), .A2(new_n289), .ZN(new_n308));
  AOI211_X1 g122(.A(KEYINPUT32), .B(new_n299), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n283), .B1(new_n298), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n311));
  XOR2_X1   g125(.A(KEYINPUT71), .B(G217), .Z(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G234), .B2(new_n269), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT73), .B(G125), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT16), .A2(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(G125), .A2(G140), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n314), .B2(G140), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  OAI211_X1 g133(.A(G146), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(G125), .A2(G140), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n216), .B1(new_n321), .B2(new_n317), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n323), .B1(new_n190), .B2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n190), .A2(G128), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(KEYINPUT23), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(new_n244), .B2(G119), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT72), .B1(new_n244), .B2(G119), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G110), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n244), .A2(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT24), .B(G110), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n332), .B1(new_n331), .B2(new_n336), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n320), .B(new_n322), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(KEYINPUT73), .A2(G125), .ZN(new_n340));
  NOR2_X1   g154(.A1(KEYINPUT73), .A2(G125), .ZN(new_n341));
  OAI21_X1  g155(.A(G140), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n317), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n319), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n316), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n216), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n320), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n334), .A2(new_n335), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n326), .A2(new_n329), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n348), .B1(new_n349), .B2(G110), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT75), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n339), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n339), .B2(new_n351), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT25), .B1(new_n359), .B2(new_n269), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NOR4_X1   g175(.A1(new_n357), .A2(new_n358), .A3(new_n361), .A4(G902), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n313), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n313), .A2(G902), .ZN(new_n364));
  XOR2_X1   g178(.A(new_n364), .B(KEYINPUT77), .Z(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT76), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n287), .A2(new_n289), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n305), .B2(new_n306), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT32), .B1(new_n374), .B2(new_n299), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n299), .B1(new_n307), .B2(new_n308), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n284), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT70), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n283), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n311), .A2(new_n372), .A3(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  OAI21_X1  g196(.A(G221), .B1(new_n382), .B2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n269), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G107), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(KEYINPUT3), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G104), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n395), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  AND2_X1   g216(.A1(KEYINPUT82), .A2(G101), .ZN(new_n403));
  NOR2_X1   g217(.A1(KEYINPUT82), .A2(G101), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n388), .A2(new_n390), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n402), .A2(new_n405), .A3(new_n393), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n398), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n402), .A3(KEYINPUT83), .A4(new_n405), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n400), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(G101), .C1(new_n392), .C2(new_n398), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n249), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT84), .B1(new_n389), .B2(G107), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n396), .A3(G104), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n419), .A3(new_n393), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n420), .A2(KEYINPUT85), .A3(G101), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT85), .B1(new_n420), .B2(G101), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n228), .A2(new_n220), .ZN(new_n425));
  INV_X1    g239(.A(new_n223), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT10), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n412), .A2(new_n415), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n220), .B1(new_n245), .B2(new_n244), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(new_n423), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n416), .A2(KEYINPUT86), .A3(new_n423), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT10), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n250), .A2(new_n251), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n427), .B1(new_n416), .B2(new_n423), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n439), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT12), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n434), .B2(new_n435), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT12), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(new_n439), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n440), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n352), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT80), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G140), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n437), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n434), .B2(new_n435), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n444), .B1(new_n458), .B2(new_n429), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n438), .B2(new_n439), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n449), .A2(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n386), .B1(new_n461), .B2(G469), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n443), .A2(KEYINPUT12), .A3(new_n444), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n447), .B1(new_n446), .B2(new_n439), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n460), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n436), .A2(new_n437), .ZN(new_n467));
  INV_X1    g281(.A(new_n429), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n439), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n458), .A2(new_n444), .A3(new_n429), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n456), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n385), .A3(new_n269), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n384), .B1(new_n462), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G214), .B1(G237), .B2(G902), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT88), .Z(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G122), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g295(.A(G113), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT5), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n189), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n481), .A2(new_n484), .B1(new_n194), .B2(new_n195), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n416), .A2(new_n423), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n414), .B1(new_n196), .B2(new_n197), .ZN(new_n487));
  INV_X1    g301(.A(new_n400), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(new_n416), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n480), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n416), .A2(new_n423), .A3(new_n485), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n479), .C1(new_n412), .C2(new_n487), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(KEYINPUT6), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT6), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n494), .B(new_n480), .C1(new_n486), .C2(new_n489), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n233), .A2(new_n314), .A3(new_n234), .ZN(new_n496));
  INV_X1    g310(.A(new_n314), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n427), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G224), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(G953), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n498), .B(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n493), .A2(new_n495), .A3(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n479), .B(KEYINPUT8), .Z(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n424), .B2(new_n485), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n481), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n194), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(new_n484), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n416), .B(new_n423), .C1(new_n508), .C2(new_n196), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT7), .B1(new_n499), .B2(G953), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n498), .A2(KEYINPUT90), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT90), .B1(new_n498), .B2(new_n511), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  OR2_X1    g329(.A1(new_n498), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n492), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n269), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n478), .B1(new_n502), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n493), .A2(new_n495), .A3(new_n501), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n492), .A2(new_n516), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n513), .B1(new_n509), .B2(new_n504), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n512), .A3(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n523), .A3(new_n269), .A4(new_n477), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n476), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n528));
  OAI21_X1  g342(.A(G131), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n259), .A2(G214), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n218), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n212), .A3(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT17), .B(G131), .C1(new_n527), .C2(new_n528), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n346), .A2(new_n534), .A3(new_n320), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(new_n212), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n527), .B2(new_n528), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT92), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n537), .B2(new_n212), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n531), .A2(new_n543), .A3(new_n526), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n342), .A2(G146), .A3(new_n343), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n322), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT91), .B(new_n538), .C1(new_n527), .C2(new_n528), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n541), .A2(new_n545), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  XOR2_X1   g363(.A(G113), .B(G122), .Z(new_n550));
  XOR2_X1   g364(.A(KEYINPUT93), .B(G104), .Z(new_n551));
  XOR2_X1   g365(.A(new_n550), .B(new_n551), .Z(new_n552));
  NAND3_X1  g366(.A1(new_n536), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n536), .A2(KEYINPUT94), .A3(new_n549), .A4(new_n552), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n536), .A2(new_n549), .ZN(new_n558));
  INV_X1    g372(.A(new_n552), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(KEYINPUT95), .A3(new_n269), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n555), .A2(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n563), .B1(new_n564), .B2(G902), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n565), .A3(G475), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n529), .A2(new_n532), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n318), .A2(KEYINPUT19), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n321), .A2(new_n317), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n568), .B1(KEYINPUT19), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n320), .B(new_n567), .C1(new_n570), .C2(G146), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n549), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n559), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n557), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n555), .A2(new_n556), .B1(new_n559), .B2(new_n572), .ZN(new_n578));
  INV_X1    g392(.A(new_n576), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT20), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n566), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G478), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(KEYINPUT15), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n312), .A2(G953), .A3(new_n382), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n244), .B2(G143), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n218), .A2(KEYINPUT13), .A3(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n244), .A2(G143), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G134), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n218), .A2(G128), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n591), .A3(new_n206), .ZN(new_n595));
  INV_X1    g409(.A(G122), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G116), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n188), .A2(G122), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n396), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n597), .A2(new_n598), .A3(new_n396), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n593), .B(new_n595), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n594), .A2(new_n591), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G134), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n595), .ZN(new_n604));
  XNOR2_X1  g418(.A(G116), .B(G122), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n396), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n188), .A2(KEYINPUT14), .A3(G122), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n597), .A2(new_n598), .ZN(new_n608));
  OAI211_X1 g422(.A(G107), .B(new_n607), .C1(new_n608), .C2(KEYINPUT14), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n601), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n601), .B2(new_n610), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n587), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n593), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n595), .B1(new_n600), .B2(new_n599), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n594), .A2(new_n591), .A3(new_n206), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n206), .B1(new_n594), .B2(new_n591), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n606), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n607), .A2(G107), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT14), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n605), .ZN(new_n622));
  OAI22_X1  g436(.A1(new_n615), .A2(new_n616), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT96), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n601), .A2(new_n610), .A3(new_n611), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n586), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n614), .A2(new_n626), .A3(new_n269), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n585), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n614), .A2(new_n626), .A3(KEYINPUT97), .A4(new_n269), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n629), .B1(new_n632), .B2(new_n585), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n352), .A2(G952), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(G234), .B2(G237), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n269), .B(new_n352), .C1(G234), .C2(G237), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT21), .B(G898), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n525), .A2(new_n583), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n474), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n381), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(new_n405), .Z(G3));
  NAND2_X1  g460(.A1(new_n460), .A2(new_n459), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n470), .B1(new_n463), .B2(new_n464), .ZN(new_n648));
  OAI211_X1 g462(.A(G469), .B(new_n647), .C1(new_n648), .C2(new_n455), .ZN(new_n649));
  INV_X1    g463(.A(new_n386), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI211_X1 g465(.A(G469), .B(G902), .C1(new_n466), .C2(new_n471), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n383), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n654));
  INV_X1    g468(.A(G472), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT98), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n371), .A2(new_n376), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(G472), .C1(new_n374), .C2(G902), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n475), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n661), .B1(new_n519), .B2(new_n524), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n614), .A2(new_n626), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(G478), .A3(new_n269), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n627), .A2(new_n584), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n566), .A2(new_n581), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n639), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n662), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n653), .A2(new_n660), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT34), .B(G104), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G6));
  AND3_X1   g487(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT99), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT99), .B1(new_n577), .B2(new_n580), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(G475), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n557), .B2(new_n560), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n677), .B1(new_n678), .B2(KEYINPUT95), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n632), .A2(new_n585), .ZN(new_n680));
  INV_X1    g494(.A(new_n629), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n679), .A2(new_n565), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n662), .A2(new_n676), .A3(new_n669), .A4(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n653), .A2(new_n660), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n396), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT100), .B(KEYINPUT35), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G9));
  INV_X1    g501(.A(new_n376), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n339), .A2(new_n351), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT36), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n356), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n689), .B(new_n691), .Z(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n366), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n363), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n656), .A2(new_n659), .A3(new_n688), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n474), .A3(new_n642), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  NAND3_X1  g513(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT99), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n581), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n636), .B1(new_n637), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n682), .A2(new_n700), .A3(new_n702), .A4(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n707));
  AOI21_X1  g521(.A(G902), .B1(new_n707), .B2(new_n521), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n477), .B1(new_n708), .B2(new_n520), .ZN(new_n709));
  INV_X1    g523(.A(new_n524), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n475), .B(new_n694), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n311), .A2(new_n474), .A3(new_n380), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  XOR2_X1   g528(.A(new_n704), .B(KEYINPUT39), .Z(new_n715));
  NAND2_X1  g529(.A1(new_n474), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(KEYINPUT40), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n302), .A2(new_n253), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n263), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT68), .B1(new_n276), .B2(new_n278), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n253), .A2(new_n187), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n720), .B(new_n269), .C1(new_n263), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G472), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n309), .B2(new_n298), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n519), .A2(new_n524), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT38), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n363), .A2(new_n693), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n633), .B1(new_n566), .B2(new_n581), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n475), .A2(new_n728), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n717), .A2(new_n718), .A3(new_n726), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G143), .ZN(G45));
  NAND2_X1  g547(.A1(new_n666), .A2(new_n667), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n582), .A2(new_n734), .A3(new_n705), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n311), .A2(new_n380), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n474), .A2(new_n662), .A3(new_n694), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT101), .B(G146), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G48));
  NAND2_X1  g555(.A1(new_n440), .A2(new_n459), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n456), .A2(new_n742), .B1(new_n465), .B2(new_n460), .ZN(new_n743));
  OAI21_X1  g557(.A(G469), .B1(new_n743), .B2(G902), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n383), .A3(new_n473), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n670), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n372), .A3(new_n311), .A4(new_n380), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT41), .B(G113), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT102), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n747), .B(new_n749), .ZN(G15));
  NOR2_X1   g564(.A1(new_n745), .A2(new_n683), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n372), .A3(new_n311), .A4(new_n380), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NAND2_X1  g567(.A1(new_n583), .A2(new_n640), .ZN(new_n754));
  INV_X1    g568(.A(new_n662), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n745), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n311), .A3(new_n380), .A4(new_n694), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  INV_X1    g572(.A(new_n745), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n257), .B1(new_n721), .B2(new_n722), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT103), .B1(new_n760), .B2(new_n286), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT103), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n256), .A2(new_n762), .A3(new_n258), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n264), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n289), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n305), .B2(new_n306), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n299), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n655), .B1(new_n296), .B2(new_n269), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n371), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n730), .A2(new_n727), .A3(new_n475), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n759), .A2(new_n669), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  AND4_X1   g586(.A1(new_n383), .A2(new_n744), .A3(new_n473), .A4(new_n662), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n735), .A2(new_n767), .A3(new_n768), .A4(new_n729), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  NOR2_X1   g590(.A1(new_n310), .A2(KEYINPUT70), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n379), .B1(new_n378), .B2(new_n283), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n473), .A2(new_n650), .A3(new_n649), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n727), .A2(new_n661), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n372), .A2(new_n780), .A3(new_n383), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n782), .A3(new_n783), .A4(new_n736), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n474), .A2(new_n372), .A3(new_n781), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT104), .B1(new_n737), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n371), .B1(new_n378), .B2(new_n283), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n735), .A2(new_n787), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n474), .A3(new_n781), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  XOR2_X1   g607(.A(new_n706), .B(KEYINPUT105), .Z(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n779), .A3(new_n782), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  NOR2_X1   g610(.A1(new_n461), .A2(KEYINPUT45), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n385), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n461), .A2(KEYINPUT45), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n650), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n473), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n801), .A2(new_n802), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n383), .B(new_n715), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT106), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n583), .A2(new_n734), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT43), .Z(new_n809));
  NAND3_X1  g623(.A1(new_n656), .A2(new_n688), .A3(new_n659), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n694), .A3(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n781), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  OAI21_X1  g632(.A(new_n383), .B1(new_n804), .B2(new_n805), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n736), .A2(new_n371), .A3(new_n781), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n779), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  AND2_X1   g641(.A1(new_n744), .A2(new_n473), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT107), .Z(new_n831));
  AOI22_X1  g645(.A1(new_n375), .A2(new_n377), .B1(G472), .B2(new_n724), .ZN(new_n832));
  OR3_X1    g646(.A1(new_n371), .A2(new_n384), .A3(new_n476), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n728), .A2(new_n808), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n828), .A2(new_n829), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n809), .A2(new_n636), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n745), .A2(new_n727), .A3(new_n661), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n789), .ZN(new_n840));
  XOR2_X1   g654(.A(new_n840), .B(KEYINPUT48), .Z(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n773), .A3(new_n769), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n635), .B(KEYINPUT117), .Z(new_n843));
  INV_X1    g657(.A(new_n668), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n838), .A2(new_n372), .A3(new_n636), .A4(new_n832), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n845), .A2(new_n582), .A3(new_n734), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n767), .A2(new_n768), .A3(new_n729), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n839), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n728), .A2(new_n475), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n837), .A2(new_n759), .A3(new_n769), .A4(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n850), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n828), .A2(new_n384), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n821), .A2(new_n822), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n837), .A2(new_n769), .A3(new_n781), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n847), .B1(new_n860), .B2(KEYINPUT51), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n860), .A2(KEYINPUT51), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n633), .A2(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(KEYINPUT108), .B(new_n629), .C1(new_n632), .C2(new_n585), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n566), .A2(new_n705), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n867), .A2(new_n674), .A3(new_n675), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n311), .A2(new_n869), .A3(new_n380), .A4(new_n694), .ZN(new_n870));
  INV_X1    g684(.A(new_n774), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n474), .A3(new_n781), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n795), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n582), .A2(new_n865), .A3(new_n866), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n525), .A2(new_n669), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n474), .A2(new_n876), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT109), .B1(new_n879), .B2(new_n697), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n525), .A2(new_n668), .A3(new_n669), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n474), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n311), .A2(new_n372), .A3(new_n380), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(new_n643), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n879), .A2(new_n697), .A3(KEYINPUT109), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT110), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n474), .A2(new_n876), .A3(new_n881), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n381), .B2(new_n644), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT109), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n867), .A2(new_n525), .A3(new_n583), .A4(new_n669), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n653), .A2(new_n891), .A3(new_n660), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n653), .A2(new_n695), .A3(new_n641), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND4_X1   g708(.A1(KEYINPUT110), .A2(new_n889), .A3(new_n886), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n875), .B1(new_n887), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT114), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n757), .A2(new_n747), .A3(new_n752), .A4(new_n771), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT115), .B(new_n898), .C1(new_n788), .C2(new_n791), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  INV_X1    g714(.A(new_n898), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n900), .B1(new_n792), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n713), .A2(new_n775), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT111), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n713), .A2(new_n775), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n739), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n770), .A2(new_n726), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT112), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n694), .A2(new_n704), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n383), .B(new_n911), .C1(new_n651), .C2(new_n652), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n780), .A2(KEYINPUT112), .A3(new_n383), .A4(new_n911), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT113), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n910), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n770), .A2(new_n726), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT113), .A2(new_n916), .A3(new_n914), .A4(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT52), .B1(new_n908), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n917), .A3(new_n914), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT113), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n913), .A2(KEYINPUT113), .A3(new_n914), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n713), .B(new_n775), .C1(new_n737), .C2(new_n738), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT52), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n920), .A2(KEYINPUT53), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n894), .A2(new_n645), .A3(new_n886), .A4(new_n882), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT110), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n889), .A2(KEYINPUT110), .A3(new_n894), .A4(new_n886), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT114), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n875), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n897), .A2(new_n903), .A3(new_n930), .A4(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n925), .A2(new_n928), .A3(new_n927), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n928), .B1(new_n925), .B2(new_n927), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n874), .B1(new_n933), .B2(new_n934), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n898), .B1(new_n788), .B2(new_n791), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT53), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n938), .A2(new_n939), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(KEYINPUT53), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n920), .A2(new_n929), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n946), .A3(new_n944), .A4(new_n943), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n953), .A3(KEYINPUT54), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n938), .A2(KEYINPUT116), .A3(new_n939), .A4(new_n947), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n863), .A2(new_n950), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n836), .B1(new_n958), .B2(new_n959), .ZN(G75));
  NOR2_X1   g774(.A1(new_n352), .A2(G952), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n936), .B1(new_n935), .B2(new_n875), .ZN(new_n963));
  AOI211_X1 g777(.A(KEYINPUT114), .B(new_n874), .C1(new_n933), .C2(new_n934), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n920), .A2(KEYINPUT53), .A3(new_n929), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n899), .A3(new_n902), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n965), .A2(new_n967), .B1(new_n946), .B2(new_n945), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n269), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT56), .B1(new_n969), .B2(G210), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n493), .A2(new_n495), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(new_n501), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT55), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n962), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(KEYINPUT119), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT120), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT120), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n970), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n977), .B2(new_n979), .ZN(G51));
  NAND2_X1  g794(.A1(new_n938), .A2(new_n947), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT54), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(KEYINPUT122), .A3(new_n948), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT122), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n984), .A3(KEYINPUT54), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n386), .B(KEYINPUT121), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT57), .Z(new_n987));
  NAND3_X1  g801(.A1(new_n983), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n472), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n969), .A2(new_n799), .A3(new_n798), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n961), .B1(new_n989), .B2(new_n990), .ZN(G54));
  AND3_X1   g805(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n962), .B1(new_n992), .B2(new_n574), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n574), .B2(new_n992), .ZN(G60));
  NAND2_X1  g808(.A1(G478), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT59), .Z(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT116), .B1(new_n968), .B2(new_n939), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n955), .A2(new_n954), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT123), .ZN(new_n1001));
  INV_X1    g815(.A(new_n665), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n996), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n983), .A2(new_n985), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n962), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1003), .A2(new_n1004), .A3(new_n1007), .ZN(G63));
  NAND2_X1  g822(.A1(G217), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT124), .Z(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT60), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n968), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n692), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n368), .A2(new_n369), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1013), .B(new_n962), .C1(new_n1015), .C2(new_n1012), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT61), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G66));
  OAI21_X1  g832(.A(G953), .B1(new_n638), .B2(new_n499), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT125), .Z(new_n1020));
  NAND2_X1  g834(.A1(new_n935), .A2(new_n901), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1020), .B1(new_n1022), .B2(G953), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n971), .B1(G898), .B2(new_n352), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(G69));
  XOR2_X1   g839(.A(new_n290), .B(new_n570), .Z(new_n1026));
  NAND2_X1  g840(.A1(G900), .A2(G953), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n807), .A2(new_n770), .A3(new_n789), .ZN(new_n1028));
  INV_X1    g842(.A(new_n817), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(new_n908), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1031), .A2(new_n795), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1030), .A2(new_n792), .A3(new_n826), .A4(new_n1032), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n1026), .B(new_n1027), .C1(new_n1033), .C2(G953), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n781), .B1(new_n877), .B2(new_n668), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n883), .A2(new_n716), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1036), .B1(new_n823), .B2(new_n825), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1031), .A2(new_n732), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  OR2_X1    g853(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1037), .A2(new_n817), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n1041), .A2(new_n352), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1034), .B1(new_n1042), .B2(new_n1026), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n352), .B1(G227), .B2(G900), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1044), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1034), .B(new_n1046), .C1(new_n1042), .C2(new_n1026), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1045), .A2(new_n1047), .ZN(G72));
  XNOR2_X1  g862(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1049));
  NAND2_X1  g863(.A1(G472), .A2(G902), .ZN(new_n1050));
  XNOR2_X1  g864(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1051), .B1(new_n1033), .B2(new_n1021), .ZN(new_n1052));
  XNOR2_X1  g866(.A(new_n277), .B(KEYINPUT127), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n961), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(new_n277), .ZN(new_n1055));
  AND3_X1   g869(.A1(new_n1055), .A2(new_n720), .A3(new_n1051), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n951), .A2(new_n953), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g871(.A(new_n1051), .B1(new_n1041), .B2(new_n1021), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1058), .A2(new_n263), .A3(new_n719), .ZN(new_n1059));
  AND3_X1   g873(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(G57));
endmodule


