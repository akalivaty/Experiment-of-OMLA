//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1329, new_n1330, new_n1331, new_n1332, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT68), .ZN(new_n238));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT69), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G226), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n247), .A2(new_n250), .A3(new_n252), .A4(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT13), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n259), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(G238), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n261), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n259), .B1(new_n255), .B2(new_n256), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n266), .A2(new_n269), .ZN(new_n273));
  OAI21_X1  g0073(.A(KEYINPUT13), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(G179), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT79), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n271), .A2(new_n274), .A3(KEYINPUT79), .A4(G179), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n262), .B1(new_n261), .B2(new_n270), .ZN(new_n280));
  NOR3_X1   g0080(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT13), .ZN(new_n281));
  OAI21_X1  g0081(.A(G169), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT14), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n284), .B(G169), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT80), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n209), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n209), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G68), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n210), .A2(G33), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(new_n214), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT11), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT11), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT78), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(KEYINPUT78), .A3(new_n303), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G68), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT12), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  INV_X1    g0111(.A(new_n308), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n289), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n308), .A2(KEYINPUT76), .A3(new_n209), .A4(new_n288), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n267), .A2(G20), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n310), .B1(new_n317), .B2(G68), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n286), .A2(new_n287), .B1(new_n306), .B2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n279), .A2(KEYINPUT80), .A3(new_n283), .A4(new_n285), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT75), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT3), .B(G33), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT71), .B1(new_n324), .B2(G1698), .ZN(new_n325));
  AND4_X1   g0125(.A1(KEYINPUT71), .A2(new_n247), .A3(new_n252), .A4(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(G238), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(G232), .A3(new_n249), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n247), .A2(new_n252), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G107), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n259), .B1(new_n327), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n266), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n260), .A2(new_n265), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(G244), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n323), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G238), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n247), .A2(new_n252), .A3(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n324), .A2(KEYINPUT71), .A3(G1698), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n328), .A2(new_n330), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n260), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT75), .A3(new_n335), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(G200), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n317), .A2(G77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT8), .B(G58), .ZN(new_n349));
  INV_X1    g0149(.A(new_n294), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n350), .B1(new_n210), .B2(new_n214), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n297), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n289), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(G77), .B2(new_n308), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT77), .B1(new_n347), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n346), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT75), .B1(new_n345), .B2(new_n335), .ZN(new_n360));
  OAI21_X1  g0160(.A(G190), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n356), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n358), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n359), .B2(new_n360), .ZN(new_n365));
  INV_X1    g0165(.A(new_n356), .ZN(new_n366));
  INV_X1    g0166(.A(G169), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n337), .A2(new_n367), .A3(new_n346), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n319), .A2(new_n306), .ZN(new_n370));
  OAI21_X1  g0170(.A(G200), .B1(new_n280), .B2(new_n281), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n271), .A2(G190), .A3(new_n274), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n322), .A2(new_n363), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT70), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n324), .A2(new_n376), .A3(G222), .A4(new_n249), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n324), .A2(G222), .A3(new_n249), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT70), .B1(new_n329), .B2(G77), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G223), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n341), .B2(new_n342), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n260), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n333), .B1(G226), .B2(new_n334), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n367), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(G179), .B2(new_n385), .ZN(new_n387));
  INV_X1    g0187(.A(new_n293), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G50), .A2(G58), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n210), .B1(new_n389), .B2(new_n295), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT8), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G58), .ZN(new_n392));
  INV_X1    g0192(.A(G58), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT8), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT73), .ZN(new_n395));
  OR3_X1    g0195(.A1(new_n393), .A2(KEYINPUT73), .A3(KEYINPUT8), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G150), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n397), .A2(new_n297), .B1(new_n398), .B2(new_n350), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT74), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n390), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI221_X1 g0201(.A(KEYINPUT74), .B1(new_n398), .B2(new_n350), .C1(new_n397), .C2(new_n297), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n388), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n291), .A2(new_n308), .A3(new_n292), .A4(new_n316), .ZN(new_n404));
  INV_X1    g0204(.A(G50), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G50), .B2(new_n308), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n387), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT9), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT9), .B1(new_n403), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT10), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n385), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(G200), .B2(new_n385), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n410), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n375), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT85), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n259), .A2(G232), .A3(new_n268), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n266), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT83), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n381), .A2(new_n249), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n248), .A2(G1698), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n247), .A2(new_n427), .A3(new_n252), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(G33), .A2(G87), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n260), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT83), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n266), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n426), .A2(new_n432), .A3(new_n416), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT84), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n259), .B1(new_n429), .B2(new_n430), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n425), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n435), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n312), .B1(new_n395), .B2(new_n396), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n395), .A2(new_n396), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT82), .B(new_n443), .C1(new_n444), .C2(new_n404), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT82), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n404), .A2(new_n444), .ZN(new_n447));
  INV_X1    g0247(.A(new_n443), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(G58), .B(G68), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(G20), .B1(G159), .B2(new_n294), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n246), .A2(G33), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n210), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT7), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(G20), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n455), .A2(new_n456), .B1(new_n329), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(KEYINPUT16), .B(new_n452), .C1(new_n458), .C2(new_n295), .ZN(new_n459));
  INV_X1    g0259(.A(new_n452), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT81), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n246), .A2(KEYINPUT81), .A3(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n252), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n457), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n456), .B1(new_n324), .B2(G20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n460), .B1(new_n467), .B2(G68), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n459), .B(new_n289), .C1(new_n468), .C2(KEYINPUT16), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n450), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n423), .B1(new_n442), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n450), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n435), .A2(new_n439), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT84), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(new_n476), .A3(KEYINPUT85), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT17), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n426), .A2(new_n434), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n438), .A2(G179), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n438), .A2(new_n425), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n367), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT18), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n484), .B(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT17), .B1(new_n472), .B2(new_n476), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n479), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n422), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n312), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n251), .A2(G1), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n388), .A2(new_n495), .A3(new_n308), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n493), .B1(new_n496), .B2(new_n492), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n456), .A2(new_n455), .B1(new_n464), .B2(new_n457), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n216), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n467), .A2(KEYINPUT87), .A3(G107), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n350), .A2(new_n214), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT86), .A2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT86), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n216), .A2(KEYINPUT6), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n492), .A2(new_n216), .ZN(new_n508));
  NOR2_X1   g0308(.A1(G97), .A2(G107), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n506), .A2(new_n507), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n502), .B1(new_n511), .B2(G20), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n500), .A2(new_n501), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n497), .B1(new_n513), .B2(new_n289), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n247), .A2(new_n252), .A3(G244), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(KEYINPUT4), .A2(G244), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n247), .A2(new_n252), .A3(new_n518), .A4(new_n249), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G283), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n247), .A2(new_n252), .A3(G250), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n249), .B1(new_n522), .B2(KEYINPUT4), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n260), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(KEYINPUT5), .B(G41), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n264), .A2(G1), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(G257), .A3(new_n259), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n267), .A2(G45), .ZN(new_n529));
  OR2_X1    g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G274), .ZN(new_n533));
  INV_X1    g0333(.A(new_n209), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(new_n258), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n524), .A2(new_n364), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n528), .A2(new_n536), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G1698), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n519), .A2(new_n520), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n517), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n539), .B1(new_n543), .B2(new_n260), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n538), .B1(new_n544), .B2(G169), .ZN(new_n545));
  OR2_X1    g0345(.A1(new_n514), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT88), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n547), .A3(G190), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n524), .A2(new_n537), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n416), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT88), .B1(new_n549), .B2(G200), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n514), .B(new_n548), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n247), .A2(new_n252), .A3(G244), .A4(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n247), .A2(new_n252), .A3(G238), .A4(new_n249), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G116), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n260), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n259), .A2(G274), .A3(new_n526), .ZN(new_n558));
  AND2_X1   g0358(.A1(G33), .A2(G41), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n529), .B(G250), .C1(new_n559), .C2(new_n209), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  NOR2_X1   g0364(.A1(G87), .A2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n503), .A2(new_n504), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT19), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n210), .B1(new_n256), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n324), .A2(new_n210), .A3(G68), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n297), .B1(new_n503), .B2(new_n504), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(KEYINPUT19), .C2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n289), .B1(new_n312), .B2(new_n352), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n293), .A2(new_n494), .A3(new_n312), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G87), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n561), .B1(new_n556), .B2(new_n260), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G190), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n564), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n576), .A2(G179), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n576), .A2(new_n367), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT89), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(G179), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT89), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n367), .C2(new_n576), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n572), .A2(new_n289), .ZN(new_n585));
  INV_X1    g0385(.A(new_n352), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n388), .A2(new_n495), .A3(new_n308), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n352), .A2(new_n312), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n573), .A2(KEYINPUT90), .A3(new_n587), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n581), .A2(new_n584), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n546), .A2(new_n552), .A3(new_n578), .A4(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n288), .A2(new_n209), .B1(G20), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(G33), .B1(new_n503), .B2(new_n504), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n520), .A2(new_n210), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(KEYINPUT20), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n312), .A2(new_n595), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n495), .A2(G116), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT91), .B1(new_n315), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT91), .ZN(new_n608));
  AOI211_X1 g0408(.A(new_n608), .B(new_n605), .C1(new_n313), .C2(new_n314), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n525), .A2(new_n526), .B1(new_n534), .B2(new_n258), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(G270), .B1(new_n532), .B2(new_n535), .ZN(new_n612));
  OAI21_X1  g0412(.A(G303), .B1(new_n453), .B2(new_n454), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n247), .A2(new_n252), .A3(G264), .A4(G1698), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n247), .A2(new_n252), .A3(G257), .A4(new_n249), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n260), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n367), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(KEYINPUT21), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n612), .A2(new_n617), .A3(G179), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT21), .B1(new_n610), .B2(new_n618), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT94), .ZN(new_n625));
  INV_X1    g0425(.A(new_n289), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n247), .A2(new_n252), .A3(new_n210), .A4(G87), .ZN(new_n627));
  NAND2_X1  g0427(.A1(KEYINPUT92), .A2(KEYINPUT22), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n324), .A2(new_n210), .A3(G87), .A4(new_n628), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n555), .A2(G20), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n210), .A2(G107), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT23), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT23), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n210), .B2(G107), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n633), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT24), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT24), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n632), .A2(new_n641), .A3(new_n638), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n626), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G13), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(G1), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n634), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(KEYINPUT93), .A3(KEYINPUT25), .ZN(new_n647));
  OR2_X1    g0447(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n648));
  NAND2_X1  g0448(.A1(KEYINPUT93), .A2(KEYINPUT25), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n645), .A2(new_n634), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n651), .B1(new_n574), .B2(G107), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n625), .B1(new_n643), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n642), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n641), .B1(new_n632), .B2(new_n638), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n289), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(KEYINPUT94), .A3(new_n652), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n247), .A2(new_n252), .A3(G257), .A4(G1698), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n247), .A2(new_n252), .A3(G250), .A4(new_n249), .ZN(new_n660));
  NAND2_X1  g0460(.A1(G33), .A2(G294), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n259), .B1(new_n662), .B2(KEYINPUT95), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT95), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n659), .A2(new_n660), .A3(new_n664), .A4(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n532), .A2(new_n260), .A3(new_n217), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(G179), .A3(new_n536), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n536), .ZN(new_n670));
  AOI211_X1 g0470(.A(new_n670), .B(new_n667), .C1(new_n663), .C2(new_n665), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n671), .B2(new_n367), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n654), .A2(new_n658), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n666), .A2(new_n416), .A3(new_n536), .A4(new_n668), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n671), .B2(G200), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n643), .A2(new_n653), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n612), .A2(new_n617), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G200), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n416), .B2(new_n678), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n610), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n624), .A2(new_n673), .A3(new_n677), .A4(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n491), .A2(new_n594), .A3(new_n683), .ZN(G372));
  NOR3_X1   g0484(.A1(new_n375), .A2(new_n421), .A3(new_n489), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n589), .B1(new_n579), .B2(new_n580), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n576), .A2(G190), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n576), .A2(new_n437), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n573), .A2(new_n575), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n582), .B1(new_n367), .B2(new_n576), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n589), .ZN(new_n693));
  AND4_X1   g0493(.A1(new_n546), .A2(new_n552), .A3(new_n677), .A4(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n666), .A2(new_n536), .A3(new_n668), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G169), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n696), .A2(new_n669), .B1(new_n657), .B2(new_n652), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n624), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n687), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n686), .A2(new_n578), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n701), .A2(new_n514), .A3(new_n545), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT96), .B1(new_n702), .B2(KEYINPUT26), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n514), .A2(new_n545), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT26), .B1(new_n704), .B2(new_n693), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT96), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(new_n593), .A3(KEYINPUT26), .A4(new_n578), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n685), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n369), .ZN(new_n712));
  AOI22_X1  g0512(.A1(new_n321), .A2(new_n320), .B1(new_n374), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n479), .A2(new_n488), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n486), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n419), .ZN(new_n716));
  INV_X1    g0516(.A(new_n420), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n409), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n711), .A2(new_n719), .ZN(G369));
  AND3_X1   g0520(.A1(new_n654), .A2(new_n658), .A3(new_n672), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n645), .A2(new_n210), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n723), .A2(new_n724), .A3(G213), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G343), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n721), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n673), .A2(new_n677), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n654), .A2(new_n658), .A3(new_n727), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n623), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n621), .A3(new_n619), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n727), .A2(new_n610), .ZN(new_n736));
  OR3_X1    g0536(.A1(new_n735), .A2(new_n736), .A3(new_n681), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n698), .A2(new_n727), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n730), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n732), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n727), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n743), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n750), .ZN(G399));
  INV_X1    g0551(.A(new_n204), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G41), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n566), .A2(G116), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n754), .A2(G1), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n207), .B2(new_n754), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT26), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n704), .A2(new_n593), .A3(new_n759), .A4(new_n578), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n704), .A2(new_n693), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n687), .B1(new_n761), .B2(KEYINPUT26), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n721), .A2(new_n735), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n546), .A2(new_n552), .A3(new_n677), .A4(new_n693), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n760), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(KEYINPUT29), .A3(new_n747), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n727), .B1(new_n700), .B2(new_n709), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(KEYINPUT29), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n727), .A2(KEYINPUT31), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n576), .A2(G179), .A3(new_n612), .A4(new_n617), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n667), .B1(new_n663), .B2(new_n665), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n771), .A2(KEYINPUT30), .A3(new_n544), .A4(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(G179), .B1(new_n612), .B2(new_n617), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n695), .A2(new_n549), .A3(new_n563), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n544), .A2(new_n620), .A3(new_n772), .A4(new_n576), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT30), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n769), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n775), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n777), .B2(new_n778), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n777), .A2(new_n783), .A3(new_n778), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n747), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n781), .B1(new_n787), .B2(KEYINPUT31), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n683), .A2(new_n594), .A3(new_n727), .ZN(new_n789));
  OAI21_X1  g0589(.A(G330), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n768), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n758), .B1(new_n792), .B2(G1), .ZN(G364));
  NOR2_X1   g0593(.A1(new_n644), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n267), .B1(new_n794), .B2(G45), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n753), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n210), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(new_n416), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n329), .B1(new_n800), .B2(G107), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n210), .A2(new_n364), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT100), .Z(new_n803));
  NOR2_X1   g0603(.A1(new_n416), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G190), .A2(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n801), .B1(new_n805), .B2(new_n393), .C1(new_n214), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n798), .A2(new_n806), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G159), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT32), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n802), .A2(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n416), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(G87), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n815), .A2(new_n405), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n808), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n813), .A2(G190), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n210), .B1(new_n804), .B2(new_n364), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n821), .A2(new_n295), .B1(new_n492), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT101), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n324), .B1(new_n810), .B2(G329), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  INV_X1    g0626(.A(G322), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n816), .C1(new_n805), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n807), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G311), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n799), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n814), .A2(G326), .ZN(new_n833));
  INV_X1    g0633(.A(G294), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n822), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT33), .B(G317), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n832), .B(new_n835), .C1(new_n820), .C2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n819), .A2(new_n824), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n209), .B1(G20), .B2(new_n367), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n797), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(G13), .A2(G33), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(G20), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n839), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n329), .A2(new_n204), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n264), .B2(new_n208), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n240), .B2(new_n264), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n752), .A2(new_n329), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n849), .A2(G355), .B1(new_n595), .B2(new_n752), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n841), .B1(new_n845), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n844), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n852), .B1(new_n739), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n797), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n740), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n739), .A2(G330), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT102), .ZN(G396));
  NAND2_X1  g0659(.A1(new_n366), .A2(new_n727), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n362), .A2(new_n361), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n357), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n369), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n712), .A2(new_n747), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n767), .B(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n797), .B1(new_n867), .B2(new_n790), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n790), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n839), .A2(new_n842), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n855), .B1(new_n214), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n369), .A2(new_n727), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n862), .B2(new_n369), .ZN(new_n873));
  AOI22_X1  g0673(.A1(G137), .A2(new_n814), .B1(new_n820), .B2(G150), .ZN(new_n874));
  INV_X1    g0674(.A(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G159), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n874), .B1(new_n805), .B2(new_n875), .C1(new_n876), .C2(new_n807), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT34), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n324), .B1(new_n809), .B2(new_n881), .C1(new_n295), .C2(new_n799), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n822), .A2(new_n393), .B1(new_n816), .B2(new_n405), .ZN(new_n883));
  NOR4_X1   g0683(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n829), .A2(G116), .B1(G283), .B2(new_n820), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n885), .A2(new_n886), .B1(new_n826), .B2(new_n815), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n886), .B2(new_n885), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT104), .Z(new_n889));
  INV_X1    g0689(.A(G311), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n329), .B1(new_n809), .B2(new_n890), .C1(new_n822), .C2(new_n492), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n817), .A2(new_n799), .B1(new_n816), .B2(new_n216), .ZN(new_n892));
  INV_X1    g0692(.A(new_n805), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(G294), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n884), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n871), .B1(new_n843), .B2(new_n873), .C1(new_n895), .C2(new_n840), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n869), .A2(new_n896), .ZN(G384));
  NOR2_X1   g0697(.A1(new_n794), .A2(new_n267), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n470), .A2(new_n725), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n484), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n478), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n459), .A2(new_n293), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT16), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n452), .B1(new_n458), .B2(new_n295), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n450), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n908), .A2(new_n909), .B1(new_n483), .B2(new_n725), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n471), .A2(new_n477), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT108), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT37), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n912), .B1(new_n911), .B2(KEYINPUT37), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n725), .B1(new_n908), .B2(new_n909), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n489), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n915), .A2(KEYINPUT38), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT38), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n487), .B1(new_n478), .B2(KEYINPUT17), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n900), .B1(new_n921), .B2(new_n486), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n484), .B(new_n900), .C1(new_n470), .C2(new_n442), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n904), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n277), .A2(new_n278), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n283), .A2(new_n285), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n287), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(new_n321), .A3(new_n370), .A4(new_n727), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n320), .A2(KEYINPUT107), .A3(new_n321), .A4(new_n727), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n370), .A2(new_n373), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n320), .B2(new_n321), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n370), .A2(new_n727), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AND4_X1   g0739(.A1(new_n546), .A2(new_n552), .A3(new_n578), .A4(new_n593), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n735), .A2(new_n681), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(new_n941), .A3(new_n731), .A4(new_n747), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n787), .A2(KEYINPUT31), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n666), .A2(new_n668), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n944), .A2(new_n549), .A3(new_n770), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT99), .B1(new_n945), .B2(KEYINPUT30), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n776), .A2(new_n946), .A3(new_n786), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n727), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT31), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n943), .A3(new_n950), .ZN(new_n951));
  AND3_X1   g0751(.A1(new_n939), .A2(new_n873), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n899), .B1(new_n926), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n939), .A2(new_n899), .A3(new_n951), .A4(new_n873), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT108), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT37), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n903), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n916), .B1(new_n921), .B2(new_n486), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n920), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n954), .B1(new_n919), .B2(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n953), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n685), .A3(new_n951), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(G330), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n962), .B1(new_n685), .B2(new_n951), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n926), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n322), .A2(new_n727), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n960), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n486), .A2(new_n725), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n864), .B(KEYINPUT106), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n767), .B2(new_n873), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n932), .A2(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n960), .A2(new_n919), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n971), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n685), .B(new_n766), .C1(KEYINPUT29), .C2(new_n767), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n719), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n979), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n898), .B1(new_n966), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n982), .B2(new_n966), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n985), .A2(G116), .A3(new_n211), .A4(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT105), .B(KEYINPUT36), .Z(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(G77), .B1(new_n393), .B2(new_n295), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n990), .A2(new_n207), .B1(G50), .B2(new_n295), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n991), .A2(G1), .A3(new_n644), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n984), .A2(new_n989), .A3(new_n992), .ZN(G367));
  AOI21_X1  g0793(.A(new_n748), .B1(new_n744), .B2(new_n745), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n546), .B(new_n552), .C1(new_n514), .C2(new_n747), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n704), .A2(new_n727), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n998), .A2(KEYINPUT42), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n546), .B1(new_n995), .B2(new_n673), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n998), .A2(KEYINPUT42), .B1(new_n747), .B2(new_n1000), .ZN(new_n1001));
  OR3_X1    g0801(.A1(new_n747), .A2(new_n691), .A3(new_n686), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n693), .B1(new_n747), .B2(new_n691), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n999), .A2(new_n1001), .B1(KEYINPUT43), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1004), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT43), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n997), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n742), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n999), .A2(new_n1001), .A3(new_n1007), .A4(new_n1006), .ZN(new_n1012));
  AND3_X1   g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1011), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n753), .B(KEYINPUT41), .Z(new_n1016));
  OAI22_X1  g0816(.A1(new_n733), .A2(new_n748), .B1(new_n698), .B2(new_n727), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(KEYINPUT44), .A3(new_n1010), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(KEYINPUT44), .B1(new_n1017), .B2(new_n1010), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT45), .B1(new_n750), .B2(new_n997), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT45), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1017), .A2(new_n1022), .A3(new_n1010), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1019), .A2(new_n1020), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n741), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1020), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1018), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n750), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1022), .B1(new_n1017), .B2(new_n1010), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(new_n1030), .A3(new_n742), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n733), .A2(new_n748), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n740), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n994), .B2(KEYINPUT109), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n994), .A2(new_n1033), .A3(KEYINPUT109), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n994), .A2(new_n1033), .A3(KEYINPUT109), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1032), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n1034), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n791), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1025), .A2(new_n1031), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1016), .B1(new_n1042), .B2(new_n792), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n795), .B(KEYINPUT110), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1015), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n234), .A2(new_n846), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n845), .B1(new_n204), .B2(new_n352), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n797), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n816), .A2(new_n393), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n329), .B(new_n1050), .C1(G137), .C2(new_n810), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n805), .B2(new_n398), .C1(new_n405), .C2(new_n807), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n799), .A2(new_n214), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n822), .A2(new_n295), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n821), .A2(new_n876), .B1(new_n815), .B2(new_n875), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n329), .B1(new_n809), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n822), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(G107), .B2(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n805), .B2(new_n826), .C1(new_n831), .C2(new_n807), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n816), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT111), .B1(new_n1062), .B2(G116), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT46), .Z(new_n1064));
  AOI22_X1  g0864(.A1(new_n814), .A2(G311), .B1(new_n800), .B2(new_n505), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n834), .B2(new_n821), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1056), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1049), .B1(new_n1070), .B2(new_n839), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n853), .B2(new_n1004), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1046), .A2(new_n1072), .ZN(G387));
  NAND2_X1  g0873(.A1(new_n229), .A2(G45), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT113), .Z(new_n1075));
  NOR2_X1   g0875(.A1(new_n349), .A2(G50), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n755), .ZN(new_n1078));
  AOI211_X1 g0878(.A(G45), .B(new_n1078), .C1(G68), .C2(G77), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n846), .B(new_n1075), .C1(new_n1077), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n849), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1081), .A2(new_n755), .B1(G107), .B2(new_n204), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n845), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n807), .A2(new_n295), .B1(new_n397), .B2(new_n821), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n816), .A2(new_n214), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n822), .A2(new_n352), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(G97), .C2(new_n800), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n324), .B1(new_n809), .B2(new_n398), .C1(new_n815), .C2(new_n876), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n893), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n324), .B1(new_n810), .B2(G326), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n822), .A2(new_n831), .B1(new_n816), .B2(new_n834), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G311), .A2(new_n820), .B1(new_n814), .B2(G322), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n805), .B2(new_n1057), .C1(new_n826), .C2(new_n807), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT49), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1092), .B1(new_n595), .B2(new_n799), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n839), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1083), .A2(new_n1103), .A3(new_n797), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n733), .B2(new_n844), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1105), .B1(new_n1106), .B2(new_n1045), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1041), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n753), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1106), .A2(new_n792), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(G393));
  NOR2_X1   g0911(.A1(new_n1024), .A2(new_n741), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n742), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n753), .A3(new_n1042), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n244), .A2(new_n846), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n845), .B1(new_n204), .B2(new_n506), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n797), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n805), .A2(new_n876), .B1(new_n398), .B2(new_n815), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT51), .Z(new_n1120));
  NOR2_X1   g0920(.A1(new_n822), .A2(new_n214), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G50), .B2(new_n820), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n295), .B2(new_n816), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n807), .A2(new_n349), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n324), .B1(new_n809), .B2(new_n875), .C1(new_n817), .C2(new_n799), .ZN(new_n1125));
  OR4_X1    g0925(.A1(new_n1120), .A2(new_n1123), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n805), .A2(new_n890), .B1(new_n1057), .B2(new_n815), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT52), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n821), .A2(new_n826), .B1(new_n595), .B2(new_n822), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G283), .B2(new_n1062), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n329), .B1(new_n809), .B2(new_n827), .C1(new_n216), .C2(new_n799), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n829), .B2(G294), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n840), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1118), .B(new_n1134), .C1(new_n844), .C2(new_n1010), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1136), .B2(new_n1045), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1115), .A2(new_n1137), .ZN(G390));
  NAND4_X1  g0938(.A1(new_n939), .A2(G330), .A3(new_n951), .A4(new_n873), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n708), .B1(new_n705), .B2(new_n706), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n702), .A2(KEYINPUT96), .A3(KEYINPUT26), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n697), .A2(new_n622), .A3(new_n623), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n686), .B1(new_n764), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n873), .B(new_n747), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n872), .B(KEYINPUT106), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n969), .B1(new_n1148), .B2(new_n939), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n968), .B2(new_n970), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n765), .A2(new_n873), .A3(new_n747), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n969), .B1(new_n1152), .B2(new_n939), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n926), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1140), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n969), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n974), .B2(new_n975), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n960), .A2(KEYINPUT39), .A3(new_n919), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT39), .B1(new_n919), .B2(new_n925), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(G330), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n780), .B1(new_n948), .B2(new_n949), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n942), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1164), .A2(new_n939), .A3(new_n873), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT115), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n865), .B1(new_n938), .B2(new_n934), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT115), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1168), .A3(new_n1164), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1161), .A2(new_n1170), .A3(new_n1154), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1156), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1045), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n842), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n870), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n797), .B1(new_n444), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n815), .A2(new_n831), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1121), .B(new_n1177), .C1(G107), .C2(new_n820), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n799), .A2(new_n295), .B1(new_n809), .B2(new_n834), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n829), .B2(new_n505), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n595), .C2(new_n805), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n329), .B1(new_n816), .B2(new_n817), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT119), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n815), .A2(new_n1184), .B1(new_n876), .B2(new_n822), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G137), .B2(new_n820), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n799), .A2(new_n405), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n329), .B(new_n1187), .C1(G125), .C2(new_n810), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(KEYINPUT54), .B(G143), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1186), .B(new_n1188), .C1(new_n807), .C2(new_n1189), .ZN(new_n1190));
  OR3_X1    g0990(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n398), .ZN(new_n1191));
  OAI21_X1  g0991(.A(KEYINPUT53), .B1(new_n816), .B2(new_n398), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(new_n805), .C2(new_n881), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1181), .A2(new_n1183), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1176), .B1(new_n1194), .B2(new_n839), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1174), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1173), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT118), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT117), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n422), .A2(new_n951), .A3(G330), .A4(new_n490), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n719), .B(new_n1201), .C1(new_n768), .C2(new_n491), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT116), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT116), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n980), .A2(new_n1204), .A3(new_n719), .A4(new_n1201), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(G330), .B(new_n873), .C1(new_n788), .C2(new_n789), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n975), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n974), .B1(new_n1208), .B2(new_n1139), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n951), .A2(G330), .A3(new_n873), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1152), .B1(new_n975), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1170), .B2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1200), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n790), .A2(new_n975), .A3(KEYINPUT115), .A4(new_n865), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1168), .B1(new_n1167), .B2(new_n1164), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1211), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1209), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1218), .A2(KEYINPUT117), .A3(new_n1205), .A4(new_n1203), .ZN(new_n1219));
  AND2_X1   g1019(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1156), .A2(new_n1171), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n754), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1213), .A2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1172), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1199), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1221), .A2(new_n1213), .A3(new_n1219), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1224), .A2(new_n1226), .A3(new_n1199), .A4(new_n753), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1198), .B1(new_n1225), .B2(new_n1228), .ZN(G378));
  INV_X1    g1029(.A(new_n421), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n725), .B1(new_n403), .B2(new_n407), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1232), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n842), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n797), .B1(G50), .B2(new_n1175), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n815), .A2(new_n595), .B1(new_n799), .B2(new_n393), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1086), .B(new_n1243), .C1(G97), .C2(new_n820), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n263), .B(new_n329), .C1(new_n809), .C2(new_n831), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1054), .B(new_n1245), .C1(new_n893), .C2(G107), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1244), .B(new_n1246), .C1(new_n352), .C2(new_n807), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT120), .Z(new_n1248));
  INV_X1    g1048(.A(KEYINPUT58), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(G33), .A2(G41), .ZN(new_n1252));
  AOI211_X1 g1052(.A(G50), .B(new_n1252), .C1(new_n329), .C2(new_n263), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(G128), .A2(new_n893), .B1(new_n829), .B2(G137), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n814), .A2(G125), .B1(new_n1059), .B2(G150), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1189), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n820), .A2(G132), .B1(new_n1062), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1259));
  INV_X1    g1059(.A(G124), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1252), .B1(new_n809), .B2(new_n1260), .C1(new_n876), .C2(new_n799), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1258), .B2(KEYINPUT59), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1253), .B1(new_n1259), .B2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1250), .A2(new_n1251), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1242), .B1(new_n1264), .B2(new_n839), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1241), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(G330), .B1(new_n953), .B2(new_n961), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1240), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n979), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1239), .B(G330), .C1(new_n953), .C2(new_n961), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1266), .B1(new_n1273), .B2(new_n1044), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1224), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n979), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT57), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1206), .B1(new_n1223), .B2(new_n1172), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n753), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1275), .B1(new_n1282), .B2(new_n1285), .ZN(G375));
  NAND2_X1  g1086(.A1(new_n975), .A2(new_n842), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n814), .A2(G132), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(KEYINPUT123), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1059), .A2(G50), .B1(new_n1062), .B2(G159), .ZN(new_n1290));
  OAI211_X1 g1090(.A(new_n1289), .B(new_n1290), .C1(new_n821), .C2(new_n1189), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n893), .A2(G137), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n807), .A2(new_n398), .ZN(new_n1293));
  OAI221_X1 g1093(.A(new_n324), .B1(new_n809), .B2(new_n1184), .C1(new_n393), .C2(new_n799), .ZN(new_n1294));
  NOR4_X1   g1094(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .A4(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1087), .B1(G97), .B2(new_n1062), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n834), .B2(new_n815), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n324), .B(new_n1053), .C1(G303), .C2(new_n810), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n831), .B2(new_n805), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT122), .ZN(new_n1300));
  OAI22_X1  g1100(.A1(new_n807), .A2(new_n216), .B1(new_n595), .B2(new_n821), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1297), .B(new_n1299), .C1(new_n1300), .C2(new_n1301), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1301), .A2(new_n1300), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1295), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1304), .A2(new_n840), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n855), .B(new_n1305), .C1(new_n295), .C2(new_n870), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1218), .A2(new_n1045), .B1(new_n1287), .B2(new_n1306), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n1223), .A2(new_n1016), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1276), .A2(KEYINPUT121), .A3(new_n1218), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT121), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1307), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  XNOR2_X1  g1114(.A(new_n1314), .B(KEYINPUT124), .ZN(G381));
  AOI21_X1  g1115(.A(new_n1197), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(G390), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(G393), .A2(G396), .ZN(new_n1319));
  INV_X1    g1119(.A(G384), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  NOR4_X1   g1121(.A1(G381), .A2(G387), .A3(new_n1317), .A4(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT57), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n754), .B1(new_n1277), .B2(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1323), .B1(new_n1284), .B2(new_n1273), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1274), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1322), .A2(new_n1327), .ZN(G407));
  INV_X1    g1128(.A(G343), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(G213), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1327), .A2(new_n1316), .A3(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(G407), .A2(G213), .A3(new_n1332), .ZN(G409));
  AND2_X1   g1133(.A1(G393), .A2(G396), .ZN(new_n1334));
  OR2_X1    g1134(.A1(new_n1334), .A2(new_n1319), .ZN(new_n1335));
  AND3_X1   g1135(.A1(new_n1046), .A2(G390), .A3(new_n1072), .ZN(new_n1336));
  AOI21_X1  g1136(.A(G390), .B1(new_n1046), .B2(new_n1072), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(new_n1318), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1334), .A2(new_n1319), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1046), .A2(G390), .A3(new_n1072), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1338), .A2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(KEYINPUT126), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1284), .A2(new_n1273), .A3(new_n1016), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1316), .B1(new_n1345), .B2(new_n1274), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1226), .A2(new_n753), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1221), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1348));
  OAI21_X1  g1148(.A(KEYINPUT118), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1197), .B1(new_n1349), .B2(new_n1227), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1346), .B1(G375), .B2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1330), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1206), .A2(new_n1212), .A3(KEYINPUT60), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n753), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1213), .A2(new_n1219), .A3(KEYINPUT60), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1354), .B1(new_n1312), .B2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1357), .A2(G384), .A3(new_n1307), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1307), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1320), .B1(new_n1356), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1331), .A2(G2897), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1358), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1361), .B1(new_n1358), .B2(new_n1360), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT61), .B1(new_n1352), .B2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1358), .A2(new_n1360), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1351), .A2(new_n1367), .A3(new_n1330), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(KEYINPUT62), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1365), .A2(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1368), .A2(KEYINPUT62), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1344), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(G378), .A2(new_n1327), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1331), .B1(new_n1373), .B2(new_n1346), .ZN(new_n1374));
  AOI21_X1  g1174(.A(KEYINPUT63), .B1(new_n1374), .B2(new_n1367), .ZN(new_n1375));
  AND3_X1   g1175(.A1(new_n1358), .A2(KEYINPUT63), .A3(new_n1360), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1351), .A2(new_n1330), .A3(new_n1376), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1377), .A2(new_n1343), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1375), .A2(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(KEYINPUT125), .B1(new_n1379), .B2(new_n1365), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1338), .A2(new_n1342), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1381), .B1(new_n1374), .B2(new_n1376), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT63), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1368), .A2(new_n1383), .ZN(new_n1384));
  AND4_X1   g1184(.A1(KEYINPUT125), .A2(new_n1365), .A3(new_n1382), .A4(new_n1384), .ZN(new_n1385));
  OAI21_X1  g1185(.A(new_n1372), .B1(new_n1380), .B2(new_n1385), .ZN(G405));
  NAND2_X1  g1186(.A1(G375), .A2(new_n1316), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1373), .A2(new_n1387), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(KEYINPUT127), .ZN(new_n1389));
  INV_X1    g1189(.A(KEYINPUT127), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1373), .A2(new_n1387), .A3(new_n1390), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1389), .A2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1392), .A2(new_n1367), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1389), .A2(new_n1366), .A3(new_n1391), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1395), .A2(new_n1381), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(new_n1393), .A2(new_n1343), .A3(new_n1394), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(G402));
endmodule


