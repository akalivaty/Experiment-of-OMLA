//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(G475), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G214), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(G143), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n194), .B(new_n198), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n197), .B(KEYINPUT83), .C1(KEYINPUT18), .C2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(KEYINPUT18), .A3(G131), .ZN(new_n201));
  AND2_X1   g015(.A1(G125), .A2(G140), .ZN(new_n202));
  NOR2_X1   g016(.A1(G125), .A2(G140), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(G146), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT18), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n195), .B(new_n206), .C1(new_n207), .C2(new_n196), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n200), .A2(new_n201), .A3(new_n205), .A4(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n197), .A3(new_n212), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT16), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  INV_X1    g031(.A(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(G125), .A2(G140), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n216), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n217), .A2(KEYINPUT16), .A3(G140), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT16), .B1(new_n202), .B2(new_n203), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n199), .A2(KEYINPUT85), .A3(KEYINPUT17), .A4(G131), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n213), .A2(new_n214), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G113), .B(G122), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n209), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n204), .B(KEYINPUT19), .ZN(new_n235));
  OR3_X1    g049(.A1(new_n235), .A2(KEYINPUT84), .A3(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n211), .A2(new_n197), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT84), .B1(new_n235), .B2(G146), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n236), .A2(new_n226), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n233), .B1(new_n239), .B2(new_n209), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n190), .B(new_n191), .C1(new_n234), .C2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT20), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n233), .B1(new_n209), .B2(new_n230), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n191), .B1(new_n234), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT86), .B(new_n191), .C1(new_n234), .C2(new_n243), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G475), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT14), .ZN(new_n250));
  INV_X1    g064(.A(G122), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(G116), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n250), .A2(new_n252), .B1(new_n253), .B2(KEYINPUT87), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT87), .A4(G122), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n250), .B2(new_n252), .ZN(new_n257));
  OAI21_X1  g071(.A(G107), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT88), .ZN(new_n259));
  XNOR2_X1  g073(.A(G116), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(G107), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G128), .B(G143), .ZN(new_n263));
  INV_X1    g077(.A(G134), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G107), .C1(new_n254), .C2(new_n257), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n259), .A2(new_n262), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(KEYINPUT13), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n198), .A2(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n269), .B(G134), .C1(KEYINPUT13), .C2(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n260), .B(new_n261), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n263), .A2(new_n264), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G217), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n188), .A2(new_n276), .A3(G953), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n268), .A2(new_n274), .A3(new_n277), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n191), .ZN(new_n282));
  INV_X1    g096(.A(G478), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n282), .B(new_n284), .Z(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n249), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G110), .B(G140), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n193), .A2(G227), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n198), .B(G146), .C1(new_n293), .C2(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n215), .A3(G143), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n293), .A2(KEYINPUT1), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n215), .A2(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n198), .A2(G146), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n292), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  AND4_X1   g115(.A1(new_n292), .A2(new_n300), .A3(new_n295), .A4(new_n294), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT10), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT3), .B1(new_n232), .B2(G107), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n261), .A3(G104), .ZN(new_n306));
  INV_X1    g120(.A(G101), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n232), .A2(G107), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n304), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n261), .A2(G104), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n232), .A2(G107), .ZN(new_n311));
  OAI21_X1  g125(.A(G101), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT75), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n309), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(KEYINPUT76), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n309), .A2(new_n312), .A3(new_n315), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n315), .B1(new_n309), .B2(new_n312), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n303), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n298), .A2(new_n299), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT0), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(new_n293), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT0), .A2(G128), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n323), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n298), .B(new_n299), .C1(new_n324), .C2(new_n293), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n304), .A2(new_n306), .A3(new_n308), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT74), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n304), .A2(new_n306), .A3(new_n333), .A4(new_n308), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(G101), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n309), .A2(KEYINPUT4), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n332), .A2(KEYINPUT4), .A3(G101), .A4(new_n334), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT11), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n264), .B2(G137), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n264), .A2(G137), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .A3(G134), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT64), .A3(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT64), .A2(G131), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(new_n344), .A3(new_n347), .A4(new_n342), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n313), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n300), .A2(new_n295), .A3(new_n294), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT10), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR4_X1   g166(.A1(new_n322), .A2(new_n339), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n314), .B2(new_n316), .ZN(new_n354));
  INV_X1    g168(.A(new_n351), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(new_n313), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n349), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT12), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT12), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n359), .B(new_n349), .C1(new_n354), .C2(new_n356), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n291), .B1(new_n353), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n337), .A2(new_n338), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n352), .B1(new_n363), .B2(new_n329), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n351), .A2(KEYINPUT67), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n296), .A2(new_n292), .A3(new_n300), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n319), .A2(new_n320), .A3(new_n318), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT76), .B1(new_n314), .B2(new_n316), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n349), .ZN(new_n373));
  INV_X1    g187(.A(new_n349), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n364), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n375), .A3(new_n290), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n362), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G469), .B1(new_n377), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n374), .B1(new_n364), .B2(new_n371), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n291), .B1(new_n353), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n375), .A2(new_n358), .A3(new_n360), .A4(new_n290), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  AND4_X1   g198(.A1(new_n379), .A2(new_n383), .A3(new_n384), .A4(new_n191), .ZN(new_n385));
  AOI21_X1  g199(.A(G902), .B1(new_n381), .B2(new_n382), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n379), .B1(new_n386), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n378), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G234), .ZN(new_n389));
  OAI211_X1 g203(.A(G952), .B(new_n193), .C1(new_n389), .C2(new_n192), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT89), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT21), .B(G898), .Z(new_n392));
  OAI211_X1 g206(.A(G902), .B(G953), .C1(new_n389), .C2(new_n192), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AND4_X1   g208(.A1(new_n189), .A2(new_n287), .A3(new_n388), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n396));
  OAI21_X1  g210(.A(G210), .B1(G237), .B2(G902), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G113), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT2), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G113), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT66), .ZN(new_n408));
  NOR3_X1   g222(.A1(new_n255), .A2(KEYINPUT5), .A3(G119), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n404), .B2(KEYINPUT5), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n407), .A2(new_n408), .B1(G113), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n369), .B2(new_n370), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n408), .ZN(new_n415));
  XOR2_X1   g229(.A(G116), .B(G119), .Z(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n400), .A3(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n363), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(KEYINPUT78), .B(new_n411), .C1(new_n369), .C2(new_n370), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XOR2_X1   g235(.A(G110), .B(G122), .Z(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n422), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n414), .A2(new_n424), .A3(new_n419), .A4(new_n420), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n423), .A2(KEYINPUT6), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT6), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT79), .B1(new_n351), .B2(G125), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n296), .A2(new_n430), .A3(new_n217), .A4(new_n300), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n429), .B(new_n431), .C1(new_n217), .C2(new_n329), .ZN(new_n432));
  INV_X1    g246(.A(G224), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(G953), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n432), .B(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n404), .A2(KEYINPUT5), .ZN(new_n437));
  INV_X1    g251(.A(new_n409), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(G113), .A3(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n415), .B(new_n439), .C1(new_n319), .C2(new_n320), .ZN(new_n440));
  INV_X1    g254(.A(new_n408), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT66), .B1(new_n403), .B2(new_n404), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n350), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n422), .A2(KEYINPUT8), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT8), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n424), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n440), .A2(new_n444), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT80), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n314), .A2(new_n316), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n450), .A2(new_n411), .B1(new_n446), .B2(new_n424), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n451), .A2(new_n452), .A3(new_n445), .A4(new_n444), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(new_n433), .B2(G953), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n432), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n330), .A2(G125), .ZN(new_n457));
  INV_X1    g271(.A(new_n455), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n457), .A2(new_n429), .A3(new_n431), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n425), .B1(new_n462), .B2(KEYINPUT81), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n449), .B2(new_n453), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n191), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n398), .B1(new_n436), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n421), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n424), .B1(new_n464), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n462), .A2(KEYINPUT81), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n426), .A2(new_n428), .A3(new_n435), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n397), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n396), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  AOI211_X1 g292(.A(KEYINPUT82), .B(new_n478), .C1(new_n468), .C2(new_n474), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n395), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT90), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n395), .B(new_n482), .C1(new_n477), .C2(new_n479), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n226), .B1(G146), .B2(new_n204), .ZN(new_n484));
  INV_X1    g298(.A(G119), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT23), .B1(new_n485), .B2(G128), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n293), .A3(G119), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n486), .A2(new_n488), .B1(new_n485), .B2(G128), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT72), .B(G110), .Z(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(G128), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n293), .A2(G119), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT24), .B(G110), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n489), .A2(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n484), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n486), .A2(new_n488), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n491), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(G110), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n227), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT71), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n227), .A2(new_n503), .A3(new_n497), .A4(new_n500), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n496), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n507), .B(new_n496), .C1(new_n502), .C2(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n193), .A2(G221), .A3(G234), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT22), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(G137), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n506), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n505), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n513), .A2(new_n507), .A3(new_n511), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n191), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n276), .B1(G234), .B2(new_n191), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT25), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n518), .B(new_n191), .C1(new_n512), .C2(new_n514), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  OR2_X1    g334(.A1(new_n512), .A2(new_n514), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n517), .A2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n345), .A2(new_n196), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n343), .A2(G134), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n342), .A2(new_n527), .A3(G131), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n526), .A2(KEYINPUT65), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT65), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(new_n355), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n346), .A2(new_n348), .B1(new_n327), .B2(new_n328), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n525), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n366), .A2(new_n367), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n526), .A2(new_n528), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(new_n418), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n535), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n415), .A2(new_n417), .ZN(new_n540));
  INV_X1    g354(.A(new_n532), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(G101), .ZN(new_n544));
  INV_X1    g358(.A(G210), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n545), .A2(G237), .A3(G953), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n544), .B(new_n546), .Z(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT31), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n542), .A2(KEYINPUT28), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n536), .A2(new_n551), .A3(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n418), .B1(new_n531), .B2(new_n532), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n547), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT68), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n548), .B2(KEYINPUT31), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT65), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n535), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n526), .A2(KEYINPUT65), .A3(new_n528), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n351), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT30), .B1(new_n564), .B2(new_n541), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n366), .A2(new_n367), .B1(new_n526), .B2(new_n528), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n566), .A2(new_n525), .A3(new_n532), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n565), .A2(new_n567), .A3(new_n540), .ZN(new_n568));
  INV_X1    g382(.A(new_n542), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(KEYINPUT68), .A3(new_n571), .A4(new_n547), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n558), .B1(new_n560), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G472), .A2(G902), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT32), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n560), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n549), .A2(new_n557), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n574), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n551), .B1(new_n536), .B2(new_n540), .ZN(new_n583));
  NOR4_X1   g397(.A1(new_n566), .A2(new_n418), .A3(KEYINPUT28), .A4(new_n532), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n547), .B(new_n554), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT69), .ZN(new_n586));
  AOI21_X1  g400(.A(KEYINPUT29), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n556), .B1(new_n568), .B2(new_n569), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n553), .A2(KEYINPUT69), .A3(new_n547), .A4(new_n554), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT70), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT70), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(new_n592), .A3(new_n588), .A4(new_n589), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n418), .B1(new_n566), .B2(new_n532), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n553), .A2(KEYINPUT29), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n595), .B2(new_n547), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n591), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n524), .B1(new_n582), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n481), .A2(new_n483), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n573), .B2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n191), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(G472), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT92), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n579), .A2(new_n574), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n603), .A2(new_n608), .A3(new_n604), .A4(G472), .ZN(new_n609));
  AND4_X1   g423(.A1(new_n388), .A2(new_n606), .A3(new_n607), .A4(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n189), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n524), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT93), .ZN(new_n614));
  INV_X1    g428(.A(new_n249), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n277), .B1(new_n268), .B2(new_n274), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n280), .B2(new_n279), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n279), .B(new_n280), .C1(KEYINPUT94), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(G478), .B(new_n191), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT95), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n282), .A2(new_n283), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n281), .B(KEYINPUT33), .C1(new_n617), .C2(new_n616), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n621), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n627), .A2(new_n628), .A3(G478), .A4(new_n191), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT96), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n624), .A2(new_n632), .A3(new_n629), .A4(new_n625), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n615), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n472), .A2(new_n397), .A3(new_n473), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n397), .B1(new_n472), .B2(new_n473), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n394), .B(new_n476), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n614), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT97), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G6));
  AOI21_X1  g456(.A(new_n478), .B1(new_n468), .B2(new_n474), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n249), .A2(new_n285), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n394), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n645), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT98), .B1(new_n638), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n614), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT35), .B(G107), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NAND3_X1  g465(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT36), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n511), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n505), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n522), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n520), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n481), .A2(new_n483), .A3(new_n653), .A4(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT37), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(G12));
  OAI21_X1  g475(.A(new_n476), .B1(new_n636), .B2(new_n637), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n582), .B2(new_n598), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n391), .B1(G900), .B2(new_n393), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT99), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n647), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n388), .A2(new_n189), .ZN(new_n667));
  INV_X1    g481(.A(new_n658), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n663), .A2(KEYINPUT100), .A3(new_n666), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT101), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n293), .ZN(G30));
  XNOR2_X1  g490(.A(new_n665), .B(KEYINPUT39), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n388), .A2(new_n189), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n249), .A2(new_n286), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n679), .B2(KEYINPUT40), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n680), .A2(new_n476), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n547), .B1(new_n542), .B2(new_n594), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n570), .B2(new_n547), .ZN(new_n685));
  OAI21_X1  g499(.A(G472), .B1(new_n685), .B2(G902), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n582), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n475), .B(KEYINPUT38), .Z(new_n689));
  NOR4_X1   g503(.A1(new_n683), .A2(new_n658), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT102), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n198), .ZN(G45));
  AOI211_X1 g506(.A(new_n615), .B(new_n665), .C1(new_n631), .C2(new_n633), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n663), .A2(new_n693), .A3(new_n669), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OR2_X1    g509(.A1(new_n386), .A2(new_n384), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n189), .B(new_n696), .C1(new_n385), .C2(new_n387), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n386), .A2(new_n384), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n290), .B1(new_n373), .B2(new_n375), .ZN(new_n701));
  AND4_X1   g515(.A1(new_n375), .A2(new_n358), .A3(new_n360), .A4(new_n290), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n384), .B(new_n191), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT77), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n386), .A2(new_n379), .A3(new_n384), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(KEYINPUT103), .A3(new_n189), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n394), .ZN(new_n709));
  AOI211_X1 g523(.A(new_n709), .B(new_n478), .C1(new_n468), .C2(new_n474), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n599), .A2(new_n708), .A3(new_n634), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  AOI21_X1  g527(.A(new_n580), .B1(new_n579), .B2(new_n574), .ZN(new_n714));
  AOI211_X1 g528(.A(KEYINPUT32), .B(new_n575), .C1(new_n577), .C2(new_n578), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n598), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n524), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n697), .A2(new_n698), .ZN(new_n718));
  AOI21_X1  g532(.A(KEYINPUT103), .B1(new_n706), .B2(new_n189), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n646), .B2(new_n648), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n255), .ZN(G18));
  AND3_X1   g536(.A1(new_n287), .A2(new_n658), .A3(new_n394), .ZN(new_n723));
  INV_X1    g537(.A(new_n697), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n643), .A3(new_n716), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  AOI21_X1  g540(.A(new_n547), .B1(new_n553), .B2(new_n594), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n577), .A2(new_n549), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n574), .B(KEYINPUT104), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n577), .B2(new_n578), .ZN(new_n732));
  INV_X1    g546(.A(G472), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n729), .A2(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n734), .A2(new_n709), .A3(new_n524), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n662), .A2(new_n681), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n708), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n734), .A2(new_n668), .ZN(new_n739));
  INV_X1    g553(.A(new_n665), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n634), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n643), .A2(new_n724), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n217), .ZN(G27));
  NOR2_X1   g558(.A1(new_n385), .A2(new_n387), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n362), .A2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(KEYINPUT105), .B(new_n291), .C1(new_n353), .C2(new_n361), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n376), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n384), .B1(new_n749), .B2(new_n191), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n189), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n468), .A2(new_n476), .A3(new_n474), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n693), .A2(new_n599), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n693), .A2(new_n599), .A3(new_n753), .A4(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G131), .ZN(G33));
  NAND3_X1  g573(.A1(new_n599), .A2(new_n753), .A3(new_n666), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND4_X1  g575(.A1(new_n747), .A2(KEYINPUT45), .A3(new_n376), .A4(new_n748), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(G469), .C1(KEYINPUT45), .C2(new_n377), .ZN(new_n763));
  NAND2_X1  g577(.A1(G469), .A2(G902), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT46), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n745), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n764), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n189), .A3(new_n678), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n249), .B1(new_n631), .B2(new_n633), .ZN(new_n770));
  AND2_X1   g584(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n652), .A3(new_n658), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n769), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n752), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n778), .B(new_n779), .C1(new_n777), .C2(new_n776), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  AOI21_X1  g595(.A(new_n611), .B1(new_n766), .B2(new_n767), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n693), .A3(new_n779), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n786), .A2(new_n716), .A3(new_n717), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NOR3_X1   g602(.A1(new_n752), .A2(new_n391), .A3(new_n697), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n775), .A2(new_n599), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT48), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n775), .A2(new_n739), .A3(new_n789), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n792), .B1(KEYINPUT116), .B2(KEYINPUT51), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n734), .A2(new_n524), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n794), .B1(new_n772), .B2(new_n774), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n697), .A2(new_n391), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n478), .A3(new_n689), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT50), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT115), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n793), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n688), .A2(new_n789), .A3(new_n717), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n631), .A2(new_n615), .A3(new_n633), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n706), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n783), .B(new_n784), .C1(new_n189), .C2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n391), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n779), .A4(new_n795), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n802), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n802), .A2(new_n813), .A3(new_n805), .A4(new_n809), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n803), .A2(new_n635), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n791), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n711), .A2(new_n737), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n648), .A2(new_n646), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n599), .A3(new_n708), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n819), .A2(KEYINPUT108), .A3(new_n821), .A4(new_n725), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n711), .A2(new_n737), .A3(new_n725), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n823), .B1(new_n824), .B2(new_n721), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(new_n758), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n635), .A2(new_n647), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n662), .A2(KEYINPUT82), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n643), .A2(new_n396), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n709), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n610), .A2(new_n612), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n659), .A2(new_n831), .A3(new_n600), .ZN(new_n832));
  INV_X1    g646(.A(new_n753), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT109), .B1(new_n741), .B2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n693), .A2(new_n739), .A3(new_n753), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n189), .A2(new_n388), .A3(new_n658), .A4(new_n740), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n287), .A3(new_n716), .A4(new_n779), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n837), .A2(new_n760), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n826), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n745), .A2(new_n750), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n688), .A2(new_n658), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n189), .A3(new_n740), .A4(new_n736), .ZN(new_n846));
  INV_X1    g660(.A(new_n743), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n674), .A2(new_n694), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n743), .B1(new_n672), .B2(new_n673), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n846), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n822), .A2(new_n825), .A3(new_n758), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n760), .A2(new_n839), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n834), .B2(new_n836), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n600), .A3(new_n659), .A4(new_n831), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT110), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n843), .A2(new_n853), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT53), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n859), .A2(new_n861), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n859), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n857), .B(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n824), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n758), .A2(new_n869), .A3(new_n821), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT113), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(KEYINPUT53), .A3(new_n853), .A4(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n866), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n795), .A2(new_n643), .A3(new_n796), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n818), .A2(new_n864), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(G952), .B(new_n193), .C1(new_n877), .C2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  OAI21_X1  g693(.A(G953), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n612), .A2(new_n476), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT107), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n806), .A2(KEYINPUT49), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(new_n770), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n687), .B1(KEYINPUT49), .B2(new_n806), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n689), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n878), .A2(new_n880), .A3(new_n886), .ZN(G75));
  AOI21_X1  g701(.A(new_n191), .B1(new_n866), .B2(new_n872), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n426), .A2(new_n428), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(new_n435), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n889), .A2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n193), .A2(G952), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT118), .Z(new_n896));
  NOR3_X1   g710(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(G51));
  NAND2_X1  g711(.A1(new_n866), .A2(new_n872), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n873), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n875), .ZN(new_n901));
  INV_X1    g715(.A(new_n898), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n902), .A2(KEYINPUT119), .A3(new_n874), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n764), .B(KEYINPUT57), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n383), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n902), .A2(new_n191), .A3(new_n763), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n895), .B1(new_n906), .B2(new_n907), .ZN(G54));
  NAND4_X1  g722(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n909));
  OR2_X1    g723(.A1(new_n234), .A2(new_n240), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n895), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .A4(new_n910), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT120), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT120), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n912), .A2(new_n917), .A3(new_n913), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(G60));
  XOR2_X1   g733(.A(new_n627), .B(KEYINPUT121), .Z(new_n920));
  AND2_X1   g734(.A1(new_n864), .A2(new_n875), .ZN(new_n921));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT59), .Z(new_n923));
  OAI21_X1  g737(.A(new_n920), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n896), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n920), .A2(new_n923), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n901), .A2(new_n903), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT60), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n898), .A2(new_n656), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n866), .B2(new_n872), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n925), .C1(new_n521), .C2(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n934), .A2(KEYINPUT122), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n934), .B2(KEYINPUT122), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G66));
  AOI21_X1  g752(.A(new_n193), .B1(new_n392), .B2(G224), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n822), .A2(new_n825), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(new_n832), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n193), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT124), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n890), .B1(G898), .B2(new_n193), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  NOR2_X1   g759(.A1(new_n565), .A2(new_n567), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(new_n235), .Z(new_n947));
  NAND2_X1  g761(.A1(G900), .A2(G953), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n758), .A2(new_n760), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n851), .A2(new_n694), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n782), .A2(new_n599), .A3(new_n678), .A4(new_n736), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n953), .A2(new_n780), .A3(new_n787), .A4(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n947), .B(new_n948), .C1(new_n955), .C2(G953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n952), .A2(new_n690), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n827), .A2(KEYINPUT125), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n679), .B1(new_n827), .B2(KEYINPUT125), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n959), .A2(new_n960), .A3(new_n599), .A4(new_n779), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n958), .A2(new_n780), .A3(new_n787), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n962), .A2(new_n193), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n956), .B1(new_n963), .B2(new_n947), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G72));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n962), .B2(new_n941), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n570), .B(KEYINPUT127), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n547), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n968), .B1(new_n955), .B2(new_n941), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n973), .A2(new_n556), .A3(new_n970), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n913), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n862), .A2(new_n863), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n976), .B1(new_n548), .B2(new_n588), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n968), .B2(new_n977), .ZN(G57));
endmodule


