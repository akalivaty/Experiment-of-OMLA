

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n680), .A2(n690), .ZN(n682) );
  NOR2_X1 U554 ( .A1(G651), .A2(n560), .ZN(n778) );
  NOR2_X1 U555 ( .A1(n560), .A2(n518), .ZN(n783) );
  BUF_X2 U556 ( .A(n873), .Z(n515) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n524), .Z(n873) );
  XOR2_X2 U558 ( .A(KEYINPUT72), .B(n616), .Z(n937) );
  XNOR2_X1 U559 ( .A(n594), .B(KEYINPUT90), .ZN(n630) );
  AND2_X1 U560 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X2 U561 ( .A1(G164), .A2(G1384), .ZN(n696) );
  NAND2_X1 U562 ( .A1(G8), .A2(n658), .ZN(n690) );
  NOR2_X1 U563 ( .A1(n685), .A2(n684), .ZN(n686) );
  INV_X1 U564 ( .A(KEYINPUT93), .ZN(n640) );
  INV_X1 U565 ( .A(KEYINPUT28), .ZN(n631) );
  NOR2_X1 U566 ( .A1(n651), .A2(n650), .ZN(n652) );
  AND2_X1 U567 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n525), .ZN(n866) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n782) );
  NAND2_X1 U570 ( .A1(G88), .A2(n782), .ZN(n517) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n560) );
  XOR2_X1 U572 ( .A(KEYINPUT64), .B(G651), .Z(n518) );
  NAND2_X1 U573 ( .A1(G75), .A2(n783), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n517), .A2(n516), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n778), .A2(G50), .ZN(n521) );
  NOR2_X1 U576 ( .A1(G543), .A2(n518), .ZN(n519) );
  XOR2_X2 U577 ( .A(KEYINPUT1), .B(n519), .Z(n779) );
  NAND2_X1 U578 ( .A1(G62), .A2(n779), .ZN(n520) );
  NAND2_X1 U579 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n523), .A2(n522), .ZN(G166) );
  NOR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  NAND2_X1 U582 ( .A1(G138), .A2(n515), .ZN(n531) );
  INV_X1 U583 ( .A(G2105), .ZN(n525) );
  AND2_X2 U584 ( .A1(n525), .A2(G2104), .ZN(n872) );
  AND2_X1 U585 ( .A1(G102), .A2(n872), .ZN(n529) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n868) );
  NAND2_X1 U587 ( .A1(G114), .A2(n868), .ZN(n527) );
  NAND2_X1 U588 ( .A1(G126), .A2(n866), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  AND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(G164) );
  NAND2_X1 U592 ( .A1(n778), .A2(G52), .ZN(n532) );
  XNOR2_X1 U593 ( .A(KEYINPUT65), .B(n532), .ZN(n540) );
  NAND2_X1 U594 ( .A1(G90), .A2(n782), .ZN(n534) );
  NAND2_X1 U595 ( .A1(G77), .A2(n783), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U597 ( .A(n535), .B(KEYINPUT9), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(KEYINPUT66), .ZN(n538) );
  NAND2_X1 U599 ( .A1(G64), .A2(n779), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U601 ( .A1(n540), .A2(n539), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G53), .A2(n778), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n541), .Z(n546) );
  NAND2_X1 U604 ( .A1(G91), .A2(n782), .ZN(n543) );
  NAND2_X1 U605 ( .A1(G78), .A2(n783), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(n544), .Z(n545) );
  NOR2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n548) );
  NAND2_X1 U609 ( .A1(G65), .A2(n779), .ZN(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U611 ( .A1(n782), .A2(G89), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n549), .B(KEYINPUT4), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G76), .A2(n783), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n552), .B(KEYINPUT5), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n778), .A2(G51), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT74), .ZN(n555) );
  NAND2_X1 U618 ( .A1(G63), .A2(n779), .ZN(n554) );
  NAND2_X1 U619 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT6), .B(n556), .Z(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U624 ( .A(G166), .ZN(G303) );
  NAND2_X1 U625 ( .A1(G87), .A2(n560), .ZN(n562) );
  NAND2_X1 U626 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n779), .A2(n563), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n778), .A2(G49), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(G288) );
  NAND2_X1 U631 ( .A1(G86), .A2(n782), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G48), .A2(n778), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n783), .A2(G73), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT2), .B(n568), .Z(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G61), .A2(n779), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(G305) );
  NAND2_X1 U639 ( .A1(n778), .A2(G47), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G60), .A2(n779), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G85), .A2(n782), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G72), .A2(n783), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(G290) );
  NAND2_X1 U646 ( .A1(G8), .A2(G166), .ZN(n579) );
  NOR2_X1 U647 ( .A1(G2090), .A2(n579), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT99), .ZN(n669) );
  NAND2_X1 U649 ( .A1(n515), .A2(G137), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G101), .A2(n872), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT23), .B(n581), .Z(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n750) );
  INV_X1 U653 ( .A(G40), .ZN(n586) );
  NAND2_X1 U654 ( .A1(G113), .A2(n868), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G125), .A2(n866), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(n749) );
  OR2_X1 U657 ( .A1(n586), .A2(n749), .ZN(n587) );
  OR2_X1 U658 ( .A1(n750), .A2(n587), .ZN(n695) );
  INV_X1 U659 ( .A(n695), .ZN(n588) );
  NAND2_X2 U660 ( .A1(n588), .A2(n696), .ZN(n658) );
  NOR2_X1 U661 ( .A1(G1966), .A2(n690), .ZN(n651) );
  XNOR2_X1 U662 ( .A(G2078), .B(KEYINPUT25), .ZN(n918) );
  NOR2_X1 U663 ( .A1(n658), .A2(n918), .ZN(n590) );
  INV_X1 U664 ( .A(n658), .ZN(n603) );
  INV_X1 U665 ( .A(G1961), .ZN(n964) );
  NOR2_X1 U666 ( .A1(n603), .A2(n964), .ZN(n589) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n639) );
  NAND2_X1 U668 ( .A1(G171), .A2(n639), .ZN(n638) );
  INV_X1 U669 ( .A(G299), .ZN(n796) );
  NAND2_X1 U670 ( .A1(n603), .A2(G2072), .ZN(n591) );
  XOR2_X1 U671 ( .A(n591), .B(KEYINPUT27), .Z(n593) );
  NAND2_X1 U672 ( .A1(G1956), .A2(n658), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n796), .A2(n630), .ZN(n629) );
  NAND2_X1 U674 ( .A1(n782), .A2(G92), .ZN(n596) );
  NAND2_X1 U675 ( .A1(G66), .A2(n779), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n778), .A2(G54), .ZN(n598) );
  NAND2_X1 U678 ( .A1(G79), .A2(n783), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U680 ( .A(KEYINPUT73), .B(n599), .Z(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U682 ( .A(KEYINPUT15), .B(n602), .ZN(n940) );
  NAND2_X1 U683 ( .A1(G1348), .A2(n658), .ZN(n605) );
  NAND2_X1 U684 ( .A1(G2067), .A2(n603), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n622) );
  NOR2_X1 U686 ( .A1(n940), .A2(n622), .ZN(n627) );
  NAND2_X1 U687 ( .A1(G56), .A2(n779), .ZN(n606) );
  XNOR2_X1 U688 ( .A(n606), .B(KEYINPUT14), .ZN(n608) );
  NAND2_X1 U689 ( .A1(G43), .A2(n778), .ZN(n607) );
  NAND2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G68), .A2(n783), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n782), .A2(G81), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U694 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT71), .ZN(n613) );
  XNOR2_X1 U696 ( .A(KEYINPUT13), .B(n613), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U698 ( .A(G1996), .ZN(n731) );
  NOR2_X1 U699 ( .A1(n658), .A2(n731), .ZN(n618) );
  XNOR2_X1 U700 ( .A(KEYINPUT26), .B(KEYINPUT91), .ZN(n617) );
  XNOR2_X1 U701 ( .A(n618), .B(n617), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n658), .A2(G1341), .ZN(n619) );
  NAND2_X1 U703 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U704 ( .A(KEYINPUT92), .B(n621), .Z(n624) );
  NAND2_X1 U705 ( .A1(n940), .A2(n622), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n937), .A2(n625), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n796), .A2(n630), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U713 ( .A(n635), .B(KEYINPUT29), .ZN(n636) );
  INV_X1 U714 ( .A(n636), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n649) );
  NOR2_X1 U716 ( .A1(G171), .A2(n639), .ZN(n646) );
  NOR2_X1 U717 ( .A1(G2084), .A2(n658), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n653), .A2(n651), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n642), .A2(G8), .ZN(n643) );
  XNOR2_X1 U721 ( .A(KEYINPUT30), .B(n643), .ZN(n644) );
  NOR2_X1 U722 ( .A1(n644), .A2(G168), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT31), .B(n647), .Z(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n657) );
  INV_X1 U726 ( .A(n657), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n652), .B(KEYINPUT94), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n653), .A2(G8), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n668) );
  AND2_X1 U730 ( .A1(G286), .A2(G8), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n665) );
  INV_X1 U732 ( .A(G8), .ZN(n663) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n690), .ZN(n660) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n658), .ZN(n659) );
  NOR2_X1 U735 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n661), .A2(G303), .ZN(n662) );
  OR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n666), .B(KEYINPUT32), .ZN(n667) );
  NAND2_X1 U739 ( .A1(n668), .A2(n667), .ZN(n674) );
  NAND2_X1 U740 ( .A1(n669), .A2(n674), .ZN(n670) );
  NAND2_X1 U741 ( .A1(n670), .A2(n690), .ZN(n694) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n673) );
  NAND2_X1 U743 ( .A1(KEYINPUT33), .A2(n673), .ZN(n671) );
  XNOR2_X1 U744 ( .A(n671), .B(KEYINPUT97), .ZN(n678) );
  NOR2_X1 U745 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n948) );
  NAND2_X1 U747 ( .A1(n674), .A2(n948), .ZN(n676) );
  NAND2_X1 U748 ( .A1(G288), .A2(G1976), .ZN(n675) );
  XOR2_X1 U749 ( .A(KEYINPUT95), .B(n675), .Z(n944) );
  NAND2_X1 U750 ( .A1(n676), .A2(n944), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n680), .A2(KEYINPUT96), .ZN(n677) );
  NOR2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U753 ( .A1(n679), .A2(n690), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT96), .B(KEYINPUT33), .Z(n681) );
  NAND2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n957) );
  NAND2_X1 U757 ( .A1(n683), .A2(n957), .ZN(n684) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT98), .ZN(n692) );
  NOR2_X1 U759 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(KEYINPUT89), .ZN(n688) );
  XNOR2_X1 U761 ( .A(n688), .B(KEYINPUT24), .ZN(n689) );
  NOR2_X1 U762 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n707) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n743) );
  XNOR2_X1 U766 ( .A(KEYINPUT37), .B(G2067), .ZN(n741) );
  NAND2_X1 U767 ( .A1(G104), .A2(n872), .ZN(n698) );
  NAND2_X1 U768 ( .A1(G140), .A2(n515), .ZN(n697) );
  NAND2_X1 U769 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U770 ( .A(KEYINPUT34), .B(n699), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n866), .A2(G128), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n700), .B(KEYINPUT84), .ZN(n702) );
  NAND2_X1 U773 ( .A1(G116), .A2(n868), .ZN(n701) );
  NAND2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U775 ( .A(KEYINPUT35), .B(n703), .Z(n704) );
  NOR2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U777 ( .A(KEYINPUT36), .B(n706), .ZN(n887) );
  NOR2_X1 U778 ( .A1(n741), .A2(n887), .ZN(n990) );
  NAND2_X1 U779 ( .A1(n743), .A2(n990), .ZN(n739) );
  AND2_X1 U780 ( .A1(n707), .A2(n739), .ZN(n730) );
  NAND2_X1 U781 ( .A1(G107), .A2(n868), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G119), .A2(n866), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n709), .A2(n708), .ZN(n714) );
  NAND2_X1 U784 ( .A1(G95), .A2(n872), .ZN(n711) );
  NAND2_X1 U785 ( .A1(G131), .A2(n515), .ZN(n710) );
  NAND2_X1 U786 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U787 ( .A(KEYINPUT85), .B(n712), .Z(n713) );
  NOR2_X1 U788 ( .A1(n714), .A2(n713), .ZN(n881) );
  INV_X1 U789 ( .A(G1991), .ZN(n919) );
  NOR2_X1 U790 ( .A1(n881), .A2(n919), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n515), .A2(G141), .ZN(n722) );
  NAND2_X1 U792 ( .A1(G117), .A2(n868), .ZN(n716) );
  NAND2_X1 U793 ( .A1(G129), .A2(n866), .ZN(n715) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U795 ( .A(KEYINPUT86), .B(n717), .ZN(n720) );
  NAND2_X1 U796 ( .A1(n872), .A2(G105), .ZN(n718) );
  XOR2_X1 U797 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  NOR2_X1 U798 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U800 ( .A(KEYINPUT87), .B(n723), .ZN(n882) );
  NOR2_X1 U801 ( .A1(n882), .A2(n731), .ZN(n724) );
  NOR2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n1000) );
  INV_X1 U803 ( .A(n743), .ZN(n726) );
  NOR2_X1 U804 ( .A1(n1000), .A2(n726), .ZN(n734) );
  XNOR2_X1 U805 ( .A(KEYINPUT88), .B(n734), .ZN(n728) );
  XNOR2_X1 U806 ( .A(G1986), .B(G290), .ZN(n950) );
  AND2_X1 U807 ( .A1(n950), .A2(n743), .ZN(n727) );
  NOR2_X1 U808 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U809 ( .A1(n730), .A2(n729), .ZN(n746) );
  XOR2_X1 U810 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n738) );
  AND2_X1 U811 ( .A1(n731), .A2(n882), .ZN(n997) );
  NOR2_X1 U812 ( .A1(G1986), .A2(G290), .ZN(n732) );
  AND2_X1 U813 ( .A1(n919), .A2(n881), .ZN(n992) );
  NOR2_X1 U814 ( .A1(n732), .A2(n992), .ZN(n733) );
  NOR2_X1 U815 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U816 ( .A(n735), .B(KEYINPUT100), .ZN(n736) );
  NOR2_X1 U817 ( .A1(n997), .A2(n736), .ZN(n737) );
  XNOR2_X1 U818 ( .A(n738), .B(n737), .ZN(n740) );
  NAND2_X1 U819 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U820 ( .A1(n741), .A2(n887), .ZN(n999) );
  NAND2_X1 U821 ( .A1(n742), .A2(n999), .ZN(n744) );
  NAND2_X1 U822 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U823 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U824 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n747) );
  XNOR2_X1 U825 ( .A(n748), .B(n747), .ZN(G329) );
  AND2_X1 U826 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U827 ( .A(G860), .ZN(n759) );
  OR2_X1 U828 ( .A1(n759), .A2(n937), .ZN(G153) );
  INV_X1 U829 ( .A(G57), .ZN(G237) );
  INV_X1 U830 ( .A(G82), .ZN(G220) );
  NOR2_X1 U831 ( .A1(n750), .A2(n749), .ZN(G160) );
  NAND2_X1 U832 ( .A1(G7), .A2(G661), .ZN(n751) );
  XNOR2_X1 U833 ( .A(n751), .B(KEYINPUT10), .ZN(n752) );
  XNOR2_X1 U834 ( .A(KEYINPUT70), .B(n752), .ZN(G223) );
  INV_X1 U835 ( .A(G223), .ZN(n818) );
  NAND2_X1 U836 ( .A1(n818), .A2(G567), .ZN(n753) );
  XOR2_X1 U837 ( .A(KEYINPUT11), .B(n753), .Z(G234) );
  INV_X1 U838 ( .A(G171), .ZN(G301) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n755) );
  INV_X1 U840 ( .A(G868), .ZN(n800) );
  NAND2_X1 U841 ( .A1(n940), .A2(n800), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(G284) );
  NAND2_X1 U843 ( .A1(n796), .A2(n800), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT75), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n800), .A2(G286), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n758), .A2(n757), .ZN(G297) );
  NAND2_X1 U847 ( .A1(n759), .A2(G559), .ZN(n760) );
  INV_X1 U848 ( .A(n940), .ZN(n890) );
  NAND2_X1 U849 ( .A1(n760), .A2(n890), .ZN(n761) );
  XNOR2_X1 U850 ( .A(n761), .B(KEYINPUT76), .ZN(n762) );
  XNOR2_X1 U851 ( .A(KEYINPUT16), .B(n762), .ZN(G148) );
  NOR2_X1 U852 ( .A1(n937), .A2(G868), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G868), .A2(n890), .ZN(n763) );
  NOR2_X1 U854 ( .A1(G559), .A2(n763), .ZN(n764) );
  NOR2_X1 U855 ( .A1(n765), .A2(n764), .ZN(G282) );
  NAND2_X1 U856 ( .A1(G99), .A2(n872), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G111), .A2(n868), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT79), .B(n768), .Z(n775) );
  NAND2_X1 U860 ( .A1(n515), .A2(G135), .ZN(n769) );
  XNOR2_X1 U861 ( .A(KEYINPUT77), .B(n769), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n866), .A2(G123), .ZN(n770) );
  XOR2_X1 U863 ( .A(KEYINPUT18), .B(n770), .Z(n771) );
  NOR2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U865 ( .A(KEYINPUT78), .B(n773), .Z(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n991) );
  XOR2_X1 U867 ( .A(G2096), .B(n991), .Z(n776) );
  NOR2_X1 U868 ( .A1(G2100), .A2(n776), .ZN(n777) );
  XOR2_X1 U869 ( .A(KEYINPUT80), .B(n777), .Z(G156) );
  NAND2_X1 U870 ( .A1(n778), .A2(G55), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G67), .A2(n779), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G93), .A2(n782), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G80), .A2(n783), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  OR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n801) );
  NAND2_X1 U877 ( .A1(n890), .A2(G559), .ZN(n797) );
  XNOR2_X1 U878 ( .A(n937), .B(n797), .ZN(n788) );
  NOR2_X1 U879 ( .A1(G860), .A2(n788), .ZN(n789) );
  XOR2_X1 U880 ( .A(n801), .B(n789), .Z(G145) );
  XNOR2_X1 U881 ( .A(KEYINPUT19), .B(G305), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n790), .B(G288), .ZN(n791) );
  XOR2_X1 U883 ( .A(n801), .B(n791), .Z(n793) );
  XNOR2_X1 U884 ( .A(G290), .B(G166), .ZN(n792) );
  XNOR2_X1 U885 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n937), .B(n794), .ZN(n795) );
  XNOR2_X1 U887 ( .A(n796), .B(n795), .ZN(n889) );
  XNOR2_X1 U888 ( .A(n889), .B(n797), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n798), .A2(G868), .ZN(n799) );
  XOR2_X1 U890 ( .A(KEYINPUT81), .B(n799), .Z(n803) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(G295) );
  NAND2_X1 U893 ( .A1(G2084), .A2(G2078), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT20), .B(n804), .Z(n805) );
  NAND2_X1 U895 ( .A1(n805), .A2(G2090), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n806), .B(KEYINPUT21), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT82), .B(n807), .ZN(n808) );
  NAND2_X1 U898 ( .A1(G2072), .A2(n808), .ZN(G158) );
  XNOR2_X1 U899 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U901 ( .A1(G220), .A2(G219), .ZN(n810) );
  XNOR2_X1 U902 ( .A(KEYINPUT22), .B(KEYINPUT83), .ZN(n809) );
  XNOR2_X1 U903 ( .A(n810), .B(n809), .ZN(n811) );
  NOR2_X1 U904 ( .A1(n811), .A2(G218), .ZN(n812) );
  NAND2_X1 U905 ( .A1(G96), .A2(n812), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n822), .ZN(n816) );
  NAND2_X1 U907 ( .A1(G69), .A2(G120), .ZN(n813) );
  NOR2_X1 U908 ( .A1(G237), .A2(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(G108), .A2(n814), .ZN(n823) );
  NAND2_X1 U910 ( .A1(G567), .A2(n823), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n843) );
  NAND2_X1 U912 ( .A1(G483), .A2(G661), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n843), .A2(n817), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(G36), .ZN(G176) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U917 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n821), .A2(n820), .ZN(G188) );
  NOR2_X1 U920 ( .A1(n823), .A2(n822), .ZN(G325) );
  XNOR2_X1 U921 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  XNOR2_X1 U922 ( .A(G1996), .B(KEYINPUT41), .ZN(n833) );
  XOR2_X1 U923 ( .A(G1981), .B(G1966), .Z(n825) );
  XNOR2_X1 U924 ( .A(G1991), .B(G1986), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U926 ( .A(G1976), .B(G1971), .Z(n827) );
  XNOR2_X1 U927 ( .A(G1961), .B(G1956), .ZN(n826) );
  XNOR2_X1 U928 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U929 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U930 ( .A(KEYINPUT108), .B(G2474), .ZN(n830) );
  XNOR2_X1 U931 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(G229) );
  XOR2_X1 U933 ( .A(G2678), .B(G2090), .Z(n835) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2072), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n836), .B(G2100), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2084), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT107), .Z(n840) );
  XNOR2_X1 U940 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(G227) );
  XOR2_X1 U943 ( .A(KEYINPUT106), .B(n843), .Z(G319) );
  NAND2_X1 U944 ( .A1(G124), .A2(n866), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n844), .B(KEYINPUT44), .ZN(n847) );
  NAND2_X1 U946 ( .A1(G112), .A2(n868), .ZN(n845) );
  XOR2_X1 U947 ( .A(KEYINPUT109), .B(n845), .Z(n846) );
  NAND2_X1 U948 ( .A1(n847), .A2(n846), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G100), .A2(n872), .ZN(n849) );
  NAND2_X1 U950 ( .A1(G136), .A2(n515), .ZN(n848) );
  NAND2_X1 U951 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U952 ( .A1(n851), .A2(n850), .ZN(G162) );
  XOR2_X1 U953 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n853) );
  XNOR2_X1 U954 ( .A(G164), .B(KEYINPUT114), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U956 ( .A(n854), .B(G162), .Z(n865) );
  XNOR2_X1 U957 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G115), .A2(n868), .ZN(n856) );
  NAND2_X1 U959 ( .A1(G127), .A2(n866), .ZN(n855) );
  NAND2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n515), .A2(G139), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT112), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G103), .A2(n872), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n1001) );
  XNOR2_X1 U967 ( .A(G160), .B(n1001), .ZN(n864) );
  XNOR2_X1 U968 ( .A(n865), .B(n864), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G130), .A2(n866), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT110), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G118), .A2(n868), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT111), .B(n869), .Z(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n878) );
  NAND2_X1 U974 ( .A1(G106), .A2(n872), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n515), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U979 ( .A(n880), .B(n879), .Z(n884) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n991), .B(n885), .Z(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U984 ( .A1(G37), .A2(n888), .ZN(G395) );
  XOR2_X1 U985 ( .A(n889), .B(G286), .Z(n892) );
  XNOR2_X1 U986 ( .A(G171), .B(n890), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U988 ( .A1(G37), .A2(n893), .ZN(G397) );
  XNOR2_X1 U989 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G229), .A2(G227), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n909) );
  XNOR2_X1 U992 ( .A(G2438), .B(G2443), .ZN(n905) );
  XOR2_X1 U993 ( .A(G2454), .B(G2430), .Z(n897) );
  XNOR2_X1 U994 ( .A(G2446), .B(KEYINPUT103), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U996 ( .A(G2451), .B(G2427), .Z(n899) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U1000 ( .A(G2435), .B(KEYINPUT104), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(n906), .A2(G14), .ZN(n912) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n912), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT115), .B(n907), .Z(n908) );
  NOR2_X1 U1006 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(G225) );
  XNOR2_X1 U1009 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n912), .ZN(G401) );
  INV_X1 U1016 ( .A(G29), .ZN(n1014) );
  XOR2_X1 U1017 ( .A(G34), .B(KEYINPUT121), .Z(n914) );
  XNOR2_X1 U1018 ( .A(G2084), .B(KEYINPUT54), .ZN(n913) );
  XNOR2_X1 U1019 ( .A(n914), .B(n913), .ZN(n931) );
  XOR2_X1 U1020 ( .A(G2090), .B(G35), .Z(n929) );
  XOR2_X1 U1021 ( .A(G2067), .B(G26), .Z(n915) );
  NAND2_X1 U1022 ( .A1(n915), .A2(G28), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(G1996), .B(G32), .ZN(n917) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n916) );
  NOR2_X1 U1025 ( .A1(n917), .A2(n916), .ZN(n923) );
  XOR2_X1 U1026 ( .A(n918), .B(G27), .Z(n921) );
  XOR2_X1 U1027 ( .A(n919), .B(G25), .Z(n920) );
  NOR2_X1 U1028 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1029 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1030 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1031 ( .A(KEYINPUT120), .B(n926), .Z(n927) );
  XNOR2_X1 U1032 ( .A(n927), .B(KEYINPUT53), .ZN(n928) );
  NAND2_X1 U1033 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n933) );
  XNOR2_X1 U1035 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n932) );
  XNOR2_X1 U1036 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n1014), .A2(n934), .ZN(n935) );
  NAND2_X1 U1038 ( .A1(n935), .A2(G11), .ZN(n936) );
  XNOR2_X1 U1039 ( .A(n936), .B(KEYINPUT123), .ZN(n1019) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n963) );
  XOR2_X1 U1041 ( .A(n937), .B(G1341), .Z(n939) );
  XNOR2_X1 U1042 ( .A(G171), .B(G1961), .ZN(n938) );
  NAND2_X1 U1043 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(G1348), .B(n940), .ZN(n941) );
  NOR2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(G1971), .A2(G303), .ZN(n943) );
  NAND2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1048 ( .A(G1956), .B(G299), .ZN(n945) );
  NOR2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(n951), .B(KEYINPUT126), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT127), .B(n954), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G168), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT124), .ZN(n956) );
  NAND2_X1 U1057 ( .A1(n957), .A2(n956), .ZN(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT125), .B(KEYINPUT57), .Z(n958) );
  XNOR2_X1 U1059 ( .A(n959), .B(n958), .ZN(n960) );
  NAND2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n988) );
  INV_X1 U1062 ( .A(G16), .ZN(n986) );
  XNOR2_X1 U1063 ( .A(G5), .B(n964), .ZN(n981) );
  XOR2_X1 U1064 ( .A(G1348), .B(KEYINPUT59), .Z(n965) );
  XNOR2_X1 U1065 ( .A(G4), .B(n965), .ZN(n967) );
  XNOR2_X1 U1066 ( .A(G20), .B(G1956), .ZN(n966) );
  NOR2_X1 U1067 ( .A1(n967), .A2(n966), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(G1341), .B(G19), .ZN(n969) );
  XNOR2_X1 U1069 ( .A(G6), .B(G1981), .ZN(n968) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1072 ( .A(n972), .B(KEYINPUT60), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n974) );
  XNOR2_X1 U1074 ( .A(G23), .B(G1976), .ZN(n973) );
  NOR2_X1 U1075 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1076 ( .A(G1986), .B(G24), .Z(n975) );
  NAND2_X1 U1077 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1078 ( .A(KEYINPUT58), .B(n977), .ZN(n978) );
  NOR2_X1 U1079 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1080 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1081 ( .A(G21), .B(G1966), .ZN(n982) );
  NOR2_X1 U1082 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1083 ( .A(KEYINPUT61), .B(n984), .ZN(n985) );
  NAND2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n1017) );
  XOR2_X1 U1086 ( .A(G160), .B(G2084), .Z(n989) );
  NOR2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1090 ( .A(KEYINPUT118), .B(n995), .ZN(n1010) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n996) );
  NOR2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1093 ( .A(KEYINPUT51), .B(n998), .Z(n1008) );
  NAND2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1001), .Z(n1003) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1002) );
  NOR2_X1 U1097 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1004), .Z(n1005) );
  NOR2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT52), .B(n1011), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(KEYINPUT55), .A2(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1105 ( .A(KEYINPUT119), .B(n1015), .Z(n1016) );
  NOR2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

