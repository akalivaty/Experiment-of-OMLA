//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT68), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT70), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n459), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(G137), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n465), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(new_n466), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR4_X1   g064(.A1(new_n471), .A2(KEYINPUT4), .A3(new_n489), .A4(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n463), .A2(G138), .A3(new_n466), .A4(new_n464), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(KEYINPUT4), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(new_n466), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n492), .A2(new_n497), .ZN(G164));
  NAND2_X1  g073(.A1(G75), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT5), .B1(new_n500), .B2(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT72), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n502), .A2(new_n503), .A3(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n505), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n510), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n508), .A2(new_n509), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(new_n516), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n500), .B1(new_n515), .B2(KEYINPUT74), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n512), .A2(new_n514), .A3(new_n529), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n528), .A2(G51), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n505), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n528), .A2(G52), .A3(new_n530), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n505), .A2(new_n515), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NOR2_X1   g116(.A1(new_n513), .A2(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT74), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(G543), .A3(new_n530), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n505), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n538), .A2(G81), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n505), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n544), .A2(G53), .A3(G543), .A4(new_n530), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  INV_X1    g144(.A(new_n567), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n528), .A2(G53), .A3(new_n530), .A4(new_n570), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n569), .B1(new_n568), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n564), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g151(.A(KEYINPUT77), .B(new_n564), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  XNOR2_X1  g154(.A(G166), .B(KEYINPUT78), .ZN(G303));
  NAND2_X1  g155(.A1(new_n546), .A2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n538), .A2(G87), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n505), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(G48), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n505), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n515), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n538), .A2(G85), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n545), .B2(new_n598), .C1(new_n599), .C2(new_n511), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n538), .A2(G92), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n538), .A2(new_n606), .A3(G92), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n505), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n546), .A2(G54), .B1(G651), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g188(.A(KEYINPUT10), .B1(new_n605), .B2(new_n607), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n603), .B1(new_n615), .B2(G868), .ZN(G284));
  OAI21_X1  g191(.A(new_n603), .B1(new_n615), .B2(G868), .ZN(G321));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(G299), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n618), .B2(G168), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n553), .A2(new_n618), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n622), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT82), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n626), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g203(.A1(new_n480), .A2(KEYINPUT84), .A3(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G135), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT84), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n479), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n629), .A2(new_n630), .A3(new_n633), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n466), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT85), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2072), .B(G2078), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n669), .A2(KEYINPUT17), .A3(new_n666), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n669), .B2(KEYINPUT17), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n670), .A2(new_n671), .A3(new_n665), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XOR2_X1   g251(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(G1956), .B(G2474), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  AND2_X1   g261(.A1(new_n681), .A2(KEYINPUT89), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n681), .A2(KEYINPUT89), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n678), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G1991), .ZN(new_n692));
  INV_X1    g267(.A(G1991), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n686), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G1996), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(G1996), .B1(new_n692), .B2(new_n694), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n697), .B2(new_n699), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n705), .B1(new_n703), .B2(new_n704), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT26), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(new_n713), .B1(G105), .B2(new_n475), .ZN(new_n714));
  INV_X1    g289(.A(G141), .ZN(new_n715));
  INV_X1    g290(.A(G129), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n714), .B1(new_n482), .B2(new_n715), .C1(new_n716), .C2(new_n479), .ZN(new_n717));
  MUX2_X1   g292(.A(G32), .B(new_n717), .S(G29), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT100), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(G301), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n720), .B1(G1961), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n554), .B2(new_n723), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1341), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G34), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n477), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G2084), .Z(new_n735));
  OR2_X1    g310(.A1(G29), .A2(G33), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT95), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n475), .A2(G103), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  AND2_X1   g314(.A1(new_n460), .A2(new_n470), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n740), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  INV_X1    g316(.A(G139), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n739), .B1(new_n466), .B2(new_n741), .C1(new_n482), .C2(new_n742), .ZN(new_n743));
  OAI221_X1 g318(.A(new_n736), .B1(new_n737), .B2(G2072), .C1(new_n743), .C2(new_n732), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n737), .A2(G2072), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NOR4_X1   g321(.A1(new_n726), .A2(new_n729), .A3(new_n735), .A4(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n732), .A2(G26), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n480), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n483), .A2(G140), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n466), .A2(G116), .ZN(new_n751));
  OAI21_X1  g326(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n748), .B1(new_n753), .B2(G29), .ZN(new_n754));
  MUX2_X1   g329(.A(new_n748), .B(new_n754), .S(KEYINPUT28), .Z(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2067), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n747), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n732), .A2(G27), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT102), .Z(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n732), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT104), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT103), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n615), .A2(new_n723), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G4), .B2(new_n723), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT93), .B(G1348), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n768), .B2(new_n766), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n757), .A2(new_n764), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n480), .A2(KEYINPUT91), .A3(G119), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n483), .A2(G131), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n781));
  INV_X1    g356(.A(G119), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n479), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(G95), .A2(G2105), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n784), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n779), .A2(new_n780), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G25), .B(new_n786), .S(G29), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT35), .B(G1991), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G1986), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n723), .A2(G24), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G290), .B2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(G288), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT33), .B(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n723), .A2(G22), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G166), .B2(new_n723), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1971), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n723), .A2(G6), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n595), .B2(new_n723), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n798), .A2(new_n801), .A3(new_n802), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n792), .A2(new_n790), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n793), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT36), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT23), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n723), .A2(G20), .ZN(new_n815));
  AOI211_X1 g390(.A(new_n814), .B(new_n815), .C1(G299), .C2(G16), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  INV_X1    g392(.A(G1956), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n723), .A2(G21), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G168), .B2(new_n723), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G1966), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n822), .A2(G1966), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT31), .B(G11), .ZN(new_n826));
  INV_X1    g401(.A(G28), .ZN(new_n827));
  AOI21_X1  g402(.A(G29), .B1(new_n827), .B2(KEYINPUT30), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(KEYINPUT30), .B2(new_n827), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n826), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n636), .A2(new_n732), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n725), .A2(G1961), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n835), .B(new_n836), .C1(new_n834), .C2(new_n833), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n824), .A2(new_n825), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT101), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n778), .A2(new_n813), .A3(new_n819), .A4(new_n839), .ZN(G150));
  INV_X1    g415(.A(G150), .ZN(G311));
  NAND2_X1  g416(.A1(new_n615), .A2(G559), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(new_n511), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n538), .A2(G93), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n544), .A2(G55), .A3(G543), .A4(new_n530), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n847), .A2(KEYINPUT106), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT106), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n554), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n553), .B(new_n846), .C1(new_n850), .C2(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n844), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XOR2_X1   g435(.A(new_n786), .B(new_n639), .Z(new_n861));
  INV_X1    g436(.A(G142), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT109), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n863), .A2(new_n466), .A3(G118), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n466), .B2(G118), .ZN(new_n865));
  OR2_X1    g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(G2104), .A3(new_n866), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n482), .A2(new_n862), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(G130), .B2(new_n480), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n861), .B(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n492), .A2(new_n497), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n717), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n753), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n743), .B(KEYINPUT108), .Z(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n871), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n870), .B1(new_n881), .B2(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n487), .B(KEYINPUT107), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(G160), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n636), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT110), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  INV_X1    g466(.A(new_n886), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n882), .A3(new_n880), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g470(.A1(new_n626), .A2(new_n855), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n626), .A2(new_n855), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT111), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n576), .A2(new_n577), .A3(new_n615), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n615), .B1(new_n576), .B2(new_n577), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT41), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n615), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n568), .A2(new_n571), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT76), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT77), .B1(new_n907), .B2(new_n564), .ZN(new_n908));
  INV_X1    g483(.A(new_n577), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n576), .A2(new_n577), .A3(new_n615), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n899), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT111), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n898), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n900), .A2(new_n901), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n896), .A2(new_n897), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n921));
  XNOR2_X1  g496(.A(G290), .B(G288), .ZN(new_n922));
  XNOR2_X1  g497(.A(G166), .B(G305), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n922), .B(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n917), .A2(new_n926), .A3(new_n919), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n921), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n921), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n851), .A2(new_n618), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(G295));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n931), .ZN(G331));
  NOR2_X1   g508(.A1(G171), .A2(KEYINPUT112), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n536), .A2(new_n537), .A3(new_n539), .A4(KEYINPUT112), .ZN(new_n935));
  NAND2_X1  g510(.A1(G168), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT113), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT113), .ZN(new_n938));
  NAND3_X1  g513(.A1(G168), .A2(new_n938), .A3(new_n935), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n854), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n852), .A3(new_n853), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n934), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n934), .A3(new_n942), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n914), .B2(new_n916), .ZN(new_n947));
  INV_X1    g522(.A(new_n945), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(new_n943), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n918), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n925), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT114), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n947), .A2(new_n925), .A3(KEYINPUT114), .A4(new_n950), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT41), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT111), .B1(new_n955), .B2(new_n915), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n902), .A2(new_n899), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n949), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n949), .A2(new_n918), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n924), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n953), .A2(new_n891), .A3(new_n954), .A4(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n951), .B2(new_n952), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n949), .B1(new_n902), .B2(new_n913), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n924), .B1(new_n965), .B2(new_n959), .ZN(new_n966));
  AND4_X1   g541(.A1(KEYINPUT43), .A2(new_n964), .A3(new_n954), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n964), .A2(new_n962), .A3(new_n954), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(G397));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n492), .B2(new_n497), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n467), .A2(G40), .A3(new_n474), .A4(new_n476), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n753), .B(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT115), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(new_n717), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(KEYINPUT46), .A3(new_n696), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n986));
  INV_X1    g561(.A(new_n980), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(new_n987), .B2(G1996), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n717), .B(new_n696), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n786), .A2(new_n788), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n992), .A2(new_n993), .B1(G2067), .B2(new_n753), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n980), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n786), .B(new_n788), .Z(new_n997));
  AOI21_X1  g572(.A(new_n987), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n987), .A2(G1986), .A3(G290), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n995), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n990), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  INV_X1    g578(.A(new_n976), .ZN(new_n1004));
  INV_X1    g579(.A(new_n979), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT121), .Z(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT119), .B(G1981), .Z(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n595), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n595), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT49), .ZN(new_n1013));
  AOI211_X1 g588(.A(G1976), .B(G288), .C1(new_n1013), .C2(new_n1006), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1010), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1007), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1013), .A2(new_n1006), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n795), .A2(G1976), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1006), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1006), .A2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1017), .A2(KEYINPUT120), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  AND2_X1   g603(.A1(G166), .A2(KEYINPUT78), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G166), .A2(KEYINPUT78), .ZN(new_n1030));
  OAI211_X1 g605(.A(KEYINPUT55), .B(G8), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT118), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND4_X1  g611(.A1(G303), .A2(new_n1036), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT45), .B(new_n975), .C1(new_n492), .C2(new_n497), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n978), .A2(new_n1039), .A3(new_n1005), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n978), .A2(new_n1039), .A3(new_n1005), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT117), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n872), .A2(new_n1046), .A3(new_n975), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n979), .B1(new_n976), .B2(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1038), .B(G8), .C1(new_n1045), .C2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1016), .B1(new_n1028), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1032), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1024), .ZN(new_n1056));
  AND4_X1   g631(.A1(KEYINPUT62), .A2(new_n1051), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1043), .B(new_n1041), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n1058), .B2(new_n763), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n763), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1049), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1060), .B1(G1961), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G171), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1966), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1043), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT122), .B(G2084), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1047), .A2(new_n1048), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(G168), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1003), .A2(KEYINPUT126), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1068), .A2(KEYINPUT51), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT51), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G8), .ZN(new_n1073));
  OAI22_X1  g648(.A1(new_n1070), .A2(new_n1071), .B1(G168), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1063), .B1(new_n1074), .B2(KEYINPUT62), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1052), .B1(new_n1057), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1053), .B(new_n1038), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1073), .A2(G286), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(KEYINPUT63), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1051), .A2(new_n1055), .A3(new_n1056), .A4(new_n1078), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1076), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1075), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1043), .B2(G1996), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n979), .B1(new_n976), .B2(new_n977), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(KEYINPUT124), .A3(new_n696), .A4(new_n1039), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1087), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT125), .B(new_n1095), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n554), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT59), .B(new_n554), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1040), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1049), .A2(new_n818), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n574), .A2(KEYINPUT57), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n904), .A2(new_n1107), .A3(new_n564), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1090), .A2(new_n1039), .A3(new_n1103), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1956), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT61), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1104), .A2(new_n1105), .A3(KEYINPUT123), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(new_n1110), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1109), .A2(KEYINPUT61), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G2067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n768), .B2(new_n1049), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n615), .B1(new_n1123), .B2(KEYINPUT60), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1101), .A2(new_n1102), .A3(new_n1120), .A4(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1118), .B1(new_n903), .B2(new_n1123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1109), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1063), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1059), .A2(G171), .A3(new_n1062), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT54), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1134), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1063), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1086), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1077), .A2(new_n1074), .A3(new_n1056), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1085), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(G290), .B(G1986), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n998), .B1(new_n980), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT116), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1002), .B1(new_n1142), .B2(new_n1145), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g721(.A(new_n457), .ZN(new_n1148));
  NOR2_X1   g722(.A1(G227), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g723(.A1(new_n660), .A2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g724(.A(new_n1150), .B(KEYINPUT127), .Z(new_n1151));
  AND2_X1   g725(.A1(new_n708), .A2(new_n1151), .ZN(new_n1152));
  AND3_X1   g726(.A1(new_n1152), .A2(new_n971), .A3(new_n894), .ZN(G308));
  NAND3_X1  g727(.A1(new_n1152), .A2(new_n971), .A3(new_n894), .ZN(G225));
endmodule


