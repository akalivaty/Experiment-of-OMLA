//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AND2_X1   g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n456), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XOR2_X1   g046(.A(new_n471), .B(KEYINPUT69), .Z(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(new_n467), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n465), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT71), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n474), .A2(G136), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT70), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n465), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n480), .B(new_n482), .C1(G124), .C2(new_n483), .ZN(G162));
  NAND2_X1  g059(.A1(new_n474), .A2(G138), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT4), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n483), .B2(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G543), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT73), .B1(new_n495), .B2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(new_n493), .A3(G543), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT72), .B(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT72), .B(G651), .Z(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(new_n503), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n495), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n505), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n511), .A2(new_n500), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(G166));
  OAI211_X1 g088(.A(G51), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  OAI211_X1 g092(.A(new_n514), .B(new_n516), .C1(new_n504), .C2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n494), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n497), .B1(new_n493), .B2(G543), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n495), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n499), .A2(new_n524), .ZN(new_n525));
  AND4_X1   g100(.A1(G63), .A2(new_n523), .A3(G651), .A4(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n518), .A2(new_n526), .ZN(G168));
  XOR2_X1   g102(.A(KEYINPUT76), .B(G90), .Z(new_n528));
  AOI22_X1  g103(.A1(new_n505), .A2(new_n528), .B1(new_n509), .B2(G52), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(G64), .A3(new_n525), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n500), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n529), .B1(new_n532), .B2(KEYINPUT75), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n534));
  AOI211_X1 g109(.A(new_n534), .B(new_n500), .C1(new_n530), .C2(new_n531), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  OAI211_X1 g111(.A(G43), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n537));
  OAI211_X1 g112(.A(G81), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G68), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n495), .ZN(new_n542));
  AOI211_X1 g117(.A(KEYINPUT74), .B(new_n494), .C1(new_n496), .C2(new_n498), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n496), .A2(new_n498), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n524), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n542), .B1(new_n546), .B2(G56), .ZN(new_n547));
  OAI211_X1 g122(.A(KEYINPUT77), .B(new_n540), .C1(new_n547), .C2(new_n500), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n523), .A2(G56), .A3(new_n525), .ZN(new_n550));
  INV_X1    g125(.A(new_n542), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n500), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n549), .B1(new_n552), .B2(new_n539), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT79), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n563));
  OAI21_X1  g138(.A(G543), .B1(new_n502), .B2(new_n503), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n507), .A2(new_n508), .ZN(new_n567));
  INV_X1    g142(.A(new_n563), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(G53), .A3(G543), .A4(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n566), .A2(new_n569), .B1(new_n505), .B2(G91), .ZN(new_n570));
  INV_X1    g145(.A(G651), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT81), .B(G65), .Z(new_n572));
  AOI22_X1  g147(.A1(new_n499), .A2(new_n572), .B1(G78), .B2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n571), .B1(new_n573), .B2(KEYINPUT82), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n574), .B1(KEYINPUT82), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  OR2_X1    g152(.A1(new_n518), .A2(new_n526), .ZN(G286));
  XOR2_X1   g153(.A(G166), .B(KEYINPUT83), .Z(G303));
  NAND2_X1  g154(.A1(new_n523), .A2(new_n525), .ZN(new_n580));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n571), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G49), .ZN(new_n583));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n583), .A2(new_n564), .B1(new_n504), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT84), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n564), .B1(new_n504), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n500), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n591), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n595), .A2(new_n500), .ZN(new_n596));
  INV_X1    g171(.A(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(new_n564), .B1(new_n504), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G290));
  OAI211_X1 g176(.A(G92), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT85), .B(G66), .Z(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n522), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(G54), .A2(new_n509), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G171), .B2(new_n610), .ZN(G284));
  OAI21_X1  g187(.A(new_n611), .B1(G171), .B2(new_n610), .ZN(G321));
  NAND2_X1  g188(.A1(G299), .A2(new_n610), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n610), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(new_n609), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n554), .B2(G868), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n468), .A2(new_n475), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  INV_X1    g201(.A(G2100), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n474), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n483), .A2(G123), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND3_X1  g210(.A1(new_n628), .A2(new_n629), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT86), .Z(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(G14), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(KEYINPUT17), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n662), .A2(new_n655), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n656), .A2(new_n655), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n661), .B(new_n664), .C1(new_n659), .C2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT89), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n675), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n677), .B(new_n680), .C1(new_n672), .C2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT91), .Z(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G6), .ZN(new_n692));
  INV_X1    g267(.A(G305), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT95), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT32), .B(G1981), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n586), .A2(new_n691), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n691), .B2(G23), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT33), .B(G1976), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G22), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT96), .Z(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n691), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT97), .B(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n700), .B2(new_n701), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n697), .A2(new_n702), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n691), .A2(G24), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n600), .B2(new_n691), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT94), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n483), .A2(G119), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G107), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G2105), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n474), .B2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n709), .B2(new_n710), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n716), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT36), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT99), .B(KEYINPUT25), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G139), .B2(new_n474), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n465), .B2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G33), .B(new_n736), .S(G29), .Z(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT100), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2072), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT101), .Z(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G32), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n474), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n483), .A2(G129), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n743), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT102), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n742), .B1(new_n749), .B2(new_n741), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT103), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n738), .A2(G2072), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n750), .B2(new_n752), .ZN(new_n756));
  AND2_X1   g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n741), .B1(KEYINPUT24), .B2(G34), .ZN(new_n758));
  OAI22_X1  g333(.A1(G160), .A2(new_n741), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n740), .A2(new_n754), .A3(new_n756), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n691), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n691), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n764), .A2(G1961), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G1961), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G29), .A2(G35), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G162), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT105), .B(KEYINPUT29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G2090), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT106), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n691), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  NAND2_X1  g353(.A1(G164), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G27), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G2078), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT31), .B(G11), .Z(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n785), .A2(KEYINPUT30), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT104), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n783), .B(new_n789), .C1(new_n741), .C2(new_n634), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  NOR2_X1   g366(.A1(G168), .A2(new_n691), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n691), .B2(G21), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n782), .B(new_n790), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n791), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n771), .B2(new_n772), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n774), .A2(new_n778), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n554), .A2(new_n691), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n691), .B2(G19), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1341), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1341), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n691), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n617), .B2(new_n691), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1348), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n741), .A2(G26), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT28), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n474), .A2(G140), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n483), .A2(G128), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n465), .A2(G116), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n807), .B1(new_n812), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2067), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n801), .A2(new_n802), .A3(new_n805), .A4(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n767), .A2(new_n797), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n730), .A2(new_n819), .ZN(G311));
  OR2_X1    g395(.A1(new_n730), .A2(new_n819), .ZN(G150));
  NOR2_X1   g396(.A1(new_n609), .A2(new_n618), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  OAI211_X1 g398(.A(G55), .B(G543), .C1(new_n502), .C2(new_n503), .ZN(new_n824));
  INV_X1    g399(.A(G93), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n504), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n546), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n500), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n548), .A2(new_n553), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT107), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n540), .B1(new_n547), .B2(new_n500), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  INV_X1    g408(.A(G67), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n580), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n826), .B1(new_n835), .B2(new_n506), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n831), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n548), .A2(new_n553), .A3(new_n829), .A4(new_n831), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n823), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT108), .ZN(new_n843));
  AOI21_X1  g418(.A(G860), .B1(new_n841), .B2(KEYINPUT39), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n829), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n748), .B(new_n491), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n474), .A2(G142), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n483), .A2(G130), .ZN(new_n851));
  OR2_X1    g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n849), .B(new_n854), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n812), .B(KEYINPUT109), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n736), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n723), .B(new_n625), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n849), .B(new_n854), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(new_n634), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G162), .ZN(new_n866));
  AOI21_X1  g441(.A(G37), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n868), .A3(new_n863), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g446(.A1(new_n836), .A2(G868), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n586), .B(KEYINPUT110), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n693), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n600), .B(G166), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT42), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n840), .B(new_n620), .Z(new_n878));
  NAND2_X1  g453(.A1(G299), .A2(new_n609), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n570), .A2(new_n575), .A3(new_n604), .A4(new_n608), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(KEYINPUT41), .A3(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n880), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n883), .B1(new_n885), .B2(new_n878), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n877), .B(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n872), .B1(new_n887), .B2(G868), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT111), .ZN(G295));
  INV_X1    g464(.A(new_n888), .ZN(G331));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n891));
  OAI21_X1  g466(.A(G286), .B1(new_n533), .B2(new_n535), .ZN(new_n892));
  INV_X1    g467(.A(new_n531), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n546), .B2(G64), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n534), .B1(new_n894), .B2(new_n500), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n895), .A2(new_n896), .A3(G168), .A4(new_n529), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n840), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n882), .A2(new_n881), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n838), .A2(new_n898), .A3(new_n839), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n884), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT113), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT113), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n874), .A2(new_n875), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n874), .A2(new_n875), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n838), .A2(new_n898), .A3(new_n839), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n898), .B1(new_n838), .B2(new_n839), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n885), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n907), .B1(new_n918), .B2(new_n906), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT113), .B1(new_n920), .B2(new_n901), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n915), .B1(new_n922), .B2(new_n876), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n905), .A2(new_n876), .A3(new_n908), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n906), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n912), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n891), .B1(new_n924), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n912), .B1(new_n919), .B2(new_n921), .ZN(new_n931));
  INV_X1    g506(.A(G37), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n915), .A2(new_n933), .B1(new_n923), .B2(new_n927), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n891), .B2(new_n934), .ZN(G397));
  AND3_X1   g510(.A1(new_n472), .A2(G40), .A3(new_n476), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n491), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(G1996), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT114), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n940), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n812), .B(G2067), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n748), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT47), .Z(new_n949));
  AND2_X1   g524(.A1(new_n748), .A2(G1996), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(new_n946), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n942), .A2(new_n749), .B1(new_n945), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n718), .A2(new_n726), .A3(new_n722), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n812), .A2(G2067), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n940), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n940), .A2(G1986), .A3(G290), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n958), .B(KEYINPUT48), .Z(new_n959));
  AOI21_X1  g534(.A(new_n726), .B1(new_n718), .B2(new_n722), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n945), .B1(new_n960), .B2(new_n953), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n952), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n949), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n936), .A2(new_n938), .A3(new_n491), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(G8), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n967));
  OAI21_X1  g542(.A(G1981), .B1(new_n593), .B2(KEYINPUT116), .ZN(new_n968));
  XOR2_X1   g543(.A(G305), .B(new_n968), .Z(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n969), .A2(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1976), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n587), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT117), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(G305), .A2(G1981), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n966), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G303), .A2(G8), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n939), .A2(new_n937), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n936), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(KEYINPUT115), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n491), .A2(new_n991), .A3(new_n938), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n936), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n772), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n981), .A2(G8), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n582), .A2(new_n585), .A3(new_n973), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n966), .A2(KEYINPUT52), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n1000), .B1(G1976), .B2(new_n587), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT52), .B1(new_n966), .B2(new_n999), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n972), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n978), .B1(new_n998), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n997), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n996), .A2(G8), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n979), .B(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n994), .A2(new_n760), .B1(new_n984), .B2(new_n791), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(new_n1010), .A3(G286), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1011), .A2(KEYINPUT63), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1005), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n994), .A2(new_n772), .B1(new_n984), .B2(new_n985), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1014), .A2(KEYINPUT118), .ZN(new_n1015));
  OAI21_X1  g590(.A(G8), .B1(new_n1014), .B2(KEYINPUT118), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1003), .A2(new_n1017), .A3(new_n997), .A4(new_n1011), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT63), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1004), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT56), .B(G2072), .Z(new_n1022));
  OAI22_X1  g597(.A1(new_n994), .A2(G1956), .B1(new_n984), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g598(.A(G299), .B(KEYINPUT57), .Z(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n994), .A2(G1348), .B1(G2067), .B2(new_n965), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g604(.A(KEYINPUT119), .B1(new_n965), .B2(G2067), .C1(new_n994), .C2(G1348), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI221_X1 g606(.A(new_n1024), .B1(new_n984), .B2(new_n1022), .C1(new_n994), .C2(G1956), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n617), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1031), .A2(KEYINPUT60), .A3(new_n609), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n609), .B1(new_n1031), .B2(KEYINPUT60), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1035), .A2(new_n1036), .B1(KEYINPUT60), .B2(new_n1031), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT58), .B(G1341), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n965), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(G1996), .B2(new_n984), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1041), .B2(new_n554), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1041), .A2(new_n554), .ZN(new_n1043));
  AND2_X1   g618(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT61), .B1(new_n1032), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1026), .B(new_n1032), .C1(new_n1046), .C2(KEYINPUT61), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1045), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1034), .B1(new_n1037), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n984), .A2(G2078), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  INV_X1    g630(.A(G1961), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1054), .A2(new_n1055), .B1(new_n1056), .B2(new_n993), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n476), .A2(KEYINPUT53), .A3(G40), .A4(new_n781), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n471), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n982), .A2(new_n983), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1057), .A2(G301), .A3(new_n1060), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n984), .A2(new_n1055), .A3(G2078), .ZN(new_n1062));
  AOI21_X1  g637(.A(G301), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1053), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT123), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1010), .B1(new_n1009), .B2(G168), .ZN(new_n1066));
  NAND2_X1  g641(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1067));
  OR2_X1    g642(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1009), .A2(new_n1010), .A3(G168), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1069), .B(new_n1070), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1057), .A2(G301), .A3(new_n1062), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT54), .B(new_n1072), .C1(new_n1073), .C2(G301), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(new_n1053), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1065), .A2(new_n1071), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1063), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1071), .A2(KEYINPUT62), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1052), .A2(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1005), .A2(new_n1017), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1021), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n600), .B(G1986), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n962), .B1(new_n940), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n964), .B1(new_n1083), .B2(new_n1085), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n1088));
  NOR2_X1   g662(.A1(G227), .A2(new_n463), .ZN(new_n1089));
  XNOR2_X1  g663(.A(new_n1089), .B(KEYINPUT125), .ZN(new_n1090));
  NAND3_X1  g664(.A1(new_n1090), .A2(new_n653), .A3(new_n689), .ZN(new_n1091));
  INV_X1    g665(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g666(.A1(new_n870), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g667(.A(new_n1088), .B1(new_n934), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n867), .B2(new_n869), .ZN(new_n1095));
  AOI21_X1  g669(.A(new_n914), .B1(new_n913), .B2(new_n925), .ZN(new_n1096));
  AND3_X1   g670(.A1(new_n925), .A2(new_n927), .A3(new_n914), .ZN(new_n1097));
  OAI211_X1 g671(.A(KEYINPUT126), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AND3_X1   g672(.A1(new_n1094), .A2(KEYINPUT127), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g673(.A(KEYINPUT127), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1100));
  NOR2_X1   g674(.A1(new_n1099), .A2(new_n1100), .ZN(G308));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1098), .ZN(G225));
endmodule


