//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G214), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(G237), .A3(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT64), .A2(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT64), .A2(G143), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  INV_X1    g010(.A(G237), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(G214), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n193), .B2(KEYINPUT85), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT18), .ZN(new_n201));
  OAI22_X1  g015(.A1(new_n195), .A2(new_n200), .B1(KEYINPUT86), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n208), .B1(new_n205), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n203), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n206), .A2(G140), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n204), .A2(G125), .ZN(new_n213));
  OAI21_X1  g027(.A(G146), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(KEYINPUT87), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n195), .B2(new_n200), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(new_n198), .A3(G214), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT64), .B(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(KEYINPUT85), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT64), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n190), .B(new_n196), .C1(new_n223), .C2(new_n194), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n201), .A2(KEYINPUT86), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n222), .A2(new_n224), .A3(G131), .A4(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n202), .A2(new_n217), .A3(new_n219), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT88), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n222), .A2(new_n224), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n218), .A2(new_n230), .B1(new_n211), .B2(new_n216), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(KEYINPUT88), .A3(new_n226), .A4(new_n202), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n222), .A2(new_n224), .A3(G131), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n219), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT16), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n212), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n205), .A2(new_n207), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT19), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n235), .B(new_n239), .C1(G146), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(G113), .B(G122), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n219), .A2(new_n249), .A3(new_n234), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n234), .A2(new_n249), .ZN(new_n251));
  AOI21_X1  g065(.A(G146), .B1(new_n236), .B2(new_n238), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n239), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n229), .A2(new_n232), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(new_n246), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n188), .B1(new_n248), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT89), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n250), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n233), .A2(new_n261), .A3(new_n246), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n246), .B1(new_n233), .B2(new_n242), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n187), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT20), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n259), .B(new_n187), .C1(new_n262), .C2(new_n263), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT90), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n248), .A2(new_n257), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n259), .A4(new_n187), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n260), .A2(new_n266), .A3(new_n268), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n233), .A2(new_n261), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n247), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT91), .B1(new_n256), .B2(new_n246), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n262), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G475), .B1(new_n277), .B2(G902), .ZN(new_n278));
  AND2_X1   g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G214), .B1(G237), .B2(G902), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT82), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n208), .A2(G143), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n193), .B2(G146), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n284), .A2(KEYINPUT0), .A3(G128), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n208), .B1(new_n191), .B2(new_n192), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n196), .A2(G146), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT0), .B(G128), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G125), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT83), .ZN(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n296), .A3(KEYINPUT1), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n295), .A2(new_n297), .B1(new_n286), .B2(new_n287), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n223), .A2(new_n196), .ZN(new_n299));
  NAND2_X1  g113(.A1(KEYINPUT64), .A2(G143), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(G146), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n293), .A2(KEYINPUT1), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n282), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n206), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT83), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(G125), .C1(new_n285), .C2(new_n290), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n198), .A2(G224), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT7), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n292), .A2(new_n306), .A3(new_n308), .A4(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G122), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT8), .ZN(new_n314));
  INV_X1    g128(.A(G107), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n317));
  OAI211_X1 g131(.A(G104), .B(new_n315), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G101), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(G104), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n245), .A2(G107), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n318), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G101), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT67), .B1(new_n328), .B2(G116), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT67), .ZN(new_n330));
  INV_X1    g144(.A(G116), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(G119), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n329), .A2(new_n332), .B1(G116), .B2(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT5), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(G116), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(G113), .C1(KEYINPUT5), .C2(new_n335), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT2), .B(G113), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n327), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n327), .B1(new_n338), .B2(new_n336), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n314), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n318), .A2(new_n322), .A3(new_n321), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n323), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n333), .B(new_n337), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n346), .A3(G101), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n327), .A2(new_n336), .A3(new_n338), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n313), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n291), .A2(new_n306), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n310), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n312), .A2(new_n341), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n309), .B(KEYINPUT84), .Z(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n291), .A2(KEYINPUT83), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n308), .A2(new_n306), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n292), .A2(new_n306), .A3(new_n308), .A4(new_n356), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n348), .A2(new_n349), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n364));
  INV_X1    g178(.A(new_n313), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n365), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT6), .A3(new_n350), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n355), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G210), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n355), .A2(new_n369), .A3(new_n371), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n281), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G478), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT15), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n299), .A2(G128), .A3(new_n300), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n293), .A2(G143), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT92), .ZN(new_n382));
  INV_X1    g196(.A(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G116), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n331), .A2(G122), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n382), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(G107), .A3(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n384), .A2(new_n385), .A3(new_n382), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n315), .B1(new_n390), .B2(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n380), .B1(new_n378), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n191), .A2(new_n192), .A3(new_n293), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT93), .B1(new_n395), .B2(KEYINPUT13), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT93), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n378), .A2(new_n397), .A3(new_n393), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n381), .B(new_n392), .C1(new_n399), .C2(new_n379), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT14), .B1(new_n383), .B2(G116), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n383), .A2(G116), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT95), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(KEYINPUT14), .B2(new_n385), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n401), .A2(new_n402), .A3(KEYINPUT95), .ZN(new_n405));
  OAI21_X1  g219(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n378), .A2(new_n380), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G134), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n381), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT94), .B(new_n315), .C1(new_n390), .C2(new_n386), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n406), .A2(new_n409), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT9), .B(G234), .ZN(new_n414));
  INV_X1    g228(.A(G217), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n414), .A2(new_n415), .A3(G953), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n400), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT96), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n400), .A2(new_n413), .A3(new_n419), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n400), .A2(new_n413), .ZN(new_n421));
  INV_X1    g235(.A(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n354), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT97), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(new_n354), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n377), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n377), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n198), .A2(G952), .ZN(new_n434));
  INV_X1    g248(.A(G234), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n197), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n354), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n279), .A2(new_n375), .A3(new_n433), .A4(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G221), .ZN(new_n443));
  INV_X1    g257(.A(new_n414), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n354), .ZN(new_n445));
  AOI21_X1  g259(.A(G146), .B1(new_n299), .B2(new_n300), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT1), .ZN(new_n447));
  OAI21_X1  g261(.A(G128), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n301), .A2(new_n282), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n448), .A2(new_n449), .B1(new_n303), .B2(KEYINPUT78), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT78), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n284), .A2(new_n451), .A3(new_n302), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n326), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT10), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT68), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n298), .B2(new_n304), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(G128), .A3(new_n297), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n286), .A2(new_n287), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT68), .A3(new_n303), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n456), .A2(new_n461), .A3(new_n327), .A4(KEYINPUT10), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n285), .A2(new_n290), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n347), .A3(new_n344), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n454), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT11), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n379), .B2(G137), .ZN(new_n467));
  INV_X1    g281(.A(G137), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(KEYINPUT11), .A3(G134), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n379), .A2(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(KEYINPUT65), .A2(G131), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n473), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n454), .A2(new_n475), .A3(new_n462), .A4(new_n464), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G140), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n198), .A2(G227), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n478), .B(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n447), .B1(new_n221), .B2(new_n208), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n449), .B1(new_n483), .B2(new_n293), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n303), .A2(KEYINPUT78), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n452), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n327), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n305), .A2(new_n326), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n473), .A2(KEYINPUT12), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n482), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT79), .B(new_n490), .C1(new_n487), .C2(new_n488), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n326), .A2(new_n303), .A3(new_n460), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT80), .B1(new_n453), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT80), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(new_n497), .A3(new_n488), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n498), .A3(new_n473), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT12), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n494), .A2(new_n501), .A3(KEYINPUT81), .ZN(new_n502));
  INV_X1    g316(.A(new_n480), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n476), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT81), .B1(new_n494), .B2(new_n501), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n481), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G469), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n354), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n354), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n475), .B1(new_n489), .B2(KEYINPUT80), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT12), .B1(new_n511), .B2(new_n498), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n491), .B1(new_n453), .B2(new_n495), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT79), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n489), .A2(new_n482), .A3(new_n491), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n476), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n517), .A2(new_n480), .B1(new_n474), .B2(new_n504), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n510), .B1(new_n518), .B2(G469), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n445), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n442), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n468), .A2(G134), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(new_n470), .A3(G131), .ZN(new_n524));
  INV_X1    g338(.A(new_n471), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(G131), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n456), .A2(new_n461), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n345), .B1(new_n463), .B2(new_n473), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n456), .A2(new_n461), .A3(KEYINPUT69), .A4(new_n526), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n463), .A2(new_n473), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n526), .B1(new_n298), .B2(new_n304), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n529), .A2(new_n533), .A3(new_n531), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(KEYINPUT30), .ZN(new_n538));
  INV_X1    g352(.A(new_n345), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n541));
  NAND3_X1  g355(.A1(new_n197), .A2(new_n198), .A3(G210), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT28), .B1(new_n530), .B2(new_n527), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n533), .A2(new_n535), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n345), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n532), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI211_X1 g371(.A(KEYINPUT72), .B(new_n552), .C1(new_n532), .C2(new_n554), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n545), .B(KEYINPUT71), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n354), .B1(new_n549), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n546), .A2(new_n548), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n529), .A2(new_n531), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n563), .A2(new_n530), .B1(new_n537), .B2(new_n345), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n551), .B(new_n562), .C1(new_n564), .C2(new_n552), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n537), .A2(new_n345), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n532), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n550), .B1(new_n568), .B2(KEYINPUT28), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n562), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G472), .B1(new_n561), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(G472), .A2(G902), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT73), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n537), .A2(KEYINPUT30), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n345), .B1(new_n576), .B2(new_n536), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(KEYINPUT31), .A3(new_n532), .A4(new_n545), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n532), .B(new_n545), .C1(new_n538), .C2(new_n539), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n575), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT32), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT32), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n532), .A2(new_n554), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT72), .B1(new_n587), .B2(new_n552), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n555), .A2(new_n556), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(new_n551), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n581), .A2(new_n578), .B1(new_n590), .B2(new_n559), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n586), .B1(new_n591), .B2(new_n575), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n573), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n328), .B2(G128), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n293), .A2(KEYINPUT23), .A3(G119), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n596), .B(new_n597), .C1(G119), .C2(new_n293), .ZN(new_n598));
  XNOR2_X1  g412(.A(G119), .B(G128), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT24), .B(G110), .Z(new_n600));
  OAI22_X1  g414(.A1(new_n598), .A2(G110), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n239), .A3(new_n215), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n598), .A2(G110), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  INV_X1    g418(.A(new_n239), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n603), .B(new_n604), .C1(new_n252), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n254), .B2(new_n603), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n602), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT22), .B(G137), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n443), .A2(new_n435), .A3(G953), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n602), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n603), .B1(new_n605), .B2(new_n252), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(KEYINPUT75), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n616), .B2(new_n606), .ZN(new_n617));
  INV_X1    g431(.A(new_n612), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n613), .A2(new_n619), .A3(new_n354), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT25), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n613), .A2(new_n619), .A3(KEYINPUT25), .A4(new_n354), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n415), .B1(G234), .B2(new_n354), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n613), .A2(new_n619), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(G902), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n593), .A2(new_n594), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n594), .B1(new_n593), .B2(new_n632), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n522), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  AND2_X1   g450(.A1(new_n579), .A2(new_n580), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n579), .A2(new_n580), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n583), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n575), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(G902), .B1(new_n582), .B2(new_n583), .ZN(new_n642));
  INV_X1    g456(.A(G472), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n521), .A2(new_n644), .A3(new_n631), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n272), .A2(new_n278), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n354), .A2(G478), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n416), .B1(new_n400), .B2(new_n413), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI221_X4 g464(.A(new_n647), .B1(new_n650), .B2(new_n417), .C1(new_n424), .C2(new_n649), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n648), .B1(KEYINPUT96), .B2(new_n417), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n652), .B2(new_n420), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT98), .B1(new_n653), .B2(G478), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT98), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n425), .A2(new_n655), .A3(new_n376), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n280), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n373), .B2(new_n374), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n659), .A2(new_n440), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n645), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  OAI21_X1  g480(.A(new_n278), .B1(new_n429), .B2(new_n431), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n260), .A2(new_n266), .A3(new_n267), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT99), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT99), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n260), .A2(new_n670), .A3(new_n266), .A4(new_n267), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n441), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n662), .B1(new_n673), .B2(KEYINPUT100), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n675), .A3(new_n441), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n645), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n617), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n629), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n626), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n442), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n521), .A2(new_n644), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  AND3_X1   g504(.A1(new_n520), .A2(new_n661), .A3(new_n684), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n437), .B1(new_n438), .B2(new_n692), .ZN(new_n693));
  AOI211_X1 g507(.A(new_n693), .B(new_n667), .C1(new_n669), .C2(new_n671), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n593), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  INV_X1    g510(.A(new_n559), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT103), .B1(new_n564), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n568), .A2(new_n699), .A3(new_n559), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n579), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n643), .B1(new_n701), .B2(new_n354), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n585), .A2(new_n592), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n373), .A2(new_n374), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT102), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n280), .A3(new_n685), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n646), .A2(new_n432), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n705), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n693), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n520), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n714), .A2(KEYINPUT40), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n221), .ZN(G45));
  INV_X1    g532(.A(new_n693), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n646), .A2(new_n658), .A3(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n691), .A2(new_n593), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND2_X1  g537(.A1(new_n507), .A2(new_n354), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n509), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n445), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n663), .A2(new_n593), .A3(new_n727), .A4(new_n632), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  NAND2_X1  g544(.A1(new_n566), .A2(new_n571), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT29), .B1(new_n540), .B2(new_n546), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n590), .B2(new_n559), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n733), .A3(new_n354), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n734), .A2(G472), .B1(new_n584), .B2(KEYINPUT32), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n631), .B1(new_n735), .B2(new_n592), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n674), .A2(new_n736), .A3(new_n676), .A4(new_n727), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  INV_X1    g552(.A(new_n445), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n739), .A3(new_n509), .A4(new_n661), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n508), .B1(new_n507), .B2(new_n354), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT81), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n512), .B2(new_n516), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n504), .A3(new_n502), .ZN(new_n746));
  AOI211_X1 g560(.A(G469), .B(G902), .C1(new_n746), .C2(new_n481), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT104), .A3(new_n739), .A4(new_n661), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n646), .A2(new_n432), .A3(new_n685), .A4(new_n440), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n742), .A2(new_n749), .A3(new_n593), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G119), .ZN(G21));
  NOR3_X1   g566(.A1(new_n740), .A2(new_n440), .A3(new_n711), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n569), .A2(new_n697), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n575), .B1(new_n582), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n639), .A2(new_n354), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n631), .B(new_n755), .C1(G472), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  AND2_X1   g573(.A1(new_n742), .A2(new_n749), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n720), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n579), .B(KEYINPUT31), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n569), .A2(new_n697), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n640), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n765), .B(new_n684), .C1(new_n642), .C2(new_n643), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n657), .B1(new_n272), .B2(new_n278), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT105), .B1(new_n767), .B2(new_n719), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n762), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n760), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n742), .A2(new_n749), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n720), .A2(new_n761), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n755), .B1(new_n756), .B2(G472), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n767), .A2(KEYINPUT105), .A3(new_n719), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n684), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT106), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n592), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n641), .A2(KEYINPUT107), .A3(new_n586), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n735), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n632), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n373), .A2(new_n374), .A3(new_n280), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n445), .B(new_n785), .C1(new_n509), .C2(new_n519), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n773), .A3(new_n775), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT42), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n762), .A2(new_n768), .A3(KEYINPUT42), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n736), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n218), .ZN(G33));
  NAND4_X1  g606(.A1(new_n736), .A2(KEYINPUT108), .A3(new_n694), .A4(new_n786), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n593), .A2(new_n694), .A3(new_n786), .A4(new_n632), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT108), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NAND2_X1  g612(.A1(new_n644), .A2(new_n684), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT109), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n279), .A2(new_n658), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT43), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT44), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n518), .A2(KEYINPUT45), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n508), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n518), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n510), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT46), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n747), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  INV_X1    g627(.A(new_n785), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n739), .A3(new_n713), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n804), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n800), .A2(KEYINPUT44), .A3(new_n803), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  OR4_X1    g633(.A1(new_n593), .A2(new_n632), .A3(new_n720), .A4(new_n785), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n813), .A2(new_n739), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n813), .A2(KEYINPUT47), .A3(new_n739), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n820), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT110), .B(G140), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(G42));
  XNOR2_X1  g641(.A(new_n726), .B(KEYINPUT111), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT49), .Z(new_n829));
  OR3_X1    g643(.A1(new_n631), .A2(new_n445), .A3(new_n281), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n830), .A2(new_n709), .A3(new_n801), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n705), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n803), .A2(new_n437), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n726), .A2(new_n445), .A3(new_n785), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n684), .A3(new_n774), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n705), .A2(new_n834), .A3(new_n632), .A4(new_n437), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n836), .A2(new_n646), .A3(new_n658), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n709), .A2(new_n280), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n727), .A2(new_n833), .A3(new_n757), .A4(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n840));
  OAI211_X1 g654(.A(new_n835), .B(new_n837), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(KEYINPUT50), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n843), .B2(new_n839), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n833), .A2(new_n757), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n823), .A2(new_n824), .ZN(new_n846));
  INV_X1    g660(.A(new_n828), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n445), .B1(new_n847), .B2(KEYINPUT117), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(KEYINPUT117), .B2(new_n847), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n814), .B(new_n845), .C1(new_n846), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n844), .A2(KEYINPUT51), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n760), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n434), .C1(new_n659), .C2(new_n836), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n833), .A2(new_n632), .A3(new_n783), .A4(new_n834), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n770), .B1(new_n760), .B2(new_n769), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n772), .A2(new_n776), .A3(KEYINPUT106), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n695), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n695), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n771), .B2(new_n777), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT112), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n684), .A2(new_n693), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n517), .A2(new_n480), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n504), .A2(new_n474), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n871), .A2(G469), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n809), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n870), .B(new_n739), .C1(new_n747), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT113), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n646), .A2(new_n432), .A3(new_n661), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n509), .A2(new_n519), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(new_n880), .A3(new_n739), .A4(new_n870), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n876), .A2(new_n704), .A3(new_n878), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n702), .B1(new_n641), .B2(new_n586), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n877), .B1(new_n885), .B2(new_n585), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(KEYINPUT114), .A3(new_n876), .A4(new_n881), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n887), .A3(new_n722), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n866), .A2(new_n869), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n864), .B2(new_n888), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n758), .A2(new_n751), .A3(new_n728), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n375), .A2(new_n441), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n279), .A2(new_n432), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n659), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n645), .A2(new_n898), .B1(new_n686), .B2(new_n687), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n635), .A3(new_n737), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n669), .A2(new_n671), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n685), .A2(new_n693), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n278), .A4(new_n433), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n592), .B2(new_n735), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n786), .B1(new_n769), .B2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n797), .A2(new_n788), .A3(new_n905), .A4(new_n790), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n893), .A2(new_n894), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n884), .A2(new_n887), .A3(new_n722), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(new_n868), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT53), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n908), .A2(KEYINPUT54), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT115), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n635), .A2(new_n899), .A3(KEYINPUT53), .ZN(new_n916));
  INV_X1    g730(.A(new_n737), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n758), .A2(new_n751), .A3(new_n728), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT116), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n895), .A2(new_n920), .A3(new_n737), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(new_n906), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n893), .A2(new_n923), .B1(new_n912), .B2(new_n894), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(new_n914), .A3(KEYINPUT115), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n861), .B1(new_n915), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(G952), .A2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n832), .B1(new_n928), .B2(new_n929), .ZN(G75));
  NOR2_X1   g744(.A1(new_n198), .A2(G952), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n868), .A2(KEYINPUT112), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n865), .B(new_n867), .C1(new_n771), .C2(new_n777), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n909), .A2(KEYINPUT52), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n923), .B1(new_n935), .B2(new_n911), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n912), .A2(new_n894), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n938), .A2(G210), .A3(G902), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT56), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n368), .A2(new_n366), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(new_n362), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n931), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT120), .B1(new_n924), .B2(new_n354), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  INV_X1    g761(.A(new_n906), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(new_n919), .A3(new_n921), .A4(new_n916), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n892), .B2(new_n891), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n909), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n892), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT53), .B1(new_n952), .B2(new_n907), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n947), .B(G902), .C1(new_n950), .C2(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n946), .A2(new_n372), .A3(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n944), .A2(KEYINPUT56), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n945), .A2(new_n957), .ZN(G51));
  XNOR2_X1  g772(.A(new_n510), .B(KEYINPUT57), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT54), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n925), .B1(new_n936), .B2(new_n937), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n507), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n946), .A2(new_n807), .A3(new_n806), .A4(new_n954), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n931), .B1(new_n963), .B2(new_n964), .ZN(G54));
  AND2_X1   g779(.A1(KEYINPUT58), .A2(G475), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n946), .A2(new_n954), .A3(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n269), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n931), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n946), .A2(new_n269), .A3(new_n954), .A4(new_n966), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G60));
  NAND2_X1  g786(.A1(new_n424), .A2(new_n649), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n650), .A2(new_n417), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n376), .A2(new_n354), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(new_n978));
  NOR2_X1   g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n960), .B2(new_n961), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n970), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n915), .A2(new_n927), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n983), .B2(new_n975), .ZN(G63));
  INV_X1    g798(.A(KEYINPUT61), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n987));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n936), .B2(new_n937), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n970), .B1(new_n990), .B2(new_n628), .ZN(new_n991));
  INV_X1    g805(.A(new_n989), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n938), .A2(new_n682), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n986), .B(new_n987), .C1(new_n991), .C2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n950), .B2(new_n953), .ZN(new_n995));
  INV_X1    g809(.A(new_n628), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n931), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n990), .A2(new_n682), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n997), .A2(KEYINPUT122), .A3(new_n985), .A4(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n994), .A2(new_n999), .ZN(G66));
  INV_X1    g814(.A(G224), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n439), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n900), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n942), .B1(G898), .B2(new_n198), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1004), .B(new_n1006), .ZN(G69));
  XNOR2_X1  g821(.A(new_n538), .B(KEYINPUT124), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n241), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n932), .A2(new_n933), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n717), .A3(new_n722), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1011), .A2(new_n1014), .A3(new_n717), .A4(new_n722), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n785), .B(new_n714), .C1(new_n659), .C2(new_n897), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1016), .B1(new_n634), .B2(new_n633), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT125), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n825), .B1(new_n816), .B2(new_n817), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1010), .B1(new_n1020), .B2(new_n198), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n791), .B1(new_n796), .B2(new_n793), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n784), .A2(new_n877), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1023), .A2(new_n739), .A3(new_n713), .A4(new_n813), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1019), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1011), .A2(new_n722), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n198), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n692), .A2(G953), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT126), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1009), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1032), .B1(new_n1021), .B2(new_n1030), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(new_n540), .A2(new_n545), .ZN(new_n1037));
  OR2_X1    g851(.A1(new_n1020), .A2(new_n900), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G472), .A2(G902), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT63), .Z(new_n1040));
  AOI21_X1  g854(.A(new_n1037), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g855(.A(new_n1040), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1042), .B1(new_n547), .B2(new_n579), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n908), .A2(new_n913), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1042), .B1(new_n1045), .B2(new_n1003), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n577), .A2(new_n532), .A3(new_n546), .ZN(new_n1047));
  OAI211_X1 g861(.A(new_n970), .B(new_n1044), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1041), .A2(new_n1048), .ZN(G57));
endmodule


