//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G236), .A2(G238), .A3(G237), .A4(G235), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OAI211_X1 g038(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n454), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT68), .Z(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n469), .B2(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(G101), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n466), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n482), .B(new_n466), .C1(new_n478), .C2(new_n479), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n475), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n470), .A2(new_n472), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT72), .Z(new_n490));
  INV_X1    g065(.A(G112), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n469), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AOI22_X1  g067(.A1(new_n488), .A2(G124), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n486), .A2(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .A3(G136), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT71), .B1(new_n495), .B2(G136), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT73), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G162));
  INV_X1    g078(.A(G126), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n470), .B2(new_n472), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n506), .B2(new_n469), .ZN(new_n507));
  OAI21_X1  g082(.A(G2105), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT4), .A2(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n470), .B2(new_n472), .ZN(new_n510));
  AND2_X1   g085(.A1(G102), .A2(G2104), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n466), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT3), .B(G2104), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G138), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G164));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT74), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .A3(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT75), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n519), .A2(KEYINPUT6), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT6), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G651), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G50), .ZN(new_n534));
  INV_X1    g109(.A(G88), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n521), .A2(new_n523), .A3(new_n529), .A4(new_n531), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n528), .A2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n529), .A2(new_n531), .A3(G51), .A4(G543), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n521), .A2(new_n523), .A3(G63), .A4(G651), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G168));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n533), .A2(new_n547), .B1(new_n548), .B2(new_n536), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n521), .A2(new_n523), .A3(G64), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n519), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n533), .A2(new_n554), .B1(new_n555), .B2(new_n536), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n521), .A2(new_n523), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n556), .B1(KEYINPUT76), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n561), .A2(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND4_X1  g145(.A1(new_n529), .A2(new_n531), .A3(G53), .A4(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n558), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  INV_X1    g151(.A(new_n536), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G91), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n576), .A3(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  OR3_X1    g155(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT77), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n543), .B2(new_n545), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G286));
  OR2_X1    g158(.A1(new_n528), .A2(new_n537), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n532), .A2(G49), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n536), .ZN(G288));
  NAND3_X1  g163(.A1(new_n521), .A2(new_n523), .A3(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n524), .A2(G86), .A3(new_n532), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n529), .A2(new_n531), .A3(G48), .A4(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n558), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n532), .A2(G543), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G47), .B1(new_n577), .B2(G85), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n599), .A2(KEYINPUT78), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n558), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n601), .A2(G54), .B1(new_n610), .B2(G651), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n536), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(KEYINPUT10), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G284));
  OAI21_X1  g193(.A(new_n607), .B1(new_n617), .B2(G868), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(KEYINPUT79), .B1(new_n621), .B2(G299), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT79), .B2(new_n620), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(KEYINPUT79), .B2(new_n620), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n617), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n617), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n488), .A2(G123), .ZN(new_n633));
  AND2_X1   g208(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n495), .A2(G135), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  OR3_X1    g213(.A1(new_n636), .A2(KEYINPUT84), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(KEYINPUT84), .B1(new_n636), .B2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n469), .A2(G2105), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n513), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT13), .ZN(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT81), .Z(new_n649));
  INV_X1    g224(.A(G2096), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n639), .A2(new_n650), .A3(new_n640), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n646), .A2(new_n647), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT80), .ZN(new_n653));
  NAND4_X1  g228(.A1(new_n642), .A2(new_n649), .A3(new_n651), .A4(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2427), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2430), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  AND3_X1   g240(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT14), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n660), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(G401));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  NOR2_X1   g247(.A1(G2072), .A2(G2078), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n444), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n674), .B(KEYINPUT17), .Z(new_n679));
  OAI211_X1 g254(.A(new_n672), .B(new_n678), .C1(new_n679), .C2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT87), .ZN(new_n681));
  INV_X1    g256(.A(new_n672), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n682), .A3(new_n677), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT88), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n672), .A2(new_n677), .A3(new_n675), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT18), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(new_n650), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G2100), .ZN(G227));
  XNOR2_X1  g264(.A(G1956), .B(G2474), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1961), .B(G1966), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1971), .B(G1976), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT19), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n693), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT20), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n690), .A2(new_n691), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n696), .B2(new_n692), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(KEYINPUT90), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT92), .Z(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n705), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(KEYINPUT102), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT97), .ZN(new_n715));
  NAND2_X1  g290(.A1(G288), .A2(G16), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT33), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G23), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n717), .B1(new_n716), .B2(new_n719), .ZN(new_n722));
  OAI21_X1  g297(.A(G1976), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1976), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n725), .A3(new_n720), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(G303), .A2(G16), .ZN(new_n729));
  INV_X1    g304(.A(G1971), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n718), .A2(G22), .ZN(new_n731));
  AND3_X1   g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(G305), .A2(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n718), .A2(G6), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT32), .B(G1981), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n740), .A2(KEYINPUT96), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n734), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n715), .B1(new_n728), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT96), .B1(new_n740), .B2(new_n741), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n748), .A2(new_n732), .A3(new_n733), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n749), .A2(KEYINPUT97), .A3(new_n727), .A4(new_n742), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(KEYINPUT34), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n718), .A2(G24), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n605), .B2(new_n718), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT95), .B(G1986), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT35), .B(G1991), .Z(new_n756));
  OR2_X1    g331(.A1(G95), .A2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(G107), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n469), .B1(new_n758), .B2(G2105), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n488), .A2(G119), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n495), .A2(G131), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n762), .A2(new_n763), .ZN(new_n766));
  OAI21_X1  g341(.A(G29), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G25), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n767), .A2(KEYINPUT94), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(KEYINPUT94), .B1(new_n767), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n756), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(new_n756), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n774), .A2(new_n775), .A3(new_n770), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n755), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n751), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(KEYINPUT34), .B1(new_n747), .B2(new_n750), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT36), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n779), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n781), .A2(new_n782), .A3(new_n751), .A4(new_n777), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n768), .A2(G35), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT100), .Z(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n502), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  OAI21_X1  g367(.A(G2090), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(KEYINPUT101), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT101), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n795), .B(G2090), .C1(new_n791), .C2(new_n792), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n768), .A2(G26), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT28), .Z(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(new_n466), .B2(G116), .ZN(new_n800));
  INV_X1    g375(.A(G104), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n466), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n488), .B2(G128), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n495), .A2(new_n804), .A3(G140), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n804), .B1(new_n495), .B2(G140), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n799), .B1(new_n807), .B2(G29), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n808), .A2(G2067), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(G2067), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n641), .A2(new_n768), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G5), .A2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT99), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G171), .B2(G16), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G1961), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT25), .Z(new_n818));
  INV_X1    g393(.A(G139), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n513), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n820));
  OAI221_X1 g395(.A(new_n818), .B1(new_n819), .B2(new_n494), .C1(new_n466), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n768), .A2(G33), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n816), .B1(G2072), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT26), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(G105), .B2(new_n643), .ZN(new_n830));
  INV_X1    g405(.A(G141), .ZN(new_n831));
  INV_X1    g406(.A(G129), .ZN(new_n832));
  OAI221_X1 g407(.A(new_n830), .B1(new_n494), .B2(new_n831), .C1(new_n832), .C2(new_n487), .ZN(new_n833));
  MUX2_X1   g408(.A(G32), .B(new_n833), .S(G29), .Z(new_n834));
  XOR2_X1   g409(.A(KEYINPUT27), .B(G1996), .Z(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n718), .A2(G21), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G168), .B2(new_n718), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(G1966), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n834), .B2(new_n835), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n815), .A2(G1961), .B1(G1966), .B2(new_n838), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n825), .A2(new_n836), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n811), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n718), .A2(G19), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(new_n564), .B2(G16), .ZN(new_n845));
  INV_X1    g420(.A(G1341), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n718), .A2(G20), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT23), .Z(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G299), .B2(G16), .ZN(new_n851));
  INV_X1    g426(.A(G1956), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n847), .A2(new_n848), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G164), .A2(G29), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(G27), .B2(G29), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(new_n443), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n443), .ZN(new_n858));
  INV_X1    g433(.A(G2084), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n768), .B1(KEYINPUT24), .B2(G34), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n860), .B1(KEYINPUT24), .B2(G34), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n484), .B2(G29), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT30), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(G28), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n768), .B1(new_n864), .B2(G28), .ZN(new_n866));
  AND2_X1   g441(.A1(KEYINPUT31), .A2(G11), .ZN(new_n867));
  NOR2_X1   g442(.A1(KEYINPUT31), .A2(G11), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n824), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n442), .ZN(new_n871));
  INV_X1    g446(.A(G1348), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n718), .A2(G4), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n872), .B(new_n873), .C1(new_n617), .C2(new_n718), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n617), .B2(new_n718), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G1348), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n862), .A2(new_n859), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n871), .A2(new_n874), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n863), .A2(new_n878), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n843), .A2(new_n854), .A3(new_n879), .ZN(new_n880));
  OR3_X1    g455(.A1(new_n791), .A2(G2090), .A3(new_n792), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n797), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n714), .B1(new_n784), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g459(.A(KEYINPUT102), .B(new_n882), .C1(new_n780), .C2(new_n783), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(G311));
  AOI21_X1  g461(.A(KEYINPUT103), .B1(new_n784), .B2(new_n883), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  AOI211_X1 g463(.A(new_n888), .B(new_n882), .C1(new_n780), .C2(new_n783), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(G150));
  AOI22_X1  g465(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n891), .A2(new_n519), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n524), .A2(G93), .A3(new_n532), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n532), .A2(G55), .A3(G543), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n894), .B1(new_n893), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n564), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n896), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n902), .A2(new_n562), .A3(new_n563), .A4(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT38), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n617), .A2(G559), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g483(.A(G860), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n908), .B2(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n899), .A2(G860), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT37), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G145));
  XNOR2_X1  g488(.A(new_n502), .B(new_n484), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(new_n641), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n762), .B(new_n833), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n495), .A2(G142), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n488), .A2(G130), .ZN(new_n919));
  OAI21_X1  g494(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n466), .A2(G118), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n922), .B2(new_n921), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n918), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(new_n645), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n807), .B(new_n517), .ZN(new_n927));
  INV_X1    g502(.A(new_n821), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n929), .A2(new_n930), .A3(new_n926), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n917), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n932), .A2(new_n917), .A3(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n915), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  INV_X1    g513(.A(new_n915), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(new_n934), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g518(.A(G305), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n605), .B(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(G166), .B(G288), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n945), .B(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT109), .B1(new_n948), .B2(KEYINPUT108), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  XOR2_X1   g529(.A(new_n904), .B(new_n627), .Z(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  INV_X1    g531(.A(G299), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n616), .ZN(new_n958));
  OAI211_X1 g533(.A(G299), .B(new_n611), .C1(new_n615), .C2(new_n614), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT107), .A4(KEYINPUT41), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT106), .B1(new_n957), .B2(new_n616), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n960), .B2(KEYINPUT106), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n962), .B(new_n963), .C1(new_n965), .C2(KEYINPUT41), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n955), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n960), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n955), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n949), .A2(new_n970), .A3(new_n952), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n954), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n969), .B1(new_n954), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(G868), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n899), .A2(new_n621), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(G295));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n975), .ZN(G331));
  XNOR2_X1  g552(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n581), .A2(G171), .A3(new_n582), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n581), .A2(G171), .A3(KEYINPUT111), .A4(new_n582), .ZN(new_n983));
  NAND2_X1  g558(.A1(G301), .A2(G168), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n900), .A3(new_n903), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n980), .A2(new_n981), .B1(G168), .B2(G301), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n904), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n968), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n985), .B(new_n904), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n966), .ZN(new_n991));
  AOI21_X1  g566(.A(G37), .B1(new_n991), .B2(new_n948), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n947), .B(new_n989), .C1(new_n966), .C2(new_n990), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n979), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n968), .B1(new_n990), .B2(new_n961), .ZN(new_n996));
  INV_X1    g571(.A(new_n986), .ZN(new_n997));
  INV_X1    g572(.A(new_n988), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT41), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n996), .B(new_n947), .C1(new_n965), .C2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n992), .ZN(new_n1001));
  OAI22_X1  g576(.A1(new_n994), .A2(new_n995), .B1(new_n1001), .B2(KEYINPUT43), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT112), .B(new_n979), .C1(new_n992), .C2(new_n993), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n978), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n1001), .B2(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n992), .A2(new_n979), .A3(new_n993), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1004), .B1(new_n1009), .B2(new_n1010), .ZN(G397));
  INV_X1    g586(.A(G1384), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n517), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(G40), .B(new_n475), .C1(new_n481), .C2(new_n483), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n1018), .A2(new_n1019), .A3(G1996), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n807), .B(G2067), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1021), .B2(new_n833), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1018), .B2(G1996), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT47), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1017), .A2(G1996), .A3(new_n833), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n833), .A2(G1996), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1017), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n762), .B(new_n775), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1017), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT48), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1025), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n765), .A2(new_n775), .A3(new_n766), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1033), .A2(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n807), .A2(G2067), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1018), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  NAND3_X1  g621(.A1(G303), .A2(new_n1046), .A3(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT55), .B1(G166), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1047), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1014), .A2(G1384), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n517), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT116), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1016), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n517), .A2(new_n1058), .A3(new_n1054), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1056), .A2(new_n1015), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n730), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1063), .B1(new_n517), .B2(new_n1012), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2090), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n517), .A2(new_n1012), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1065), .A2(new_n1066), .A3(new_n1057), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1060), .B2(new_n730), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n1053), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1981), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n592), .A2(new_n1073), .A3(new_n593), .A4(new_n594), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n1075));
  INV_X1    g650(.A(G86), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n594), .B1(new_n536), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n519), .B1(new_n589), .B2(new_n590), .ZN(new_n1078));
  OAI21_X1  g653(.A(G1981), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1075), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G305), .A2(KEYINPUT120), .A3(G1981), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT49), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT49), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1080), .A2(new_n1086), .A3(new_n1081), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G288), .A2(new_n725), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT52), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1089), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n725), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1091), .A2(G8), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(KEYINPUT63), .A3(new_n1090), .A4(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1057), .A2(new_n1055), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT45), .B1(new_n517), .B2(new_n1012), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT121), .B(G2084), .Z(new_n1100));
  NAND4_X1  g675(.A1(new_n1065), .A2(new_n1057), .A3(new_n1068), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G286), .A2(new_n1049), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1095), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1072), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1060), .A2(new_n730), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT117), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n1069), .A3(new_n1062), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1109), .A2(G8), .B1(new_n1050), .B2(new_n1047), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1045), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1088), .A2(new_n1090), .A3(new_n1094), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1067), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1013), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n517), .A2(new_n1063), .A3(new_n1012), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1115), .A2(new_n1057), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1066), .A2(new_n1117), .B1(new_n1060), .B2(new_n730), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1113), .B1(new_n1118), .B2(new_n1049), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1104), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1072), .A2(new_n1112), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT63), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1113), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(KEYINPUT122), .A3(new_n1072), .A4(new_n1105), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1111), .A2(new_n1123), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1099), .A2(G168), .A3(new_n1101), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(G168), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1132), .A3(G8), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT62), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1060), .B2(G2078), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(G2078), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1015), .A2(new_n1057), .A3(new_n1055), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1057), .A2(new_n1068), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n1141), .B2(new_n1064), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1065), .A2(new_n1143), .A3(new_n1057), .A4(new_n1068), .ZN(new_n1144));
  AOI21_X1  g719(.A(G1961), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(G171), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1072), .A2(new_n1112), .A3(new_n1119), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1131), .A2(new_n1149), .A3(new_n1133), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1135), .A2(new_n1147), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(G288), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1088), .A2(new_n725), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1084), .B1(new_n1153), .B2(new_n1074), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1072), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1155), .B2(new_n1112), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1127), .A2(new_n1151), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1158));
  INV_X1    g733(.A(G1961), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(G40), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n480), .B2(G2105), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT125), .A3(new_n475), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1138), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT125), .B1(new_n1162), .B2(new_n475), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1166), .A2(new_n1056), .A3(new_n1015), .A4(new_n1059), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n517), .A2(new_n1054), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1098), .B1(new_n1058), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1171), .A2(KEYINPUT126), .A3(new_n1056), .A4(new_n1166), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1160), .A2(new_n1173), .A3(G301), .A4(new_n1137), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1146), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT54), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1160), .A2(new_n1173), .A3(new_n1137), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(G171), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1171), .A2(new_n443), .A3(new_n1057), .A4(new_n1056), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n1158), .A2(new_n1159), .B1(new_n1180), .B2(new_n1136), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1139), .A2(G301), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1176), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1179), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1177), .A2(new_n1148), .A3(new_n1184), .A4(new_n1134), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n1188));
  AOI21_X1  g763(.A(G1348), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1091), .A2(G2067), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1158), .B2(new_n872), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n616), .B1(new_n1192), .B2(KEYINPUT60), .ZN(new_n1193));
  NOR4_X1   g768(.A1(new_n1189), .A2(new_n1188), .A3(new_n617), .A4(new_n1190), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1191), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(KEYINPUT58), .B(G1341), .Z(new_n1196));
  NAND2_X1  g771(.A1(new_n1091), .A2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(new_n1060), .B2(G1996), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n565), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(KEYINPUT123), .A2(KEYINPUT57), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT57), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OR3_X1    g782(.A1(G299), .A2(new_n1204), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g783(.A1(G299), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  XOR2_X1   g785(.A(KEYINPUT56), .B(G2072), .Z(new_n1211));
  NOR2_X1   g786(.A1(new_n1060), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1016), .B1(new_n1013), .B2(new_n1114), .ZN(new_n1213));
  AOI21_X1  g788(.A(G1956), .B1(new_n1213), .B2(new_n1116), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1210), .B1(new_n1212), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1213), .A2(new_n1116), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n852), .ZN(new_n1217));
  INV_X1    g792(.A(new_n1210), .ZN(new_n1218));
  OAI211_X1 g793(.A(new_n1217), .B(new_n1218), .C1(new_n1060), .C2(new_n1211), .ZN(new_n1219));
  AOI21_X1  g794(.A(KEYINPUT61), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1203), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1215), .A2(new_n1219), .A3(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1195), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g798(.A(new_n1215), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1219), .A2(new_n617), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1192), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g802(.A1(new_n1185), .A2(new_n1186), .B1(new_n1223), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1157), .B1(new_n1187), .B2(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n605), .B(G1986), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1033), .B(new_n1035), .C1(new_n1018), .C2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1044), .B1(new_n1229), .B2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g807(.A1(new_n669), .A2(new_n464), .ZN(new_n1234));
  NOR3_X1   g808(.A1(G227), .A2(G229), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g809(.A(new_n942), .B(new_n1235), .C1(new_n1002), .C2(new_n1003), .ZN(G225));
  INV_X1    g810(.A(G225), .ZN(G308));
endmodule


