//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT91), .ZN(new_n211));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(KEYINPUT15), .B2(new_n212), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  INV_X1    g015(.A(G36gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(KEYINPUT15), .A3(new_n212), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(new_n215), .B2(new_n219), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n207), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  XOR2_X1   g024(.A(new_n225), .B(KEYINPUT92), .Z(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n206), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n224), .A2(KEYINPUT18), .A3(new_n227), .A4(new_n228), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n220), .B(new_n206), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n226), .B(KEYINPUT93), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT13), .Z(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n231), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT11), .ZN(new_n239));
  INV_X1    g038(.A(G169gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT12), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n231), .A2(new_n243), .A3(new_n232), .A4(new_n236), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT36), .ZN(new_n249));
  NAND2_X1  g048(.A1(G227gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT28), .ZN(new_n252));
  INV_X1    g051(.A(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT65), .A2(G183gat), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT27), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT27), .B(G183gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n252), .B1(new_n261), .B2(new_n253), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT66), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n253), .B1(new_n265), .B2(new_n258), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT65), .B(G183gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n258), .B1(new_n268), .B2(KEYINPUT27), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n264), .B(new_n267), .C1(new_n269), .C2(new_n254), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n240), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n275), .A2(new_n278), .B1(G183gat), .B2(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n270), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n268), .B2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n277), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT64), .B1(new_n274), .B2(KEYINPUT23), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n271), .B1(new_n277), .B2(new_n288), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n290), .B2(new_n289), .ZN(new_n295));
  INV_X1    g094(.A(G183gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n253), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT25), .B1(new_n285), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n294), .A2(KEYINPUT25), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G113gat), .ZN(new_n300));
  INV_X1    g099(.A(G120gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT1), .ZN(new_n303));
  NAND2_X1  g102(.A1(G113gat), .A2(G120gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G127gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G134gat), .ZN(new_n308));
  INV_X1    g107(.A(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G127gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT68), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT68), .B1(new_n308), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n306), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n309), .ZN(new_n315));
  NAND2_X1  g114(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(G127gat), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n305), .A2(new_n317), .A3(new_n308), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(KEYINPUT69), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT68), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n309), .A2(G127gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n307), .A2(G134gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT68), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n305), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n305), .A2(new_n317), .A3(new_n308), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n320), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n280), .A2(new_n299), .A3(new_n319), .A4(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n280), .A2(new_n299), .B1(new_n319), .B2(new_n328), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n280), .A2(new_n299), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n328), .A2(new_n319), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n333), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n251), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  INV_X1    g139(.A(G71gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT71), .B(G99gat), .Z(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND3_X1  g143(.A1(new_n337), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n344), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n336), .B(KEYINPUT32), .C1(new_n338), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n334), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT70), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n331), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n251), .A2(KEYINPUT34), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n329), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n332), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n356), .A2(KEYINPUT73), .A3(new_n351), .A4(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n350), .A2(new_n250), .A3(new_n351), .A4(new_n329), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT34), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n359), .A2(KEYINPUT72), .A3(KEYINPUT34), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT72), .B1(new_n359), .B2(KEYINPUT34), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n368), .A2(new_n358), .B1(new_n345), .B2(new_n347), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n249), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n364), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n368), .A2(new_n347), .A3(new_n345), .A4(new_n358), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(KEYINPUT36), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  AND2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT81), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G155gat), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n382));
  NAND2_X1  g181(.A1(G155gat), .A2(G162gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G141gat), .B(G148gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT2), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(G155gat), .B2(G162gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT80), .B(KEYINPUT2), .ZN(new_n391));
  NAND2_X1  g190(.A1(G141gat), .A2(G148gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G141gat), .ZN(new_n396));
  INV_X1    g195(.A(G148gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n392), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n391), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT78), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT78), .B1(new_n379), .B2(new_n380), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n383), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n390), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n406), .A2(KEYINPUT74), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(KEYINPUT74), .ZN(new_n408));
  XNOR2_X1  g207(.A(G197gat), .B(G204gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G211gat), .B(G218gat), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n407), .A2(new_n411), .A3(new_n408), .A4(new_n409), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT29), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n405), .B1(new_n415), .B2(KEYINPUT3), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n375), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n391), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT79), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n399), .B1(new_n398), .B2(new_n392), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n404), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n422), .A2(new_n423), .B1(new_n385), .B2(new_n389), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT29), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n413), .A2(new_n414), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n416), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  OAI221_X1 g228(.A(new_n416), .B1(new_n417), .B2(new_n375), .C1(new_n426), .C2(new_n427), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(G22gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n430), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT86), .B(G22gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n431), .B(new_n434), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n429), .B2(new_n430), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT87), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n435), .A2(new_n436), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n443), .A2(new_n441), .ZN(new_n444));
  OAI22_X1  g243(.A1(new_n439), .A2(new_n442), .B1(new_n444), .B2(new_n434), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT5), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n313), .A2(new_n318), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n424), .B2(new_n425), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n395), .A2(new_n400), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n404), .B1(new_n452), .B2(new_n419), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n388), .B(new_n386), .C1(new_n378), .C2(new_n384), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT3), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n449), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n328), .A2(new_n424), .A3(new_n457), .A4(new_n319), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n424), .B2(new_n450), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n326), .A2(new_n327), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n405), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n463), .A2(KEYINPUT82), .A3(new_n457), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n456), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n405), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n422), .A2(new_n423), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n467), .A3(new_n390), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n447), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n448), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n390), .B(new_n425), .C1(new_n401), .C2(new_n404), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n462), .A3(new_n472), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n328), .A2(new_n424), .A3(KEYINPUT4), .A4(new_n319), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n405), .A2(new_n462), .B1(new_n457), .B2(new_n470), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n465), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G1gat), .B(G29gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT0), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(G57gat), .ZN(new_n481));
  INV_X1    g280(.A(G85gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n465), .A2(new_n477), .A3(new_n483), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT83), .B1(new_n488), .B2(new_n486), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT84), .B1(new_n478), .B2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n491), .B(new_n483), .C1(new_n465), .C2(new_n477), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n488), .A2(KEYINPUT83), .A3(new_n486), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n427), .ZN(new_n496));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n333), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n280), .B2(new_n299), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n333), .A2(new_n498), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT29), .B1(new_n280), .B2(new_n299), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n503), .B(new_n427), .C1(new_n498), .C2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G64gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(G92gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n502), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n502), .A2(new_n505), .A3(KEYINPUT76), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n502), .A2(new_n505), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n508), .ZN(new_n518));
  INV_X1    g317(.A(new_n508), .ZN(new_n519));
  AOI211_X1 g318(.A(KEYINPUT75), .B(new_n519), .C1(new_n502), .C2(new_n505), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n502), .A2(new_n505), .A3(new_n519), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n521), .A2(KEYINPUT77), .A3(new_n509), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT77), .B1(new_n521), .B2(new_n509), .ZN(new_n523));
  OAI221_X1 g322(.A(new_n515), .B1(new_n518), .B2(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n446), .B1(new_n495), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n374), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n374), .A2(KEYINPUT88), .A3(new_n525), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT82), .B1(new_n463), .B2(new_n457), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n459), .A2(new_n460), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n458), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n447), .B1(new_n533), .B2(new_n473), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT39), .B1(new_n469), .B2(new_n470), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n483), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g335(.A(KEYINPUT39), .B(new_n447), .C1(new_n533), .C2(new_n473), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n533), .A2(new_n456), .B1(new_n471), .B2(new_n476), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(new_n483), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n536), .A2(new_n537), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT40), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n544));
  NAND3_X1  g343(.A1(new_n502), .A2(new_n505), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n508), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n502), .B2(new_n505), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n546), .A2(KEYINPUT38), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n521), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT6), .B1(new_n539), .B2(new_n483), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n485), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n487), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(KEYINPUT89), .A3(new_n485), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT38), .B1(new_n546), .B2(new_n548), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n551), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n558), .A3(new_n445), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n528), .A2(new_n529), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n365), .A2(new_n369), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n515), .B1(new_n518), .B2(new_n520), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n522), .A2(new_n523), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n488), .A2(new_n486), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT83), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n485), .A2(new_n491), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n478), .A2(KEYINPUT84), .A3(new_n484), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n494), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n540), .A2(KEYINPUT6), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n565), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n561), .A2(new_n445), .A3(new_n564), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n445), .A2(new_n371), .A3(new_n372), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n554), .B1(new_n566), .B2(new_n540), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n556), .A3(new_n572), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n522), .A2(new_n523), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n517), .A2(new_n508), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT75), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n517), .A2(new_n516), .A3(new_n508), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n580), .A2(new_n581), .B1(new_n513), .B2(new_n514), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n565), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n574), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n248), .B1(new_n560), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT7), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n482), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G99gat), .B(G106gat), .Z(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT97), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G57gat), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT95), .B1(new_n601), .B2(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n603));
  INV_X1    g402(.A(G64gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(G57gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n602), .B(new_n605), .C1(G57gat), .C2(new_n604), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT96), .ZN(new_n607));
  NAND2_X1  g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  OR2_X1    g407(.A1(G71gat), .A2(G78gat), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT9), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G57gat), .B(G64gat), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n608), .B(new_n609), .C1(new_n613), .C2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n612), .A2(new_n614), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n595), .A2(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n595), .A2(KEYINPUT99), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n596), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n598), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n600), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n616), .B2(new_n621), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G176gat), .ZN(new_n632));
  INV_X1    g431(.A(G204gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n626), .A2(new_n637), .A3(new_n627), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n629), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n635), .B1(new_n639), .B2(new_n634), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n626), .B2(new_n627), .ZN(new_n643));
  INV_X1    g442(.A(new_n627), .ZN(new_n644));
  AOI211_X1 g443(.A(KEYINPUT100), .B(new_n644), .C1(new_n623), .C2(new_n625), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n630), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n634), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(KEYINPUT101), .A3(new_n635), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n206), .B1(new_n617), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n296), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n653));
  NAND2_X1  g452(.A1(G231gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n657));
  XOR2_X1   g456(.A(G127gat), .B(G155gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G211gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n656), .A2(new_n661), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT41), .ZN(new_n666));
  XNOR2_X1  g465(.A(G190gat), .B(G218gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n600), .B1(new_n221), .B2(new_n223), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n624), .A2(new_n220), .B1(KEYINPUT41), .B2(new_n665), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT98), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n675), .B1(new_n673), .B2(new_n677), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n669), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n668), .A3(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n650), .A2(new_n664), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n589), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n571), .A2(new_n572), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(G1gat), .Z(G1324gat));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n564), .ZN(new_n693));
  INV_X1    g492(.A(G8gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(KEYINPUT103), .B(G8gat), .C1(new_n688), .C2(new_n564), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  AND3_X1   g497(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n693), .B2(new_n698), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n695), .B(new_n696), .C1(new_n699), .C2(new_n700), .ZN(G1325gat));
  OAI21_X1  g500(.A(G15gat), .B1(new_n688), .B2(new_n374), .ZN(new_n702));
  INV_X1    g501(.A(new_n561), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n688), .B2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n688), .A2(new_n445), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(new_n684), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n560), .B2(new_n585), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n525), .A2(KEYINPUT104), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n446), .B(new_n713), .C1(new_n495), .C2(new_n524), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n712), .A2(new_n374), .A3(new_n559), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n709), .B1(new_n715), .B2(new_n585), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n718));
  OAI22_X1  g517(.A1(new_n710), .A2(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(new_n664), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n650), .A2(new_n248), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(G29gat), .B1(new_n722), .B2(new_n689), .ZN(new_n723));
  INV_X1    g522(.A(new_n664), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(new_n650), .A3(new_n709), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n587), .B2(new_n588), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n216), .A3(new_n495), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(KEYINPUT45), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(KEYINPUT45), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n723), .B1(new_n729), .B2(new_n730), .ZN(G1328gat));
  AND3_X1   g530(.A1(new_n727), .A2(new_n217), .A3(new_n524), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT46), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  OAI21_X1  g534(.A(G36gat), .B1(new_n722), .B2(new_n564), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n727), .A2(new_n738), .A3(new_n561), .ZN(new_n739));
  INV_X1    g538(.A(new_n374), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n719), .A2(new_n740), .A3(new_n664), .A4(new_n721), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n739), .B2(new_n742), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT47), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n739), .A2(new_n742), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n747), .A2(new_n751), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n722), .B2(new_n445), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n727), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(G50gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n446), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n727), .A2(new_n754), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n753), .B(KEYINPUT48), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  AND3_X1   g562(.A1(new_n648), .A2(KEYINPUT101), .A3(new_n635), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT101), .B1(new_n648), .B2(new_n635), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n247), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n767), .A2(new_n724), .A3(new_n709), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n715), .A2(new_n585), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n689), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(new_n601), .ZN(G1332gat));
  INV_X1    g573(.A(new_n772), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n564), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n777), .B(new_n778), .Z(G1333gat));
  AOI21_X1  g578(.A(new_n341), .B1(new_n775), .B2(new_n740), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n772), .A2(G71gat), .A3(new_n703), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT109), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT109), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(KEYINPUT50), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n775), .A2(new_n446), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G78gat), .ZN(G1335gat));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n771), .A2(new_n792), .A3(new_n684), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n664), .A2(new_n248), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n716), .A2(new_n792), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n716), .B2(new_n792), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n574), .A2(new_n584), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n564), .A2(new_n689), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n713), .B1(new_n801), .B2(new_n446), .ZN(new_n802));
  AOI211_X1 g601(.A(KEYINPUT104), .B(new_n445), .C1(new_n564), .C2(new_n689), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n541), .A2(KEYINPUT40), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(new_n485), .A3(new_n538), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n446), .B1(new_n806), .B2(new_n524), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(new_n558), .B1(new_n370), .B2(new_n373), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n800), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT110), .B1(new_n809), .B2(new_n709), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n799), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n798), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n766), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n482), .A3(new_n495), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n720), .A2(new_n767), .ZN(new_n816));
  OAI21_X1  g615(.A(G85gat), .B1(new_n816), .B2(new_n689), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1336gat));
  OAI21_X1  g617(.A(G92gat), .B1(new_n816), .B2(new_n564), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n650), .A2(new_n593), .A3(new_n524), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT111), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n819), .B(new_n824), .C1(new_n813), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1337gat));
  INV_X1    g625(.A(G99gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n814), .A2(new_n827), .A3(new_n561), .ZN(new_n828));
  OAI21_X1  g627(.A(G99gat), .B1(new_n816), .B2(new_n374), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1338gat));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n445), .A2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n799), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n799), .B2(new_n810), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n650), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n719), .A2(new_n446), .A3(new_n664), .A4(new_n767), .ZN(new_n838));
  AOI22_X1  g637(.A1(new_n837), .A2(KEYINPUT112), .B1(G106gat), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n812), .A2(new_n840), .A3(new_n650), .A4(new_n834), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n832), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(G106gat), .ZN(new_n843));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n831), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n837), .A2(KEYINPUT112), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(new_n841), .A3(new_n843), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(KEYINPUT114), .A3(new_n845), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(G1339gat));
  NAND2_X1  g651(.A1(new_n685), .A2(new_n248), .ZN(new_n853));
  XOR2_X1   g652(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n636), .A2(new_n638), .A3(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n626), .B2(new_n627), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n623), .A2(new_n644), .A3(new_n625), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n634), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT55), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n856), .A2(new_n860), .A3(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n635), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n227), .B1(new_n224), .B2(new_n228), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n233), .A2(new_n235), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n242), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n246), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n684), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n864), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n764), .B2(new_n765), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n650), .A2(KEYINPUT117), .A3(new_n871), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n247), .A2(new_n635), .A3(new_n865), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n878), .B1(new_n862), .B2(new_n863), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(new_n709), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n853), .B1(new_n881), .B2(new_n724), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n495), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n883), .A2(new_n575), .A3(new_n524), .ZN(new_n884));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884), .B2(new_n247), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n882), .A2(new_n445), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n703), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n689), .A2(new_n524), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n882), .A2(KEYINPUT118), .A3(new_n445), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n248), .A2(new_n300), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(G1340gat));
  AOI21_X1  g692(.A(G120gat), .B1(new_n884), .B2(new_n650), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n766), .A2(new_n301), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n894), .B1(new_n891), .B2(new_n895), .ZN(G1341gat));
  AOI21_X1  g695(.A(KEYINPUT119), .B1(new_n884), .B2(new_n724), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(G127gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n884), .A2(KEYINPUT119), .A3(new_n724), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n664), .A2(new_n307), .ZN(new_n900));
  AOI22_X1  g699(.A1(new_n898), .A2(new_n899), .B1(new_n891), .B2(new_n900), .ZN(G1342gat));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n315), .A3(new_n316), .A4(new_n684), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT56), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n684), .A3(new_n889), .A4(new_n890), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n905), .B2(G134gat), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n903), .B(new_n904), .C1(new_n906), .C2(new_n907), .ZN(G1343gat));
  NOR2_X1   g707(.A1(new_n740), .A2(new_n445), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n883), .A2(new_n524), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n396), .A3(new_n247), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n874), .A2(KEYINPUT121), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n650), .A2(new_n916), .A3(new_n871), .ZN(new_n917));
  INV_X1    g716(.A(new_n861), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n878), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n873), .B1(new_n920), .B2(new_n709), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n914), .B1(new_n921), .B2(new_n724), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n870), .B1(new_n642), .B2(new_n649), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n923), .A2(new_n916), .B1(new_n918), .B2(new_n878), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n684), .B1(new_n924), .B2(new_n915), .ZN(new_n925));
  OAI211_X1 g724(.A(KEYINPUT122), .B(new_n664), .C1(new_n925), .C2(new_n873), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n853), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n913), .B1(new_n927), .B2(new_n446), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n374), .A2(new_n889), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n882), .A2(new_n446), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(KEYINPUT57), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n928), .A2(new_n931), .A3(new_n248), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n912), .B1(new_n932), .B2(new_n396), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT58), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n935), .B(new_n912), .C1(new_n932), .C2(new_n396), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(G1344gat));
  NAND3_X1  g736(.A1(new_n911), .A2(new_n397), .A3(new_n650), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n930), .A2(KEYINPUT57), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n687), .A2(new_n248), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n921), .A2(new_n724), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n913), .B(new_n446), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n650), .A3(new_n929), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n939), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n928), .A2(new_n931), .A3(new_n766), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(KEYINPUT59), .A3(new_n397), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n938), .B1(new_n946), .B2(new_n948), .ZN(G1345gat));
  NAND3_X1  g748(.A1(new_n911), .A2(new_n379), .A3(new_n724), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n928), .A2(new_n931), .A3(new_n664), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n379), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT123), .B(new_n950), .C1(new_n951), .C2(new_n379), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  NOR2_X1   g755(.A1(new_n910), .A2(new_n524), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n709), .A2(G162gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n882), .A2(new_n495), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n928), .A2(new_n931), .A3(new_n709), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n961), .B2(new_n380), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n964), .B(new_n960), .C1(new_n961), .C2(new_n380), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n495), .A2(new_n564), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n888), .A2(new_n890), .A3(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n240), .A3(new_n248), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n882), .A2(new_n689), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n575), .A2(new_n564), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(G169gat), .B1(new_n972), .B2(new_n247), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n969), .A2(new_n973), .ZN(G1348gat));
  OAI21_X1  g773(.A(G176gat), .B1(new_n968), .B2(new_n766), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n276), .A3(new_n650), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1349gat));
  NAND4_X1  g776(.A1(new_n888), .A2(new_n724), .A3(new_n890), .A4(new_n967), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n268), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n972), .A2(new_n261), .A3(new_n724), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT60), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT60), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n979), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1350gat));
  AND4_X1   g784(.A1(new_n253), .A2(new_n970), .A3(new_n684), .A4(new_n971), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT126), .ZN(new_n987));
  OAI21_X1  g786(.A(G190gat), .B1(new_n968), .B2(new_n709), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g789(.A(KEYINPUT61), .B(G190gat), .C1(new_n968), .C2(new_n709), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(G1351gat));
  INV_X1    g791(.A(G197gat), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n910), .A2(new_n564), .ZN(new_n994));
  AND4_X1   g793(.A1(new_n993), .A2(new_n970), .A3(new_n247), .A4(new_n994), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  XNOR2_X1  g795(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n374), .A2(new_n967), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  AND3_X1   g798(.A1(new_n940), .A2(new_n943), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n1000), .A2(new_n247), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n997), .B1(new_n993), .B2(new_n1001), .ZN(G1352gat));
  AND2_X1   g801(.A1(new_n970), .A2(new_n994), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1003), .A2(new_n633), .A3(new_n650), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n944), .A2(new_n650), .A3(new_n999), .ZN(new_n1007));
  OAI211_X1 g806(.A(new_n1005), .B(new_n1006), .C1(new_n633), .C2(new_n1007), .ZN(G1353gat));
  NAND3_X1  g807(.A1(new_n1003), .A2(new_n660), .A3(new_n724), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1000), .A2(new_n724), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT63), .B1(new_n1010), .B2(G211gat), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT63), .ZN(new_n1012));
  AOI211_X1 g811(.A(new_n1012), .B(new_n660), .C1(new_n1000), .C2(new_n724), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1009), .B1(new_n1011), .B2(new_n1013), .ZN(G1354gat));
  AOI21_X1  g813(.A(G218gat), .B1(new_n1003), .B2(new_n684), .ZN(new_n1015));
  AND2_X1   g814(.A1(new_n684), .A2(G218gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1015), .B1(new_n1000), .B2(new_n1016), .ZN(G1355gat));
endmodule


