//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954;
  INV_X1    g000(.A(G43gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT87), .B(G50gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G43gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n202), .A2(G50gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n203), .A2(KEYINPUT15), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT85), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n211), .A2(KEYINPUT14), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT85), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n215), .A2(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n220), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT88), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n225), .B(new_n226), .C1(G1gat), .C2(new_n223), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n227), .B(G8gat), .C1(new_n226), .C2(new_n225), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n223), .A2(G1gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(new_n229), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n217), .A2(new_n219), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT91), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(KEYINPUT18), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT93), .B1(new_n241), .B2(new_n238), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(new_n242), .Z(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(new_n243), .ZN(new_n250));
  OR2_X1    g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(KEYINPUT18), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G169gat), .B(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n261), .A3(new_n251), .A4(new_n252), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(KEYINPUT94), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT94), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n253), .A2(new_n264), .A3(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(KEYINPUT95), .A3(new_n265), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273));
  INV_X1    g072(.A(G211gat), .ZN(new_n274));
  INV_X1    g073(.A(G218gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g076(.A(G211gat), .B(G218gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT78), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G155gat), .B2(G162gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(G155gat), .B2(G162gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G155gat), .B(G162gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT2), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(new_n288), .A3(new_n283), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n281), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT3), .B1(new_n279), .B2(new_n303), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n290), .A2(KEYINPUT79), .A3(new_n299), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT79), .B1(new_n290), .B2(new_n299), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n306), .B2(new_n300), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n311), .A2(new_n312), .B1(new_n305), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G78gat), .B(G106gat), .Z(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G22gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n314), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G226gat), .ZN(new_n320));
  INV_X1    g119(.A(G233gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n323), .A2(KEYINPUT26), .ZN(new_n324));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(KEYINPUT26), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT28), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT28), .B1(new_n329), .B2(new_n330), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n327), .B(new_n328), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(KEYINPUT23), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n323), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(KEYINPUT23), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n328), .A2(new_n341), .A3(KEYINPUT24), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT67), .ZN(new_n344));
  AND2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n340), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n330), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n344), .A3(new_n328), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n345), .A2(KEYINPUT67), .A3(new_n343), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n336), .A3(new_n339), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT68), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  AND2_X1   g157(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT66), .A2(G176gat), .ZN(new_n360));
  OAI211_X1 g159(.A(KEYINPUT23), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n336), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n351), .A2(new_n330), .A3(KEYINPUT65), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G183gat), .B2(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n345), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n328), .B1(new_n371), .B2(new_n343), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT25), .B1(new_n363), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n334), .B1(new_n357), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n322), .B1(new_n375), .B2(new_n303), .ZN(new_n376));
  INV_X1    g175(.A(new_n322), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n367), .A2(new_n370), .A3(new_n372), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n337), .B1(new_n378), .B2(new_n362), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n379), .A2(new_n356), .A3(new_n350), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n380), .B2(new_n334), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n281), .ZN(new_n383));
  INV_X1    g182(.A(new_n281), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n376), .B2(new_n381), .ZN(new_n385));
  XOR2_X1   g184(.A(G8gat), .B(G36gat), .Z(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(G92gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(G64gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n383), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT30), .ZN(new_n392));
  INV_X1    g191(.A(new_n385), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n376), .A2(new_n384), .A3(new_n381), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n392), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT69), .ZN(new_n397));
  INV_X1    g196(.A(G134gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n399), .A2(KEYINPUT1), .A3(G127gat), .ZN(new_n400));
  INV_X1    g199(.A(G127gat), .ZN(new_n401));
  INV_X1    g200(.A(G120gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(G113gat), .ZN(new_n403));
  INV_X1    g202(.A(G113gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G120gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n398), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(G127gat), .B1(new_n399), .B2(KEYINPUT1), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n401), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(G134gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n375), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n410), .A2(new_n411), .A3(G134gat), .ZN(new_n415));
  AOI21_X1  g214(.A(G134gat), .B1(new_n410), .B2(new_n411), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n380), .A2(new_n417), .A3(new_n334), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G227gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n321), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n397), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n421), .ZN(new_n423));
  AOI211_X1 g222(.A(KEYINPUT69), .B(new_n423), .C1(new_n414), .C2(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT32), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G15gat), .B(G43gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  AOI21_X1  g229(.A(new_n425), .B1(KEYINPUT33), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n380), .A2(new_n417), .A3(new_n334), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n417), .B1(new_n380), .B2(new_n334), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n421), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT69), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n397), .A3(new_n421), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT70), .B1(new_n439), .B2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT70), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT32), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n441), .B(new_n442), .C1(new_n437), .C2(new_n438), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n430), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n433), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n441), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n439), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n433), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n432), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n414), .A2(new_n423), .A3(new_n418), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT34), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(KEYINPUT74), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT73), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n431), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT74), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n455), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n319), .B(new_n396), .C1(new_n457), .C2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n417), .B1(new_n309), .B2(new_n307), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n290), .A2(new_n299), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n413), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(G225gat), .B(G233gat), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n290), .A2(KEYINPUT79), .A3(new_n299), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT3), .B1(new_n468), .B2(new_n308), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n413), .A3(new_n302), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n413), .C2(new_n465), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n417), .B2(new_n300), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n300), .A2(new_n409), .A3(new_n474), .A4(new_n412), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n473), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT5), .B(new_n467), .C1(new_n472), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n476), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n473), .A4(new_n470), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G1gat), .B(G29gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G85gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT0), .B(G57gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  AOI21_X1  g288(.A(KEYINPUT6), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n484), .ZN(new_n491));
  INV_X1    g290(.A(new_n489), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(KEYINPUT6), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n453), .A2(new_n455), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n460), .A2(new_n456), .ZN(new_n501));
  INV_X1    g300(.A(new_n318), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n317), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n480), .A2(new_n504), .A3(new_n484), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n480), .B2(new_n484), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n492), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n493), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n490), .B1(new_n508), .B2(KEYINPUT6), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n396), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n500), .A2(new_n501), .A3(new_n503), .A4(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n463), .A2(new_n499), .B1(new_n498), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n513), .B1(new_n393), .B2(new_n394), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT83), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT83), .B(new_n513), .C1(new_n393), .C2(new_n394), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n383), .A2(KEYINPUT37), .A3(new_n385), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(new_n390), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT38), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n393), .A2(new_n394), .A3(new_n513), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n515), .B2(new_n514), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT38), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n390), .A4(new_n517), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(new_n395), .A3(new_n520), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n491), .A2(KEYINPUT82), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n480), .A2(new_n504), .A3(new_n484), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT39), .ZN(new_n529));
  INV_X1    g328(.A(new_n470), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n475), .A2(new_n481), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n482), .A2(KEYINPUT39), .A3(new_n470), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n473), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT39), .B(new_n473), .C1(new_n464), .C2(new_n466), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n534), .A2(new_n492), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n528), .A2(new_n492), .B1(new_n537), .B2(KEYINPUT40), .ZN(new_n538));
  OR3_X1    g337(.A1(new_n534), .A2(new_n492), .A3(new_n536), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT81), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT40), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT81), .B1(new_n537), .B2(KEYINPUT40), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n538), .A2(new_n542), .A3(new_n396), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n503), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n319), .B1(new_n497), .B2(new_n396), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT36), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n457), .B2(new_n462), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n500), .B2(new_n501), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n547), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n271), .B1(new_n512), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT21), .ZN(new_n555));
  XOR2_X1   g354(.A(G71gat), .B(G78gat), .Z(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n556), .A2(KEYINPUT96), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(KEYINPUT96), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n559), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n239), .B1(new_n555), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(new_n351), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G211gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n569), .B(new_n571), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n555), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT97), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n572), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(G85gat), .A2(G92gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT7), .ZN(new_n580));
  INV_X1    g379(.A(G99gat), .ZN(new_n581));
  INV_X1    g380(.A(G106gat), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT8), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n580), .B(new_n583), .C1(G85gat), .C2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G99gat), .B(G106gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  NAND2_X1  g385(.A1(new_n222), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT98), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n220), .A2(new_n586), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n222), .A2(new_n590), .A3(new_n586), .ZN(new_n591));
  NAND3_X1  g390(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  OR3_X1    g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n596), .A2(new_n597), .B1(new_n595), .B2(new_n593), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT100), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n598), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n598), .A2(new_n599), .A3(new_n603), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n578), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n586), .A2(new_n565), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n586), .B(new_n565), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n612), .A2(KEYINPUT102), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT102), .B1(new_n612), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(G230gat), .A3(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n621), .B(KEYINPUT101), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n612), .A2(new_n613), .ZN(new_n624));
  INV_X1    g423(.A(new_n621), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n617), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n554), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n497), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  INV_X1    g433(.A(new_n396), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n224), .A2(new_n233), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n641), .B(new_n642), .C1(new_n233), .C2(new_n636), .ZN(G1325gat));
  INV_X1    g442(.A(G15gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n549), .A2(new_n552), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n631), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n500), .A2(new_n501), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n644), .B2(new_n650), .ZN(G1326gat));
  NOR2_X1   g450(.A1(new_n631), .A2(new_n503), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT43), .B(G22gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1327gat));
  NAND2_X1  g453(.A1(new_n553), .A2(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n547), .B(new_n656), .C1(new_n549), .C2(new_n552), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n512), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n596), .A2(new_n597), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n593), .A2(new_n595), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n663), .A3(new_n602), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n604), .A3(KEYINPUT104), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT104), .B1(new_n664), .B2(new_n604), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n658), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n553), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n457), .A2(new_n462), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n672), .A2(new_n503), .A3(new_n635), .A4(new_n499), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n511), .A2(new_n498), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n607), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n577), .A2(new_n627), .ZN(new_n679));
  INV_X1    g478(.A(new_n266), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n496), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n554), .A2(new_n607), .A3(new_n679), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n685), .A2(G29gat), .A3(new_n496), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(KEYINPUT45), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(KEYINPUT45), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n684), .B1(new_n687), .B2(new_n688), .ZN(G1328gat));
  OR2_X1    g488(.A1(new_n685), .A2(new_n635), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n691));
  OAI22_X1  g490(.A1(new_n690), .A2(G36gat), .B1(new_n691), .B2(KEYINPUT46), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(KEYINPUT105), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G36gat), .B1(new_n683), .B2(new_n635), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n691), .B(KEYINPUT46), .C1(new_n690), .C2(G36gat), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(G1329gat));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n678), .A2(new_n645), .A3(new_n682), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n685), .A2(G43gat), .A3(new_n648), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(KEYINPUT106), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n678), .A2(new_n704), .A3(new_n645), .A4(new_n682), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(G43gat), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n701), .A2(new_n698), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT107), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(G1330gat));
  AOI211_X1 g509(.A(new_n503), .B(new_n681), .C1(new_n670), .C2(new_n677), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT108), .B1(new_n711), .B2(new_n204), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n685), .A2(new_n503), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n204), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n678), .A2(new_n319), .A3(new_n682), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n716));
  INV_X1    g515(.A(new_n204), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT109), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n678), .A2(new_n723), .A3(new_n319), .A4(new_n682), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n720), .B1(new_n713), .B2(new_n204), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n725), .A2(KEYINPUT110), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n721), .B1(new_n727), .B2(new_n728), .ZN(G1331gat));
  AND2_X1   g528(.A1(new_n658), .A2(new_n608), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n680), .A2(new_n628), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n496), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n732), .A2(new_n635), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  NOR2_X1   g541(.A1(new_n732), .A2(new_n648), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n645), .A2(G71gat), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n743), .A2(G71gat), .B1(new_n732), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n745), .B(new_n746), .Z(G1334gat));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n503), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT113), .B(G78gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1335gat));
  NAND3_X1  g549(.A1(new_n678), .A2(new_n578), .A3(new_n731), .ZN(new_n751));
  INV_X1    g550(.A(G85gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n496), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n658), .A2(new_n266), .A3(new_n607), .A4(new_n578), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n497), .A3(new_n627), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n757), .B2(new_n752), .ZN(G1336gat));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  OAI21_X1  g558(.A(G92gat), .B1(new_n751), .B2(new_n635), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n627), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n635), .A2(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n755), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n754), .A2(new_n765), .A3(KEYINPUT51), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n767), .A2(new_n627), .A3(new_n762), .A4(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n769), .A2(new_n760), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n770), .B2(new_n759), .ZN(G1337gat));
  OAI21_X1  g570(.A(G99gat), .B1(new_n751), .B2(new_n646), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n649), .A2(new_n581), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n761), .B2(new_n773), .ZN(G1338gat));
  OR2_X1    g573(.A1(new_n751), .A2(new_n503), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G106gat), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n628), .A2(G106gat), .A3(new_n503), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT53), .B1(new_n756), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n767), .A2(new_n768), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n780), .A2(new_n777), .B1(new_n775), .B2(G106gat), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  NOR4_X1   g582(.A1(new_n578), .A2(new_n607), .A3(new_n680), .A4(new_n627), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n248), .A2(KEYINPUT116), .A3(new_n250), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT116), .B1(new_n248), .B2(new_n250), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n240), .A2(new_n242), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(G229gat), .A3(G233gat), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT117), .B(new_n262), .C1(new_n790), .C2(new_n258), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792));
  INV_X1    g591(.A(new_n262), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n258), .B1(new_n787), .B2(new_n789), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n614), .B2(new_n615), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n612), .A2(new_n613), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(KEYINPUT54), .A3(new_n624), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n621), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .A4(new_n621), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n804), .A2(KEYINPUT115), .A3(new_n626), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n804), .B2(new_n626), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n796), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n666), .B2(new_n667), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n627), .B(new_n262), .C1(new_n790), .C2(new_n258), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n807), .B2(new_n266), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n664), .A2(new_n604), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT104), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n811), .A2(new_n814), .A3(new_n665), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n784), .B1(new_n816), .B2(new_n578), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(new_n648), .A3(new_n319), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n818), .A2(new_n497), .A3(new_n635), .ZN(new_n819));
  OAI21_X1  g618(.A(G113gat), .B1(new_n819), .B2(new_n271), .ZN(new_n820));
  INV_X1    g619(.A(new_n735), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n822), .A2(new_n463), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n404), .A3(new_n680), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(G1340gat));
  OAI21_X1  g624(.A(G120gat), .B1(new_n819), .B2(new_n628), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n402), .A3(new_n627), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n823), .B2(new_n577), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n819), .A2(new_n401), .A3(new_n578), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  NAND3_X1  g630(.A1(new_n823), .A2(new_n398), .A3(new_n607), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n833));
  OAI21_X1  g632(.A(G134gat), .B1(new_n819), .B2(new_n812), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(KEYINPUT56), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(G1343gat));
  NOR3_X1   g635(.A1(new_n645), .A2(new_n496), .A3(new_n396), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n577), .B1(new_n809), .B2(new_n815), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n838), .B(new_n319), .C1(new_n839), .C2(new_n784), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n804), .A2(new_n626), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n268), .A2(new_n269), .A3(new_n803), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n607), .B1(new_n843), .B2(new_n810), .ZN(new_n844));
  INV_X1    g643(.A(new_n809), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n578), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n784), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n503), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n837), .B(new_n840), .C1(new_n848), .C2(new_n838), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n271), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n645), .A2(new_n503), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n822), .A2(new_n635), .A3(new_n270), .A4(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n850), .B(new_n851), .C1(G141gat), .C2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G141gat), .B1(new_n849), .B2(new_n266), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n822), .A2(new_n635), .A3(new_n852), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n294), .A4(new_n270), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT118), .B1(new_n853), .B2(G141gat), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n854), .B1(new_n860), .B2(new_n851), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n856), .A2(new_n295), .A3(new_n627), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n810), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n812), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n808), .A2(new_n607), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n577), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n629), .A2(new_n270), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n838), .B(new_n319), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT57), .B1(new_n817), .B2(new_n503), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n627), .A3(new_n837), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n863), .B1(new_n872), .B2(G148gat), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n863), .B(G148gat), .C1(new_n849), .C2(new_n628), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n862), .B1(new_n873), .B2(new_n875), .ZN(G1345gat));
  NOR3_X1   g675(.A1(new_n849), .A2(new_n291), .A3(new_n578), .ZN(new_n877));
  AOI21_X1  g676(.A(G155gat), .B1(new_n856), .B2(new_n577), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n292), .A3(new_n607), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G162gat), .B1(new_n849), .B2(new_n668), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1347gat));
  NAND2_X1  g683(.A1(new_n672), .A2(new_n503), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n817), .B2(new_n497), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT120), .B(new_n496), .C1(new_n839), .C2(new_n784), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n889), .A2(new_n358), .A3(new_n396), .A4(new_n680), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n821), .A2(new_n396), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT122), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n649), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(KEYINPUT123), .A3(new_n649), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n816), .A2(new_n578), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n319), .B1(new_n900), .B2(new_n847), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n270), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G169gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n892), .A2(new_n904), .ZN(G1348gat));
  AND2_X1   g704(.A1(new_n889), .A2(new_n396), .ZN(new_n906));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906), .B2(new_n627), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n628), .A2(new_n360), .A3(new_n359), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n902), .B2(new_n908), .ZN(G1349gat));
  NAND4_X1  g708(.A1(new_n901), .A2(new_n577), .A3(new_n897), .A4(new_n898), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n899), .A2(KEYINPUT124), .A3(new_n577), .A4(new_n901), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(G183gat), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n889), .A2(new_n329), .A3(new_n396), .A4(new_n577), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(KEYINPUT125), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT60), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT125), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1350gat));
  NAND2_X1  g719(.A1(new_n902), .A2(new_n607), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G190gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n668), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n330), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n924), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n921), .A2(G190gat), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n894), .A2(new_n646), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n871), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n271), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n852), .A2(new_n396), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n888), .B2(new_n887), .ZN(new_n937));
  INV_X1    g736(.A(G197gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(new_n680), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n934), .A2(new_n939), .ZN(G1352gat));
  INV_X1    g739(.A(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n937), .A2(new_n941), .A3(new_n627), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n937), .A2(new_n944), .A3(new_n941), .A4(new_n627), .ZN(new_n945));
  AND3_X1   g744(.A1(new_n871), .A2(new_n627), .A3(new_n932), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n943), .B(new_n945), .C1(new_n941), .C2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n937), .A2(new_n274), .A3(new_n577), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n869), .A2(new_n577), .A3(new_n870), .A4(new_n932), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT63), .B1(new_n949), .B2(G211gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1354gat));
  OAI21_X1  g751(.A(G218gat), .B1(new_n933), .B2(new_n812), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n275), .A3(new_n926), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


