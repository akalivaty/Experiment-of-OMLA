

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578;

  XNOR2_X1 U320 ( .A(G120GAT), .B(n399), .ZN(n288) );
  XNOR2_X1 U321 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n411) );
  XNOR2_X1 U322 ( .A(n412), .B(n411), .ZN(n413) );
  NOR2_X1 U323 ( .A1(n420), .A2(n419), .ZN(n421) );
  NOR2_X1 U324 ( .A1(n505), .A2(n425), .ZN(n563) );
  INV_X1 U325 ( .A(G190GAT), .ZN(n445) );
  XNOR2_X1 U326 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U327 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(G29GAT), .B(KEYINPUT7), .Z(n290) );
  XNOR2_X1 U329 ( .A(G43GAT), .B(G36GAT), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n290), .B(n289), .ZN(n292) );
  XOR2_X1 U331 ( .A(G50GAT), .B(KEYINPUT8), .Z(n291) );
  XOR2_X1 U332 ( .A(n292), .B(n291), .Z(n393) );
  INV_X1 U333 ( .A(n393), .ZN(n310) );
  XOR2_X1 U334 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n294) );
  XNOR2_X1 U335 ( .A(G99GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(G85GAT), .B(n295), .Z(n406) );
  XOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT79), .Z(n357) );
  XOR2_X1 U339 ( .A(KEYINPUT10), .B(n357), .Z(n297) );
  XNOR2_X1 U340 ( .A(G134GAT), .B(G218GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(n406), .B(n298), .Z(n300) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n302) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(KEYINPUT65), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U348 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n304) );
  XNOR2_X1 U349 ( .A(G162GAT), .B(KEYINPUT78), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U353 ( .A(n310), .B(n309), .Z(n546) );
  XOR2_X1 U354 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n312) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n350) );
  XOR2_X1 U357 ( .A(n350), .B(G71GAT), .Z(n314) );
  NAND2_X1 U358 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U360 ( .A(G176GAT), .B(KEYINPUT20), .Z(n316) );
  XNOR2_X1 U361 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U363 ( .A(n318), .B(n317), .Z(n327) );
  XNOR2_X1 U364 ( .A(G127GAT), .B(G134GAT), .ZN(n319) );
  XNOR2_X1 U365 ( .A(n319), .B(KEYINPUT0), .ZN(n320) );
  XOR2_X1 U366 ( .A(n320), .B(KEYINPUT86), .Z(n322) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(G120GAT), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n341) );
  XOR2_X1 U369 ( .A(G183GAT), .B(G190GAT), .Z(n324) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G99GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U372 ( .A(n341), .B(n325), .ZN(n326) );
  XOR2_X1 U373 ( .A(n327), .B(n326), .Z(n521) );
  INV_X1 U374 ( .A(n521), .ZN(n511) );
  XOR2_X1 U375 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n443) );
  XOR2_X1 U376 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT91), .B(KEYINPUT4), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n345) );
  XOR2_X1 U379 ( .A(G85GAT), .B(G155GAT), .Z(n331) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(G148GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U382 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n333) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U385 ( .A(n335), .B(n334), .Z(n343) );
  XOR2_X1 U386 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n337) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(G162GAT), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n436) );
  XOR2_X1 U389 ( .A(n436), .B(KEYINPUT93), .Z(n339) );
  NAND2_X1 U390 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U394 ( .A(n345), .B(n344), .ZN(n518) );
  INV_X1 U395 ( .A(n518), .ZN(n505) );
  INV_X1 U396 ( .A(KEYINPUT54), .ZN(n424) );
  XOR2_X1 U397 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n347) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(G218GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n437) );
  XOR2_X1 U400 ( .A(KEYINPUT80), .B(G211GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(G8GAT), .B(G183GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n437), .B(n368), .ZN(n361) );
  XOR2_X1 U404 ( .A(n350), .B(KEYINPUT94), .Z(n352) );
  NAND2_X1 U405 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT95), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(n356), .B(n355), .Z(n359) );
  XOR2_X1 U411 ( .A(G176GAT), .B(G64GAT), .Z(n399) );
  XNOR2_X1 U412 ( .A(n357), .B(n399), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U414 ( .A(n361), .B(n360), .Z(n507) );
  INV_X1 U415 ( .A(n507), .ZN(n422) );
  XOR2_X1 U416 ( .A(G22GAT), .B(G155GAT), .Z(n426) );
  XOR2_X1 U417 ( .A(KEYINPUT82), .B(KEYINPUT85), .Z(n363) );
  XNOR2_X1 U418 ( .A(G127GAT), .B(G64GAT), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U420 ( .A(n426), .B(n364), .Z(n366) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U423 ( .A(n367), .B(KEYINPUT81), .Z(n370) );
  XNOR2_X1 U424 ( .A(n368), .B(KEYINPUT14), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U426 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n379) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G1GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n375), .B(KEYINPUT68), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT13), .B(G57GAT), .Z(n377) );
  XNOR2_X1 U433 ( .A(G71GAT), .B(G78GAT), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n398) );
  XNOR2_X1 U435 ( .A(n382), .B(n398), .ZN(n378) );
  XOR2_X1 U436 ( .A(n379), .B(n378), .Z(n573) );
  XNOR2_X1 U437 ( .A(n573), .B(KEYINPUT111), .ZN(n558) );
  XOR2_X1 U438 ( .A(KEYINPUT67), .B(KEYINPUT29), .Z(n381) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G8GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n392) );
  XOR2_X1 U441 ( .A(G113GAT), .B(n382), .Z(n384) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(G141GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n385), .B(G197GAT), .Z(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n387) );
  NAND2_X1 U446 ( .A1(G229GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U447 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U448 ( .A(KEYINPUT69), .B(n388), .ZN(n389) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n564) );
  XNOR2_X1 U452 ( .A(G106GAT), .B(G204GAT), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n395), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U454 ( .A(n427), .B(KEYINPUT75), .Z(n397) );
  NAND2_X1 U455 ( .A1(G230GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n402) );
  XNOR2_X1 U457 ( .A(KEYINPUT33), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n400), .B(n288), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n404) );
  XNOR2_X1 U461 ( .A(KEYINPUT74), .B(KEYINPUT31), .ZN(n403) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n568) );
  INV_X1 U465 ( .A(KEYINPUT64), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n568), .B(n409), .ZN(n410) );
  XOR2_X1 U467 ( .A(KEYINPUT41), .B(n410), .Z(n524) );
  INV_X1 U468 ( .A(n524), .ZN(n555) );
  NOR2_X1 U469 ( .A1(n564), .A2(n555), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n558), .A2(n413), .ZN(n414) );
  NAND2_X1 U471 ( .A1(n546), .A2(n414), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n415), .B(KEYINPUT47), .ZN(n420) );
  XOR2_X1 U473 ( .A(KEYINPUT70), .B(n564), .Z(n548) );
  INV_X1 U474 ( .A(n546), .ZN(n532) );
  XOR2_X1 U475 ( .A(KEYINPUT36), .B(n532), .Z(n576) );
  NOR2_X1 U476 ( .A1(n576), .A2(n573), .ZN(n416) );
  XNOR2_X1 U477 ( .A(KEYINPUT45), .B(n416), .ZN(n417) );
  NAND2_X1 U478 ( .A1(n417), .A2(n568), .ZN(n418) );
  NOR2_X1 U479 ( .A1(n548), .A2(n418), .ZN(n419) );
  XNOR2_X1 U480 ( .A(KEYINPUT48), .B(n421), .ZN(n517) );
  NOR2_X1 U481 ( .A1(n422), .A2(n517), .ZN(n423) );
  XNOR2_X1 U482 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n441) );
  XOR2_X1 U486 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U489 ( .A(G78GAT), .B(G211GAT), .Z(n433) );
  XNOR2_X1 U490 ( .A(G50GAT), .B(KEYINPUT90), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U492 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n454) );
  NAND2_X1 U496 ( .A1(n563), .A2(n454), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n443), .B(n442), .ZN(n444) );
  NAND2_X1 U498 ( .A1(n511), .A2(n444), .ZN(n554) );
  NOR2_X1 U499 ( .A1(n546), .A2(n554), .ZN(n448) );
  XNOR2_X1 U500 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n446) );
  NAND2_X1 U501 ( .A1(n568), .A2(n548), .ZN(n479) );
  NOR2_X1 U502 ( .A1(n532), .A2(n573), .ZN(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT16), .B(n449), .ZN(n465) );
  XNOR2_X1 U504 ( .A(n507), .B(KEYINPUT96), .ZN(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT27), .B(n450), .Z(n457) );
  XOR2_X1 U506 ( .A(n454), .B(KEYINPUT28), .Z(n513) );
  NOR2_X1 U507 ( .A1(n457), .A2(n513), .ZN(n519) );
  NAND2_X1 U508 ( .A1(n521), .A2(n519), .ZN(n451) );
  NAND2_X1 U509 ( .A1(n451), .A2(n505), .ZN(n463) );
  NAND2_X1 U510 ( .A1(n511), .A2(n507), .ZN(n452) );
  NAND2_X1 U511 ( .A1(n454), .A2(n452), .ZN(n453) );
  XOR2_X1 U512 ( .A(KEYINPUT25), .B(n453), .Z(n461) );
  NOR2_X1 U513 ( .A1(n511), .A2(n454), .ZN(n455) );
  XOR2_X1 U514 ( .A(KEYINPUT97), .B(n455), .Z(n456) );
  XNOR2_X1 U515 ( .A(KEYINPUT26), .B(n456), .ZN(n562) );
  INV_X1 U516 ( .A(n562), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n458), .A2(n457), .ZN(n537) );
  XNOR2_X1 U518 ( .A(KEYINPUT98), .B(n537), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n505), .A2(n459), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n476) );
  INV_X1 U522 ( .A(n476), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n493) );
  NOR2_X1 U524 ( .A1(n479), .A2(n493), .ZN(n473) );
  NAND2_X1 U525 ( .A1(n473), .A2(n505), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT34), .ZN(n467) );
  XNOR2_X1 U527 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  XOR2_X1 U528 ( .A(G8GAT), .B(KEYINPUT99), .Z(n469) );
  NAND2_X1 U529 ( .A1(n473), .A2(n507), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(G1325GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n471) );
  NAND2_X1 U532 ( .A1(n473), .A2(n511), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(n472), .ZN(G1326GAT) );
  XOR2_X1 U535 ( .A(G22GAT), .B(KEYINPUT101), .Z(n475) );
  NAND2_X1 U536 ( .A1(n473), .A2(n513), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n475), .B(n474), .ZN(G1327GAT) );
  XOR2_X1 U538 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n483) );
  NOR2_X1 U539 ( .A1(n576), .A2(n476), .ZN(n477) );
  NAND2_X1 U540 ( .A1(n573), .A2(n477), .ZN(n478) );
  XOR2_X1 U541 ( .A(KEYINPUT37), .B(n478), .Z(n504) );
  NOR2_X1 U542 ( .A1(n504), .A2(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(n490) );
  NAND2_X1 U545 ( .A1(n490), .A2(n505), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U547 ( .A(G29GAT), .B(n484), .Z(G1328GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n486) );
  NAND2_X1 U549 ( .A1(n490), .A2(n507), .ZN(n485) );
  XNOR2_X1 U550 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(n487), .ZN(G1329GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n511), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n488), .B(KEYINPUT40), .ZN(n489) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NAND2_X1 U555 ( .A1(n490), .A2(n513), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n491), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n492), .ZN(G1331GAT) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n495) );
  NAND2_X1 U559 ( .A1(n524), .A2(n564), .ZN(n503) );
  NOR2_X1 U560 ( .A1(n503), .A2(n493), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n505), .A2(n499), .ZN(n494) );
  XNOR2_X1 U562 ( .A(n495), .B(n494), .ZN(G1332GAT) );
  XOR2_X1 U563 ( .A(G64GAT), .B(KEYINPUT107), .Z(n497) );
  NAND2_X1 U564 ( .A1(n499), .A2(n507), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NAND2_X1 U566 ( .A1(n499), .A2(n511), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n501) );
  NAND2_X1 U569 ( .A1(n499), .A2(n513), .ZN(n500) );
  XNOR2_X1 U570 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(n502), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n504), .A2(n503), .ZN(n514) );
  NAND2_X1 U573 ( .A1(n505), .A2(n514), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n506), .ZN(G1336GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n509) );
  NAND2_X1 U576 ( .A1(n514), .A2(n507), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(n510), .ZN(G1337GAT) );
  NAND2_X1 U579 ( .A1(n514), .A2(n511), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U581 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(KEYINPUT44), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  XOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT113), .Z(n523) );
  NOR2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n519), .A2(n536), .ZN(n520) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n533), .A2(n548), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT114), .Z(n526) );
  NAND2_X1 U591 ( .A1(n533), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n530) );
  NAND2_X1 U596 ( .A1(n533), .A2(n558), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U598 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  XOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NOR2_X1 U603 ( .A1(n564), .A2(n545), .ZN(n538) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n538), .Z(G1344GAT) );
  NOR2_X1 U605 ( .A1(n545), .A2(n555), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n540) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  NOR2_X1 U610 ( .A1(n573), .A2(n545), .ZN(n543) );
  XOR2_X1 U611 ( .A(KEYINPUT118), .B(n543), .Z(n544) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n547), .Z(G1347GAT) );
  INV_X1 U615 ( .A(n554), .ZN(n559) );
  AND2_X1 U616 ( .A1(n559), .A2(n548), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n553) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n552) );
  XNOR2_X1 U622 ( .A(n553), .B(n552), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(n557), .B(n556), .Z(G1349GAT) );
  XOR2_X1 U625 ( .A(G183GAT), .B(KEYINPUT123), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n575) );
  NOR2_X1 U629 ( .A1(n564), .A2(n575), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U633 ( .A1(n575), .A2(n568), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

