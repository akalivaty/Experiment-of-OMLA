//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT69), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT69), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G953), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G227), .ZN(new_n198));
  XOR2_X1   g012(.A(G110), .B(G140), .Z(new_n199));
  XOR2_X1   g013(.A(new_n198), .B(new_n199), .Z(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n206), .B2(G146), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n204), .A2(KEYINPUT64), .A3(G143), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n208), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT10), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT84), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G104), .ZN(new_n224));
  INV_X1    g038(.A(G104), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT84), .A3(G107), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n225), .A2(G107), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(KEYINPUT83), .B(KEYINPUT3), .C1(new_n225), .C2(G107), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n227), .A2(new_n228), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n223), .A2(G104), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n205), .A2(new_n207), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n202), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n234), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n221), .A2(new_n237), .B1(new_n242), .B2(new_n220), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n205), .A2(new_n207), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n212), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n233), .A2(new_n226), .A3(new_n224), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n252));
  OR2_X1    g066(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n223), .A2(G104), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n250), .B(G101), .C1(new_n251), .C2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n257), .B(G101), .C1(new_n251), .C2(new_n255), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n234), .A3(KEYINPUT4), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n232), .A2(new_n233), .A3(new_n226), .A4(new_n224), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n260), .B2(G101), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n249), .B(new_n256), .C1(new_n259), .C2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G134), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n267), .B2(KEYINPUT11), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT11), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n265), .B(new_n269), .C1(new_n266), .C2(G137), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(KEYINPUT11), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n266), .A2(G137), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n270), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n243), .A2(new_n262), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT64), .B1(new_n204), .B2(G143), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n209), .A2(new_n206), .A3(G146), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n280), .A2(new_n281), .B1(G143), .B2(new_n204), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n213), .A2(new_n215), .B1(new_n205), .B2(KEYINPUT1), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n238), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n242), .B1(new_n237), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n285), .A2(KEYINPUT12), .A3(new_n277), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT12), .B1(new_n285), .B2(new_n277), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n279), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n279), .A2(new_n200), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n243), .A2(new_n262), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n277), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n201), .A2(new_n288), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n192), .B1(new_n292), .B2(G469), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n279), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n201), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n279), .B(new_n200), .C1(new_n286), .C2(new_n287), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT73), .B(G902), .Z(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n190), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n189), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT20), .ZN(new_n302));
  INV_X1    g116(.A(G237), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n206), .A2(KEYINPUT90), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n197), .A2(G214), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n194), .A2(new_n196), .A3(G214), .A4(new_n303), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT90), .A3(new_n206), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G131), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n307), .A3(new_n274), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(G125), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  INV_X1    g127(.A(G140), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(G125), .A2(G140), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(new_n312), .B2(G140), .ZN(new_n317));
  OAI211_X1 g131(.A(G146), .B(new_n315), .C1(new_n317), .C2(new_n313), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n320));
  AOI22_X1  g134(.A1(new_n317), .A2(KEYINPUT19), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n204), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n311), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n305), .A2(new_n307), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n308), .A2(KEYINPUT18), .A3(G131), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n204), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n327), .A2(KEYINPUT91), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT91), .B1(new_n327), .B2(new_n328), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n325), .B(new_n326), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n323), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G113), .B(G122), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n225), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT17), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n309), .A2(new_n337), .A3(new_n310), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n308), .A2(KEYINPUT17), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n318), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n313), .A2(new_n314), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT75), .A2(G125), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT75), .A2(G125), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(KEYINPUT75), .A2(G125), .ZN(new_n348));
  OAI21_X1  g162(.A(G140), .B1(new_n348), .B2(new_n344), .ZN(new_n349));
  INV_X1    g163(.A(new_n316), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n347), .B1(new_n351), .B2(KEYINPUT16), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT76), .A3(G146), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n313), .B1(new_n349), .B2(new_n350), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n204), .B1(new_n354), .B2(new_n347), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n342), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n334), .B(new_n331), .C1(new_n340), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n336), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G475), .A2(G902), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n302), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n302), .A3(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(new_n357), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n355), .B1(new_n318), .B2(new_n341), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT76), .B1(new_n352), .B2(G146), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n338), .A3(new_n339), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n334), .B1(new_n367), .B2(new_n331), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n191), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n361), .A2(new_n362), .B1(G475), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n197), .ZN(new_n371));
  INV_X1    g185(.A(new_n298), .ZN(new_n372));
  NAND2_X1  g186(.A1(G234), .A2(G237), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT21), .B(G898), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n373), .A2(G952), .A3(new_n193), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n206), .A2(G128), .ZN(new_n380));
  XOR2_X1   g194(.A(new_n380), .B(KEYINPUT13), .Z(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT66), .B(G128), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G143), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G134), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n266), .A3(new_n380), .ZN(new_n386));
  XNOR2_X1  g200(.A(G116), .B(G122), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(new_n223), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n390));
  INV_X1    g204(.A(G116), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n391), .B2(G122), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n390), .B1(new_n391), .B2(G122), .ZN(new_n394));
  OAI21_X1  g208(.A(G107), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n387), .A2(new_n223), .ZN(new_n398));
  INV_X1    g212(.A(new_n386), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n266), .B1(new_n383), .B2(new_n380), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n389), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G217), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n187), .A2(new_n403), .A3(G953), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(KEYINPUT94), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n405), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n389), .C1(new_n397), .C2(new_n401), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n298), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G478), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  OAI221_X1 g227(.A(new_n298), .B1(KEYINPUT15), .B2(new_n411), .C1(new_n406), .C2(new_n409), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n370), .A2(new_n379), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n301), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G214), .B1(G237), .B2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  XOR2_X1   g234(.A(KEYINPUT2), .B(G113), .Z(new_n421));
  XNOR2_X1  g235(.A(G116), .B(G119), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT2), .B(G113), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n391), .A2(G119), .ZN(new_n425));
  INV_X1    g239(.A(G119), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G116), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n424), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n256), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n259), .B2(new_n261), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n430), .B(KEYINPUT86), .C1(new_n259), .C2(new_n261), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n422), .A2(KEYINPUT5), .ZN(new_n435));
  INV_X1    g249(.A(G113), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n425), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n438), .B1(new_n421), .B2(new_n422), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n234), .A3(new_n236), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n433), .A2(new_n434), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G110), .B(G122), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n433), .A2(new_n442), .A3(new_n434), .A4(new_n440), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n193), .A2(G224), .ZN(new_n447));
  INV_X1    g261(.A(new_n248), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n245), .B(new_n312), .C1(new_n282), .C2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n447), .B(new_n449), .C1(new_n219), .C2(new_n312), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n312), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n284), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n447), .B1(new_n453), .B2(new_n449), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(new_n456), .A3(new_n443), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n447), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n451), .B2(new_n454), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n449), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n459), .A3(new_n447), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n440), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n439), .A2(new_n234), .A3(KEYINPUT87), .A4(new_n236), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n465), .B(new_n466), .C1(new_n237), .C2(new_n439), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n442), .B(KEYINPUT8), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n461), .A2(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n445), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT88), .B1(new_n470), .B2(new_n191), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(G902), .C1(new_n469), .C2(new_n445), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n458), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT89), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n458), .B(new_n477), .C1(new_n471), .C2(new_n473), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n420), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n418), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n403), .B1(new_n298), .B2(G234), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT24), .B(G110), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT74), .B1(new_n426), .B2(G128), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n216), .B2(new_n426), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n382), .A2(KEYINPUT74), .A3(G119), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n382), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT23), .B1(new_n202), .B2(G119), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n426), .B2(G128), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(G110), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n364), .B2(new_n365), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n486), .A2(new_n487), .A3(new_n484), .ZN(new_n496));
  XNOR2_X1  g310(.A(KEYINPUT77), .B(G110), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AND4_X1   g313(.A1(new_n495), .A2(new_n499), .A3(new_n318), .A4(new_n328), .ZN(new_n500));
  INV_X1    g314(.A(new_n328), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n501), .B1(new_n352), .B2(G146), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n495), .B1(new_n502), .B2(new_n499), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n494), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT79), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT79), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n494), .B(new_n506), .C1(new_n500), .C2(new_n503), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n197), .A2(G221), .A3(G234), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G137), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n503), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n502), .A2(new_n495), .A3(new_n499), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n513), .A2(new_n514), .B1(new_n356), .B2(new_n493), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT80), .B1(new_n515), .B2(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n505), .A2(KEYINPUT80), .A3(new_n507), .A4(new_n511), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT25), .B1(new_n519), .B2(new_n298), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n521), .B(new_n372), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n483), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n483), .A2(G902), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n524), .B(KEYINPUT81), .Z(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n529), .B(KEYINPUT72), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  INV_X1    g347(.A(new_n276), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n274), .B1(new_n268), .B2(new_n270), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n249), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n266), .A2(G137), .ZN(new_n537));
  OAI21_X1  g351(.A(G131), .B1(new_n537), .B2(new_n264), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n284), .A2(new_n276), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n533), .B1(new_n540), .B2(new_n429), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n429), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n276), .A2(new_n538), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT68), .B1(new_n544), .B2(new_n219), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n284), .A2(new_n546), .A3(new_n276), .A4(new_n538), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n536), .A3(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(new_n429), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n543), .B1(new_n533), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n197), .A2(G210), .A3(new_n303), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT27), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT26), .B(G101), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n545), .A2(KEYINPUT30), .A3(new_n536), .A4(new_n547), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT67), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n540), .B2(new_n560), .ZN(new_n561));
  AOI211_X1 g375(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n536), .C2(new_n539), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n429), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT31), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(new_n550), .A4(new_n555), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n565), .A2(new_n566), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n557), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n550), .A3(new_n555), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT70), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT31), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n570), .B2(KEYINPUT31), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n532), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G472), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT29), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n543), .B(new_n577), .C1(new_n533), .C2(new_n550), .ZN(new_n578));
  INV_X1    g392(.A(new_n541), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n548), .B(new_n429), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(KEYINPUT28), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n555), .B(new_n578), .C1(new_n581), .C2(new_n577), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n563), .A2(new_n577), .A3(new_n550), .A4(new_n556), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n583), .A2(new_n298), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n576), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n551), .A2(new_n556), .ZN(new_n587));
  INV_X1    g401(.A(new_n558), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n276), .A2(new_n538), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n277), .A2(new_n249), .B1(new_n589), .B2(new_n284), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT67), .B1(new_n590), .B2(KEYINPUT30), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n540), .A2(new_n559), .A3(new_n560), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n549), .B1(new_n593), .B2(new_n429), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n594), .A2(KEYINPUT71), .A3(new_n564), .A4(new_n555), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n565), .A2(new_n566), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n570), .A2(KEYINPUT31), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT70), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT31), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n530), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n575), .B(new_n586), .C1(new_n602), .C2(KEYINPUT32), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n528), .A2(KEYINPUT82), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT82), .B1(new_n528), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n482), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n474), .A2(new_n475), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n458), .B(new_n476), .C1(new_n471), .C2(new_n473), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n419), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n369), .A2(G475), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n358), .A2(new_n302), .A3(new_n359), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(new_n614), .B2(new_n360), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n410), .A2(new_n411), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT96), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n402), .B2(new_n405), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n406), .A2(new_n409), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n402), .A2(new_n405), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n621), .A2(new_n617), .A3(KEYINPUT33), .A4(new_n408), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n298), .A2(G478), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n378), .B2(new_n376), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n420), .B1(new_n474), .B2(new_n475), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT95), .A3(new_n609), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n612), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n523), .A2(new_n526), .A3(new_n300), .ZN(new_n631));
  INV_X1    g445(.A(new_n530), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n569), .B2(new_n574), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n372), .B1(new_n597), .B2(new_n601), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n633), .B1(new_n634), .B2(new_n576), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  OAI211_X1 g453(.A(new_n613), .B(new_n415), .C1(new_n614), .C2(new_n360), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n379), .B(KEYINPUT97), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n612), .A2(new_n629), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n636), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  OAI21_X1  g461(.A(new_n298), .B1(new_n569), .B2(new_n574), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n602), .B1(G472), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n505), .A2(new_n507), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n511), .A2(KEYINPUT36), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n650), .B(new_n651), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n525), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n523), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n649), .A2(new_n481), .A3(new_n418), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AND3_X1   g471(.A1(new_n628), .A2(KEYINPUT95), .A3(new_n609), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT95), .B1(new_n628), .B2(new_n609), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n633), .A2(new_n531), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n597), .A2(new_n601), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n585), .B1(new_n662), .B2(new_n532), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n301), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n374), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n378), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n370), .A2(new_n665), .A3(new_n415), .A4(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n668), .ZN(new_n670));
  OAI21_X1  g484(.A(KEYINPUT98), .B1(new_n640), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n664), .A3(new_n654), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XNOR2_X1  g488(.A(new_n668), .B(KEYINPUT39), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n300), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n615), .A2(new_n415), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n419), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n654), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n594), .A2(new_n556), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n191), .B1(new_n580), .B2(new_n555), .ZN(new_n687));
  OAI21_X1  g501(.A(G472), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT99), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n661), .A2(new_n575), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n479), .A2(new_n480), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT38), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n684), .A2(new_n685), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n679), .A2(new_n693), .A3(new_n683), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G143), .ZN(G45));
  NOR2_X1   g512(.A1(new_n626), .A2(new_n670), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n660), .A2(new_n664), .A3(new_n654), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  AOI21_X1  g515(.A(new_n527), .B1(new_n661), .B2(new_n663), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n297), .A2(new_n298), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n188), .A3(new_n299), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n630), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND3_X1  g523(.A1(new_n644), .A2(new_n702), .A3(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR3_X1   g525(.A1(new_n658), .A2(new_n659), .A3(new_n705), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n417), .B1(new_n523), .B2(new_n653), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(KEYINPUT102), .A3(new_n603), .A4(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n603), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n612), .A2(new_n629), .A3(new_n706), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  NOR2_X1   g534(.A1(new_n680), .A2(new_n642), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n612), .A2(new_n629), .A3(new_n706), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n648), .A2(G472), .ZN(new_n723));
  OAI221_X1 g537(.A(new_n598), .B1(new_n555), .B2(new_n581), .C1(new_n567), .C2(new_n568), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n632), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n526), .A3(new_n523), .A4(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n722), .A2(new_n726), .A3(KEYINPUT103), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(KEYINPUT103), .B1(new_n722), .B2(new_n726), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  AND3_X1   g545(.A1(new_n654), .A2(new_n723), .A3(new_n725), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n712), .A2(new_n732), .A3(new_n699), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n661), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n633), .A2(KEYINPUT104), .A3(new_n531), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n737), .A3(new_n663), .ZN(new_n738));
  AND4_X1   g552(.A1(new_n419), .A2(new_n300), .A3(new_n479), .A4(new_n480), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n739), .A2(new_n699), .A3(KEYINPUT42), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n740), .A3(new_n528), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n528), .A2(new_n603), .A3(new_n699), .A4(new_n739), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NAND4_X1  g560(.A1(new_n528), .A2(new_n603), .A3(new_n672), .A4(new_n739), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  AOI21_X1  g562(.A(KEYINPUT43), .B1(new_n370), .B2(KEYINPUT106), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n370), .A2(new_n625), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n370), .B(new_n625), .C1(KEYINPUT106), .C2(KEYINPUT43), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n635), .A4(new_n654), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n692), .A2(new_n420), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n288), .A2(new_n201), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n289), .A2(new_n291), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n292), .A2(KEYINPUT45), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(G469), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n762), .A2(new_n763), .A3(KEYINPUT105), .A4(G469), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n192), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n299), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n188), .B(new_n675), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n754), .A2(new_n773), .A3(new_n755), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n753), .A2(new_n635), .A3(new_n654), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n757), .A2(new_n772), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  NAND3_X1  g593(.A1(new_n755), .A2(new_n527), .A3(new_n699), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n603), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n188), .B1(new_n769), .B2(new_n770), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(KEYINPUT47), .B(new_n188), .C1(new_n769), .C2(new_n770), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n719), .A2(new_n606), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n692), .A2(new_n419), .A3(new_n641), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT108), .ZN(new_n791));
  AOI211_X1 g605(.A(new_n420), .B(new_n642), .C1(new_n479), .C2(new_n480), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n626), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n626), .A2(new_n793), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n640), .A2(KEYINPUT109), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n640), .A2(KEYINPUT109), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n636), .B(new_n791), .C1(new_n794), .C2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n707), .A3(new_n710), .A4(new_n655), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT103), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n612), .A2(new_n629), .A3(new_n706), .A4(new_n721), .ZN(new_n802));
  INV_X1    g616(.A(new_n726), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n727), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n789), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n523), .A2(new_n300), .A3(new_n653), .A4(new_n668), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n660), .A2(new_n691), .A3(new_n807), .A4(new_n681), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n733), .A2(new_n673), .A3(new_n700), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n612), .A2(new_n629), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n523), .A2(new_n653), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n664), .C1(new_n672), .C2(new_n699), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n808), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n370), .A2(new_n416), .A3(new_n668), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n818), .B1(new_n523), .B2(new_n653), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n603), .A3(new_n300), .A4(new_n755), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n648), .A2(G472), .B1(new_n632), .B2(new_n724), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n739), .A3(new_n654), .A4(new_n699), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n747), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n744), .B2(new_n741), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n817), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n702), .A2(KEYINPUT82), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n528), .A2(new_n603), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT82), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n482), .B1(new_n714), .B2(new_n718), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n523), .A2(new_n526), .A3(new_n300), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n791), .A2(new_n649), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n626), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n692), .A2(new_n793), .A3(new_n419), .A4(new_n641), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n798), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n528), .A2(new_n603), .A3(new_n706), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n612), .A2(new_n629), .A3(new_n643), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n835), .A2(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n612), .A2(new_n629), .A3(new_n627), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n655), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n833), .A2(new_n824), .A3(new_n844), .A4(new_n730), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT111), .A3(KEYINPUT53), .A4(new_n817), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n789), .A2(new_n800), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n730), .A4(new_n824), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n845), .A2(KEYINPUT110), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n817), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n827), .A2(new_n847), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT112), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n827), .A2(new_n847), .ZN(new_n857));
  INV_X1    g671(.A(new_n851), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n817), .B1(new_n845), .B2(KEYINPUT110), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT112), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT54), .ZN(new_n863));
  INV_X1    g677(.A(new_n817), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n853), .B1(new_n864), .B2(new_n845), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n825), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(KEYINPUT54), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n738), .A2(new_n528), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n755), .A2(new_n377), .A3(new_n706), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n752), .B2(new_n751), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT48), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n869), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n870), .A2(new_n691), .A3(new_n527), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n836), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(G952), .A3(new_n193), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n869), .B2(new_n871), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n803), .A2(new_n377), .A3(new_n753), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n717), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n880), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n784), .A2(new_n786), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n704), .A2(new_n299), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n188), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n755), .B(new_n883), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT51), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n615), .A2(new_n625), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n732), .A2(new_n871), .B1(new_n876), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n706), .A2(new_n420), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n693), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n693), .B2(new_n892), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n880), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT50), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(KEYINPUT50), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n880), .C1(new_n893), .C2(new_n894), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n890), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n875), .B(new_n882), .C1(new_n888), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n903), .B(new_n890), .C1(new_n897), .C2(new_n899), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n902), .A2(new_n904), .A3(new_n887), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n856), .A2(new_n863), .A3(new_n868), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(G952), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n193), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n885), .B(KEYINPUT49), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n420), .A2(new_n912), .A3(new_n189), .A4(new_n750), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n527), .A2(new_n913), .A3(new_n691), .A4(new_n693), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(G75));
  NAND2_X1  g729(.A1(new_n371), .A2(new_n909), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT119), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n866), .A2(new_n372), .ZN(new_n920));
  OAI211_X1 g734(.A(KEYINPUT118), .B(new_n919), .C1(new_n920), .C2(new_n475), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n446), .A2(new_n457), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT117), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n455), .B(KEYINPUT55), .Z(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n925), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(G51));
  XNOR2_X1  g742(.A(new_n192), .B(KEYINPUT57), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n865), .A2(new_n825), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n855), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n867), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n297), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n866), .A2(new_n372), .A3(new_n766), .A4(new_n767), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n918), .B1(new_n933), .B2(new_n934), .ZN(G54));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n920), .A2(new_n358), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n358), .B1(new_n920), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n918), .B1(new_n937), .B2(new_n938), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  NOR2_X1   g755(.A1(new_n623), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n931), .B2(new_n867), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n917), .ZN(new_n944));
  INV_X1    g758(.A(new_n941), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n855), .B1(new_n857), .B2(new_n860), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n868), .B1(new_n946), .B2(new_n862), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n945), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n949), .B2(new_n623), .ZN(G63));
  OAI21_X1  g764(.A(new_n917), .B1(KEYINPUT121), .B2(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n930), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n955), .B2(new_n652), .ZN(new_n956));
  NAND2_X1  g770(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n517), .B(new_n518), .C1(new_n930), .C2(new_n954), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n956), .B2(new_n958), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  INV_X1    g775(.A(new_n375), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n193), .B1(new_n962), .B2(G224), .ZN(new_n963));
  INV_X1    g777(.A(new_n806), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n197), .ZN(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n923), .B1(new_n966), .B2(new_n371), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  XNOR2_X1  g782(.A(new_n593), .B(new_n321), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n812), .A2(new_n680), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n772), .A2(new_n869), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n778), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n815), .A2(new_n733), .ZN(new_n975));
  AND4_X1   g789(.A1(new_n745), .A2(new_n787), .A3(new_n747), .A4(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n371), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n197), .A2(G900), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n969), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT124), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n626), .B1(new_n796), .B2(new_n797), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n832), .A2(new_n675), .A3(new_n739), .A4(new_n981), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n787), .A2(new_n778), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n694), .A2(new_n696), .A3(new_n733), .A4(new_n815), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT62), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n984), .B2(KEYINPUT62), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT62), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n697), .A2(new_n975), .A3(KEYINPUT122), .A4(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n984), .B2(KEYINPUT62), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n980), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n987), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT62), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n990), .A2(new_n992), .ZN(new_n998));
  NAND4_X1  g812(.A1(new_n997), .A2(KEYINPUT124), .A3(new_n998), .A4(new_n983), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n371), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n979), .B1(new_n1000), .B2(new_n969), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n197), .B1(G227), .B2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1002), .B(KEYINPUT125), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G72));
  INV_X1    g818(.A(new_n686), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n994), .A2(new_n999), .A3(new_n806), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n594), .A2(new_n556), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1011), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT127), .Z(new_n1013));
  NOR2_X1   g827(.A1(new_n854), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n974), .A2(new_n976), .A3(new_n806), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1011), .B1(new_n1015), .B2(new_n1008), .ZN(new_n1016));
  NOR4_X1   g830(.A1(new_n1009), .A2(new_n1014), .A3(new_n918), .A4(new_n1016), .ZN(G57));
endmodule


