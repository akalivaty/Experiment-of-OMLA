//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  AND2_X1   g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  INV_X1    g0010(.A(G97), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n202), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n209), .B(new_n213), .C1(G87), .C2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G107), .A2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G50), .A2(G226), .ZN(new_n217));
  NAND4_X1  g0017(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n208), .B(new_n221), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT67), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G264), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G303), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n252), .B1(new_n253), .B2(new_n251), .C1(new_n255), .C2(new_n212), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT71), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n223), .A2(KEYINPUT71), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT5), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n270), .A2(new_n258), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G270), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G116), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n282), .A2(new_n222), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n277), .A2(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n278), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G283), .ZN(new_n286));
  INV_X1    g0086(.A(G20), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n286), .B(new_n287), .C1(G33), .C2(new_n211), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n282), .A2(new_n222), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(new_n287), .C2(G116), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n290), .A2(new_n291), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n281), .B1(new_n280), .B2(new_n285), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n276), .A2(new_n295), .A3(G169), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT21), .ZN(new_n297));
  AND4_X1   g0097(.A1(G179), .A2(new_n263), .A3(new_n273), .A4(new_n275), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n296), .A2(new_n297), .B1(new_n298), .B2(new_n295), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n295), .A2(G169), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT97), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT21), .A4(new_n276), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT97), .B1(new_n296), .B2(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n276), .A2(G200), .ZN(new_n304));
  INV_X1    g0104(.A(new_n295), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n276), .ZN(new_n307));
  AND4_X1   g0107(.A1(new_n299), .A2(new_n302), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT74), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n309), .A2(G20), .A3(G33), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT74), .B1(new_n287), .B2(new_n248), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G50), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n248), .A2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n316), .A2(new_n202), .B1(new_n287), .B2(G68), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n289), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT11), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n277), .A2(G20), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n321), .A2(new_n289), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(KEYINPUT12), .B1(new_n278), .B2(G68), .ZN(new_n324));
  OR3_X1    g0124(.A1(new_n278), .A2(KEYINPUT12), .A3(G68), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n277), .B1(G41), .B2(G45), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n271), .ZN(new_n330));
  INV_X1    g0130(.A(G226), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n254), .ZN(new_n332));
  INV_X1    g0132(.A(G232), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G1698), .ZN(new_n334));
  AND2_X1   g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NOR2_X1   g0135(.A1(KEYINPUT3), .A2(G33), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n332), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n330), .B1(new_n339), .B2(new_n262), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n258), .A2(new_n329), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT69), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n329), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(G238), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT81), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n340), .A2(KEYINPUT81), .A3(new_n345), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(KEYINPUT13), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT82), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n340), .A2(new_n345), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n348), .A2(new_n351), .A3(KEYINPUT13), .A4(new_n349), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n328), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n346), .A2(KEYINPUT13), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n353), .B1(new_n340), .B2(new_n345), .ZN(new_n359));
  OAI21_X1  g0159(.A(G169), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT14), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT14), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(G169), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n327), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n340), .A2(KEYINPUT81), .A3(new_n345), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT81), .B1(new_n340), .B2(new_n345), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n366), .A2(new_n367), .A3(new_n353), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT82), .B1(new_n346), .B2(KEYINPUT13), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n356), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G190), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n358), .A2(new_n359), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n327), .B1(G200), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n374), .A3(KEYINPUT83), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT83), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n306), .B1(new_n355), .B2(new_n356), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n326), .B(new_n319), .C1(new_n372), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n365), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT84), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT84), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n365), .A2(new_n375), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n343), .A2(new_n344), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G226), .ZN(new_n387));
  INV_X1    g0187(.A(new_n330), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G222), .A2(G1698), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n254), .A2(G223), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n251), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n335), .A2(new_n336), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n202), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT70), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n391), .A2(KEYINPUT70), .A3(new_n393), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n262), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n387), .B(new_n388), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n397), .A2(G179), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT72), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(KEYINPUT8), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT8), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n402), .A2(KEYINPUT72), .A3(G58), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(G58), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n402), .A2(KEYINPUT73), .A3(G58), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n316), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G150), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n312), .A2(new_n411), .B1(new_n287), .B2(new_n201), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n289), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n279), .A2(new_n313), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT75), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n283), .A2(new_n415), .A3(new_n278), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT75), .B1(new_n279), .B2(new_n289), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(new_n417), .A3(G50), .A4(new_n320), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G169), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n397), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n398), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n413), .A2(new_n418), .A3(KEYINPUT9), .A4(new_n414), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n423), .B(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n419), .A2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n396), .A2(new_n394), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(G190), .A3(new_n388), .A4(new_n387), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n397), .A2(G200), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT10), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n429), .A2(new_n430), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n423), .A2(new_n424), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n423), .A2(new_n424), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n435), .B1(new_n441), .B2(new_n427), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n422), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n386), .A2(G244), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n388), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n251), .A2(G238), .A3(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI221_X1 g0249(.A(new_n448), .B1(new_n449), .B2(new_n251), .C1(new_n255), .C2(new_n333), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n262), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(KEYINPUT76), .A3(new_n388), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n328), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n321), .A2(new_n289), .A3(new_n202), .ZN(new_n455));
  NOR2_X1   g0255(.A1(G20), .A2(G33), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT74), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n400), .A2(KEYINPUT8), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n405), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g0260(.A(KEYINPUT15), .B(G87), .Z(new_n461));
  AOI22_X1  g0261(.A1(new_n461), .A2(new_n315), .B1(G20), .B2(G77), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n283), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n455), .B(new_n463), .C1(new_n202), .C2(new_n279), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n420), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n454), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n465), .B1(new_n466), .B2(G200), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT77), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n469), .A2(KEYINPUT77), .B1(new_n306), .B2(new_n466), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT80), .B1(new_n443), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n468), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n464), .B1(new_n453), .B2(new_n378), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT77), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n476), .A2(new_n477), .B1(G190), .B2(new_n453), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n475), .B1(new_n478), .B2(new_n470), .ZN(new_n479));
  XNOR2_X1  g0279(.A(new_n432), .B(new_n436), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n422), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n385), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT87), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT16), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n249), .A2(new_n287), .A3(new_n250), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT7), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n287), .A4(new_n250), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n322), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G58), .B(G68), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G20), .ZN(new_n492));
  INV_X1    g0292(.A(G159), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n312), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n485), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT7), .B1(new_n392), .B2(new_n287), .ZN(new_n496));
  INV_X1    g0296(.A(new_n489), .ZN(new_n497));
  OAI21_X1  g0297(.A(G68), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n457), .A2(G159), .B1(new_n491), .B2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(KEYINPUT16), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(new_n500), .A3(new_n289), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT85), .A4(new_n289), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n407), .B(new_n408), .C1(new_n401), .C2(new_n403), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n416), .A3(new_n417), .A4(new_n320), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n404), .A2(new_n409), .A3(new_n279), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT86), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n331), .A2(G1698), .ZN(new_n515));
  OAI221_X1 g0315(.A(new_n515), .B1(G223), .B2(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G87), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n516), .A2(new_n517), .B1(new_n260), .B2(new_n261), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n341), .A2(new_n333), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n518), .A2(new_n519), .A3(new_n330), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n306), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(G200), .B2(new_n520), .ZN(new_n522));
  AND4_X1   g0322(.A1(KEYINPUT17), .A2(new_n505), .A3(new_n514), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n513), .B1(new_n503), .B2(new_n504), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT17), .B1(new_n524), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n484), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n505), .A2(new_n514), .A3(new_n522), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(KEYINPUT17), .A3(new_n522), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(KEYINPUT87), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n505), .A2(new_n514), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n518), .A2(new_n330), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n533), .B2(new_n519), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n520), .A2(G179), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT18), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n524), .B2(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n526), .A2(new_n531), .A3(new_n541), .ZN(new_n542));
  XOR2_X1   g0342(.A(new_n542), .B(KEYINPUT88), .Z(new_n543));
  NAND2_X1  g0343(.A1(new_n483), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n254), .C1(new_n335), .C2(new_n336), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n248), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n262), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT99), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n274), .A2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n549), .A2(KEYINPUT99), .A3(new_n262), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n552), .A2(new_n273), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n553), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n272), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n555), .A2(G190), .B1(new_n557), .B2(G200), .ZN(new_n558));
  INV_X1    g0358(.A(new_n285), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n278), .A2(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n561), .B(KEYINPUT25), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n287), .B(G87), .C1(new_n335), .C2(new_n336), .ZN(new_n563));
  OAI21_X1  g0363(.A(KEYINPUT22), .B1(new_n563), .B2(KEYINPUT98), .ZN(new_n564));
  AOI21_X1  g0364(.A(G20), .B1(new_n249), .B2(new_n250), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT98), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(G87), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n315), .A2(G116), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n287), .A2(G107), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT23), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT24), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n569), .A2(KEYINPUT24), .A3(new_n570), .A4(new_n572), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n289), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n558), .A2(new_n560), .A3(new_n562), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n560), .A3(new_n562), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n555), .A2(G169), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n557), .A2(G179), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n210), .A2(G1698), .ZN(new_n584));
  OAI221_X1 g0384(.A(new_n584), .B1(G238), .B2(G1698), .C1(new_n335), .C2(new_n336), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n248), .B2(new_n280), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n262), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n277), .A2(G45), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n258), .A2(G250), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n265), .A2(G274), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT95), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(KEYINPUT95), .A3(new_n590), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n587), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n461), .A2(new_n278), .ZN(new_n596));
  INV_X1    g0396(.A(G87), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n285), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g0398(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n599));
  NAND2_X1  g0399(.A1(new_n338), .A2(new_n287), .ZN(new_n600));
  NOR2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n597), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n565), .A2(G68), .ZN(new_n604));
  XNOR2_X1  g0404(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n316), .B2(new_n211), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n596), .B(new_n598), .C1(new_n289), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n589), .A2(new_n590), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT95), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n592), .B1(new_n586), .B2(new_n262), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n595), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n607), .A2(new_n289), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n559), .A2(new_n461), .ZN(new_n616));
  INV_X1    g0416(.A(new_n596), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n587), .B(new_n328), .C1(new_n591), .C2(new_n593), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(G169), .C2(new_n612), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n578), .A2(new_n583), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n279), .A2(new_n211), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n285), .B2(new_n211), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n449), .B1(new_n488), .B2(new_n489), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n312), .A2(new_n202), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n625), .A2(KEYINPUT91), .B1(new_n626), .B2(KEYINPUT89), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n626), .A2(KEYINPUT89), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT6), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n211), .A2(new_n449), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n629), .B1(new_n630), .B2(new_n601), .ZN(new_n631));
  NAND2_X1  g0431(.A1(KEYINPUT6), .A2(G97), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT90), .B1(new_n632), .B2(G107), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n632), .A2(KEYINPUT90), .A3(G107), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G20), .ZN(new_n636));
  OAI21_X1  g0436(.A(G107), .B1(new_n496), .B2(new_n497), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT91), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n627), .A2(new_n628), .A3(new_n636), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n624), .B1(new_n640), .B2(new_n289), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n272), .B1(new_n274), .B2(G257), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT93), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n251), .A2(G244), .A3(new_n254), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT4), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n644), .A2(new_n286), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT94), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT94), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n251), .A2(new_n651), .A3(G250), .A4(G1698), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n643), .A2(KEYINPUT93), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n648), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n262), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n642), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G169), .ZN(new_n658));
  OAI211_X1 g0458(.A(G179), .B(new_n642), .C1(new_n655), .C2(new_n656), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n641), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT92), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n636), .B1(new_n625), .B2(KEYINPUT91), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT91), .B(G107), .C1(new_n496), .C2(new_n497), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n457), .A2(KEYINPUT89), .A3(G77), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n283), .B1(new_n666), .B2(new_n628), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n661), .B1(new_n667), .B2(new_n624), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n641), .A2(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n642), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n650), .A2(new_n652), .ZN(new_n672));
  INV_X1    g0472(.A(new_n654), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n643), .A2(KEYINPUT93), .B1(G33), .B2(G283), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n647), .A4(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n675), .B2(new_n262), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n306), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(G200), .B2(new_n676), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n660), .B1(new_n670), .B2(new_n678), .ZN(new_n679));
  AND4_X1   g0479(.A1(new_n308), .A2(new_n545), .A3(new_n622), .A4(new_n679), .ZN(G372));
  NOR2_X1   g0480(.A1(new_n641), .A2(KEYINPUT92), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n661), .B(new_n624), .C1(new_n640), .C2(new_n289), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT26), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n659), .B1(new_n676), .B2(new_n420), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n683), .A2(new_n684), .A3(new_n621), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n657), .A2(G190), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n676), .A2(G200), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n681), .A2(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n641), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n689), .A2(new_n578), .A3(new_n614), .A4(new_n691), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n299), .A2(new_n583), .A3(new_n303), .A4(new_n302), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n620), .B(new_n686), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n660), .A2(new_n621), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n684), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n545), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n422), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n371), .A2(new_n374), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n475), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n365), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n526), .A3(new_n531), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n541), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n704), .B2(new_n480), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(G369));
  INV_X1    g0506(.A(new_n308), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n708));
  INV_X1    g0508(.A(G13), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OR3_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .A3(G1), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT27), .B1(new_n711), .B2(G1), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n305), .A2(new_n717), .ZN(new_n718));
  MUX2_X1   g0518(.A(new_n707), .B(new_n708), .S(new_n718), .Z(new_n719));
  INV_X1    g0519(.A(G330), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n578), .A2(new_n583), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n579), .A2(new_n716), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n579), .A2(new_n582), .A3(new_n716), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n708), .A2(new_n716), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n579), .A2(new_n582), .A3(new_n717), .ZN(new_n730));
  INV_X1    g0530(.A(new_n722), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(G399));
  NOR2_X1   g0533(.A1(new_n602), .A2(G116), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n206), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n735), .A2(new_n737), .A3(new_n277), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n740));
  INV_X1    g0540(.A(new_n737), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n740), .C1(new_n226), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT101), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  AND4_X1   g0545(.A1(new_n684), .A2(new_n621), .A3(new_n685), .A4(new_n690), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n668), .A2(new_n621), .A3(new_n685), .A4(new_n669), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(KEYINPUT26), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n748), .B(new_n620), .C1(new_n693), .C2(new_n692), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n745), .B1(new_n749), .B2(new_n717), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n745), .B(new_n717), .C1(new_n694), .C2(new_n696), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n679), .A2(new_n308), .A3(new_n622), .A4(new_n717), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n594), .A2(new_n556), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n676), .A2(new_n298), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n676), .A2(new_n298), .A3(KEYINPUT30), .A4(new_n756), .ZN(new_n760));
  INV_X1    g0560(.A(new_n557), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n657), .A2(new_n328), .A3(new_n276), .A4(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n759), .B(new_n760), .C1(new_n612), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n716), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n755), .A2(KEYINPUT31), .A3(new_n764), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n764), .A2(KEYINPUT31), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n765), .A2(G330), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n754), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n744), .B1(new_n770), .B2(G1), .ZN(G364));
  INV_X1    g0571(.A(new_n721), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n277), .B1(new_n710), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n737), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n719), .A2(new_n720), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n772), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n719), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n227), .A2(new_n264), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n736), .A2(new_n251), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(new_n240), .C2(new_n264), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n251), .A2(new_n206), .ZN(new_n786));
  XOR2_X1   g0586(.A(G355), .B(KEYINPUT102), .Z(new_n787));
  OAI221_X1 g0587(.A(new_n785), .B1(G116), .B2(new_n206), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(KEYINPUT103), .A2(G169), .ZN(new_n789));
  NAND2_X1  g0589(.A1(KEYINPUT103), .A2(G169), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(G20), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n223), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT104), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n781), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n287), .A2(G179), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n799), .A2(new_n306), .A3(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n449), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n799), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n392), .B(new_n801), .C1(G87), .C2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT106), .Z(new_n805));
  AND3_X1   g0605(.A1(new_n328), .A2(new_n378), .A3(KEYINPUT105), .ZN(new_n806));
  AOI21_X1  g0606(.A(KEYINPUT105), .B1(new_n328), .B2(new_n378), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n287), .B1(new_n809), .B2(G190), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G97), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n287), .A2(new_n328), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n813), .A2(new_n306), .A3(new_n378), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n808), .A2(new_n287), .A3(G190), .ZN(new_n815));
  AOI21_X1  g0615(.A(KEYINPUT32), .B1(new_n815), .B2(G159), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n815), .A2(KEYINPUT32), .A3(G159), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n812), .B1(new_n202), .B2(new_n814), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n813), .A2(G190), .A3(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n813), .A2(new_n306), .A3(G200), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G50), .A2(new_n820), .B1(new_n822), .B2(G68), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n813), .A2(G190), .A3(new_n378), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n400), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n805), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n251), .B1(new_n827), .B2(G322), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n253), .B2(new_n802), .C1(new_n829), .C2(new_n814), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n815), .A2(G329), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n820), .A2(G326), .B1(new_n822), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n548), .C2(new_n810), .ZN(new_n834));
  INV_X1    g0634(.A(new_n800), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n830), .B(new_n834), .C1(G283), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n796), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n782), .A2(new_n798), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n778), .B1(new_n776), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT107), .ZN(G396));
  OAI211_X1 g0640(.A(new_n479), .B(new_n717), .C1(new_n694), .C2(new_n696), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n697), .A2(new_n717), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n468), .A2(new_n716), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n471), .A2(new_n472), .B1(new_n464), .B2(new_n717), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(new_n468), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(new_n768), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n768), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n776), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n843), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n478), .A2(new_n470), .B1(new_n465), .B2(new_n716), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n475), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n779), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G143), .A2(new_n827), .B1(new_n822), .B2(G150), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n820), .A2(G137), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n493), .C2(new_n814), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT34), .Z(new_n857));
  AOI21_X1  g0657(.A(new_n392), .B1(new_n811), .B2(G58), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n803), .A2(G50), .B1(new_n835), .B2(G68), .ZN(new_n859));
  INV_X1    g0659(.A(G132), .ZN(new_n860));
  INV_X1    g0660(.A(new_n815), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n821), .A2(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n392), .B1(new_n814), .B2(new_n280), .C1(new_n548), .C2(new_n824), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(G107), .B2(new_n803), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n815), .A2(G311), .ZN(new_n867));
  AOI22_X1  g0667(.A1(G303), .A2(new_n820), .B1(new_n835), .B2(G87), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n866), .A2(new_n812), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI22_X1  g0669(.A1(new_n857), .A2(new_n862), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n796), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n796), .A2(new_n779), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n202), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n853), .A2(new_n775), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n849), .A2(new_n874), .ZN(G384));
  AND2_X1   g0675(.A1(new_n765), .A2(new_n766), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n327), .A2(new_n716), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n381), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n365), .A2(new_n700), .A3(new_n877), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT108), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT108), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n876), .A2(new_n845), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n509), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n714), .B1(new_n501), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n542), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n527), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n505), .A2(new_n514), .B1(new_n536), .B2(new_n714), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT37), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n501), .A2(new_n886), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n887), .B1(new_n537), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n894), .B2(new_n527), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  INV_X1    g0698(.A(new_n890), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n892), .B1(new_n899), .B2(new_n527), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(new_n891), .ZN(new_n901));
  INV_X1    g0701(.A(new_n714), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n532), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n523), .A2(new_n525), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n903), .B1(new_n904), .B2(new_n541), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n898), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT40), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n885), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n888), .B2(new_n896), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(KEYINPUT110), .B(new_n911), .C1(new_n885), .C2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n888), .A2(new_n896), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n898), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n897), .ZN(new_n919));
  AND3_X1   g0719(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n883), .B1(new_n879), .B2(new_n880), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n921), .A3(new_n852), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n919), .A2(new_n876), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT110), .B1(new_n923), .B2(new_n911), .ZN(new_n924));
  OAI211_X1 g0724(.A(G330), .B(new_n910), .C1(new_n916), .C2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n483), .A2(new_n543), .A3(new_n767), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n911), .B1(new_n885), .B2(new_n914), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n909), .B1(new_n930), .B2(new_n915), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n545), .A3(new_n876), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n897), .A2(new_n934), .A3(new_n906), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT109), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n897), .A2(new_n938), .A3(new_n906), .A4(new_n934), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n365), .A2(new_n716), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n541), .A2(new_n902), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n882), .A2(new_n884), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n850), .B2(new_n841), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n944), .B1(new_n946), .B2(new_n919), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n933), .B(new_n948), .Z(new_n949));
  INV_X1    g0749(.A(new_n752), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n543), .B(new_n483), .C1(new_n950), .C2(new_n750), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n705), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n949), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n277), .B2(new_n710), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n280), .B1(new_n635), .B2(KEYINPUT35), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n955), .B(new_n225), .C1(KEYINPUT35), .C2(new_n635), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  OAI21_X1  g0757(.A(G77), .B1(new_n400), .B2(new_n322), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n958), .A2(new_n226), .B1(G50), .B2(new_n322), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n959), .A2(G1), .A3(new_n709), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n957), .A3(new_n960), .ZN(G367));
  INV_X1    g0761(.A(new_n679), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n732), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n679), .B1(new_n670), .B2(new_n717), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n683), .A2(new_n685), .A3(new_n716), .ZN(new_n966));
  AND2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n691), .B1(new_n967), .B2(new_n583), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n717), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n608), .A2(new_n717), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n621), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n620), .B2(new_n971), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT43), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n976));
  OR3_X1    g0776(.A1(new_n970), .A2(KEYINPUT43), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(KEYINPUT111), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n729), .B2(new_n967), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n732), .A2(new_n730), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n967), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n981), .A3(new_n967), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT44), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n985), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n987), .A2(new_n988), .A3(new_n983), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n982), .A2(new_n967), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n729), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n732), .A2(new_n728), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT113), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n721), .B1(KEYINPUT113), .B2(new_n995), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n769), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n737), .B(KEYINPUT41), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n773), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n729), .A2(new_n967), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n976), .A2(new_n1003), .A3(new_n977), .A4(new_n978), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n980), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(G303), .A2(new_n827), .B1(new_n820), .B2(G311), .ZN(new_n1006));
  INV_X1    g0806(.A(G317), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n810), .B2(new_n449), .C1(new_n1007), .C2(new_n861), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n802), .A2(new_n280), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(KEYINPUT46), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G97), .B2(new_n835), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n251), .B1(new_n1009), .B2(KEYINPUT46), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(new_n548), .C2(new_n821), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n814), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1008), .B(new_n1013), .C1(G283), .C2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n1014), .B1(new_n827), .B2(G150), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G143), .A2(new_n820), .B1(new_n803), .B2(G58), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n800), .A2(new_n202), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n392), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT114), .B(G137), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n815), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n322), .B2(new_n810), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1020), .B(new_n1023), .C1(G159), .C2(new_n822), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n796), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n781), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n973), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n461), .A2(new_n736), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n784), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n797), .B(new_n1030), .C1(new_n235), .C2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n775), .A3(new_n1029), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1005), .A2(new_n1033), .ZN(G387));
  OR2_X1    g0834(.A1(new_n770), .A2(new_n998), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n770), .A2(new_n998), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n737), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n784), .B1(new_n232), .B2(new_n264), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n786), .A2(new_n734), .ZN(new_n1039));
  AOI211_X1 g0839(.A(G45), .B(new_n735), .C1(G68), .C2(G77), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n459), .A2(new_n313), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT50), .Z(new_n1042));
  AOI22_X1  g0842(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n206), .A2(G107), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n797), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n726), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1045), .B1(new_n1046), .B2(new_n1028), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n819), .A2(KEYINPUT115), .A3(new_n493), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT115), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n820), .B2(G159), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1048), .B(new_n1050), .C1(G77), .C2(new_n803), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n811), .A2(new_n461), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n827), .A2(G50), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n251), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n506), .A2(new_n822), .B1(new_n1014), .B2(G68), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT116), .Z(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n211), .B2(new_n800), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1054), .B(new_n1057), .C1(G150), .C2(new_n815), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT117), .Z(new_n1059));
  OAI22_X1  g0859(.A1(new_n824), .A2(new_n1007), .B1(new_n814), .B2(new_n253), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT118), .Z(new_n1061));
  INV_X1    g0861(.A(G322), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1061), .B1(new_n829), .B2(new_n821), .C1(new_n1062), .C2(new_n819), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT119), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT48), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n863), .B2(new_n810), .C1(new_n548), .C2(new_n802), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT49), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n815), .A2(G326), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1068), .B(new_n392), .C1(new_n280), .C2(new_n800), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1059), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1047), .B1(new_n1070), .B2(new_n796), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n1071), .A2(new_n775), .B1(new_n774), .B2(new_n998), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1037), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT120), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1037), .A2(KEYINPUT120), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n1076), .ZN(G393));
  NOR2_X1   g0877(.A1(new_n993), .A2(new_n994), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n729), .B1(new_n990), .B2(new_n992), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1036), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n993), .A2(new_n770), .A3(new_n998), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n737), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n776), .B1(new_n967), .B2(new_n781), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n797), .B1(new_n211), .B2(new_n206), .C1(new_n245), .C2(new_n1031), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n824), .A2(new_n829), .B1(new_n819), .B2(new_n1007), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT52), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1085), .A2(new_n1086), .B1(G294), .B2(new_n1014), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n251), .B(new_n801), .C1(G283), .C2(new_n803), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n1089), .B1(new_n280), .B2(new_n810), .C1(new_n1062), .C2(new_n861), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(G303), .C2(new_n822), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1014), .A2(new_n459), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n824), .A2(new_n493), .B1(new_n819), .B2(new_n411), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT51), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1092), .B1(new_n313), .B2(new_n821), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n811), .A2(G77), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n392), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n803), .A2(G68), .B1(new_n835), .B2(G87), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1095), .B(new_n1099), .C1(G143), .C2(new_n815), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n796), .B1(new_n1091), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1083), .A2(new_n1084), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n774), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1082), .A2(new_n1104), .ZN(G390));
  AOI21_X1  g0905(.A(new_n942), .B1(new_n897), .B2(new_n906), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n749), .A2(new_n479), .A3(new_n717), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1107), .A2(new_n850), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1106), .B1(new_n1108), .B2(new_n945), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n841), .A2(new_n850), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n920), .A2(new_n921), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n942), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1109), .B1(new_n940), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n767), .A3(new_n845), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1109), .B(new_n1114), .C1(new_n940), .C2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n774), .A3(new_n1117), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n940), .A2(new_n780), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI22_X1  g0920(.A1(new_n822), .A2(new_n1021), .B1(new_n1014), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n810), .B2(new_n493), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT121), .ZN(new_n1123));
  INV_X1    g0923(.A(G125), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1123), .B(new_n251), .C1(new_n1124), .C2(new_n861), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(G128), .A2(new_n820), .B1(new_n827), .B2(G132), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n313), .B2(new_n800), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n803), .A2(G150), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1125), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n392), .B1(new_n802), .B2(new_n597), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT123), .Z(new_n1132));
  AOI22_X1  g0932(.A1(G116), .A2(new_n827), .B1(new_n835), .B2(G68), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G97), .A2(new_n1014), .B1(new_n822), .B2(G107), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1132), .B(new_n1133), .C1(KEYINPUT122), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT122), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1137), .B(new_n1096), .C1(new_n548), .C2(new_n861), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(G283), .C2(new_n820), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n796), .B1(new_n1130), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n872), .A2(new_n409), .A3(new_n404), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1119), .A2(new_n775), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1118), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT124), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n845), .A2(new_n765), .A3(G330), .A4(new_n766), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n945), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1114), .A2(new_n1108), .A3(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1110), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n922), .A2(new_n767), .B1(new_n945), .B2(new_n1147), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n951), .A2(new_n705), .A3(new_n926), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1146), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n951), .A2(new_n705), .A3(new_n926), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1114), .A2(new_n1148), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1110), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1158), .B2(new_n1149), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1116), .A2(new_n1159), .A3(new_n1117), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n737), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1118), .A2(KEYINPUT124), .A3(new_n1142), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1145), .A2(new_n1161), .A3(new_n1162), .ZN(G378));
  NAND2_X1  g0963(.A1(new_n419), .A2(new_n902), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n443), .B(new_n1164), .Z(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n776), .B1(new_n1167), .B2(new_n779), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n872), .A2(new_n313), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n796), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G116), .A2(new_n820), .B1(new_n1014), .B2(new_n461), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n827), .A2(G107), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1171), .A2(new_n266), .A3(new_n392), .A4(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G97), .A2(new_n822), .B1(new_n803), .B2(G77), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n810), .B2(new_n322), .C1(new_n863), .C2(new_n861), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(G58), .C2(new_n835), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT58), .Z(new_n1177));
  OAI21_X1  g0977(.A(new_n313), .B1(new_n335), .B2(G41), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n811), .A2(G150), .B1(new_n803), .B2(new_n1120), .ZN(new_n1179));
  INV_X1    g0979(.A(G128), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n824), .A2(new_n1180), .B1(new_n819), .B2(new_n1124), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(G137), .B2(new_n1014), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n860), .C2(new_n821), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT59), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n815), .A2(G124), .ZN(new_n1185));
  AOI21_X1  g0985(.A(G33), .B1(new_n835), .B2(G159), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1184), .A2(new_n266), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1177), .A2(new_n1178), .A3(new_n1187), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1168), .B(new_n1169), .C1(new_n1170), .C2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT125), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n948), .A2(new_n1167), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1165), .B(new_n1166), .Z(new_n1192));
  NAND3_X1  g0992(.A1(new_n943), .A2(new_n947), .A3(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1191), .A2(G330), .A3(new_n931), .A4(new_n1193), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n943), .A2(new_n947), .A3(new_n1192), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1192), .B1(new_n943), .B2(new_n947), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n925), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1194), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1190), .B1(new_n774), .B2(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1194), .A2(new_n1197), .B1(new_n1153), .B2(new_n1160), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n737), .B1(new_n1200), .B2(KEYINPUT57), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1160), .A2(new_n1153), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1199), .B1(new_n1201), .B2(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n945), .A2(new_n779), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n821), .A2(new_n280), .B1(new_n819), .B2(new_n548), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(G107), .B2(new_n1014), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT126), .Z(new_n1208));
  AOI211_X1 g1008(.A(new_n1018), .B(new_n1208), .C1(G97), .C2(new_n803), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n815), .A2(G303), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n811), .A2(new_n461), .B1(G283), .B2(new_n827), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1209), .A2(new_n392), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n811), .A2(G50), .B1(G128), .B2(new_n815), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n822), .A2(new_n1120), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n251), .B1(new_n814), .B2(new_n411), .C1(new_n860), .C2(new_n819), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G159), .B2(new_n803), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n827), .A2(new_n1021), .B1(new_n835), .B2(G58), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1170), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n776), .B(new_n1219), .C1(new_n322), .C2(new_n872), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1152), .A2(new_n774), .B1(new_n1205), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1000), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1221), .B1(new_n1222), .B2(new_n1159), .ZN(G381));
  NAND2_X1  g1023(.A1(new_n1198), .A2(new_n774), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT125), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1189), .B(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n925), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1191), .A2(new_n1193), .B1(new_n931), .B2(G330), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1202), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT57), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n741), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1227), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G378), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1236), .A2(G384), .A3(G381), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1005), .A2(new_n1082), .A3(new_n1104), .A4(new_n1033), .ZN(new_n1238));
  INV_X1    g1038(.A(G396), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1075), .A2(new_n1239), .A3(new_n1076), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(G407));
  OAI211_X1 g1042(.A(G407), .B(G213), .C1(G343), .C2(new_n1236), .ZN(G409));
  INV_X1    g1043(.A(G213), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1244), .A2(G343), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1000), .B(new_n1202), .C1(new_n1228), .C2(new_n1229), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1235), .A2(new_n1199), .A3(new_n1247), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1114), .A2(new_n1108), .A3(new_n1148), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1150), .B1(new_n1114), .B2(new_n1148), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT60), .B1(new_n1253), .B2(new_n1156), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1250), .B1(new_n1254), .B2(new_n1159), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(KEYINPUT60), .A3(new_n1156), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n737), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT60), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(KEYINPUT127), .A3(new_n1154), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1255), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1261), .A2(G384), .A3(new_n1221), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1261), .B2(new_n1221), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1245), .A2(G2897), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1259), .A2(KEYINPUT127), .A3(new_n1154), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1259), .B2(new_n1154), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1256), .A2(new_n737), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1221), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(G384), .A3(new_n1221), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1264), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1266), .A2(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT61), .B1(new_n1249), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(G375), .A2(G378), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1247), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1245), .B1(new_n1279), .B2(new_n1235), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1278), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT62), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1277), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G387), .A2(G390), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1238), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1240), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1286), .A2(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1278), .A2(new_n1280), .A3(new_n1282), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT63), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(new_n1249), .B2(new_n1276), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1297), .B(new_n1298), .C1(new_n1300), .C2(new_n1296), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1295), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(new_n1236), .A2(new_n1278), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1282), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1303), .A2(new_n1282), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1293), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1306), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1308), .A2(new_n1294), .A3(new_n1304), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(G402));
endmodule


