//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n218), .B2(new_n220), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT65), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n216), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n256));
  OAI21_X1  g0056(.A(G58), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT71), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT8), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT71), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(G58), .C1(new_n255), .C2(new_n256), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n254), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n253), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n210), .A2(G1), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n202), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n272), .A2(new_n274), .B1(new_n202), .B2(new_n271), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n264), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT67), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT69), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(G1698), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  OAI21_X1  g0092(.A(KEYINPUT69), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n279), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT68), .B(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G222), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n296), .A2(new_n297), .B1(new_n224), .B2(new_n289), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n278), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  AOI21_X1  g0101(.A(G1), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n278), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  INV_X1    g0104(.A(new_n216), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n303), .A2(G226), .B1(new_n307), .B2(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G179), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n277), .B(new_n310), .C1(new_n311), .C2(new_n309), .ZN(new_n312));
  XOR2_X1   g0112(.A(new_n277), .B(KEYINPUT9), .Z(new_n313));
  INV_X1    g0113(.A(new_n309), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G190), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n309), .A2(G200), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n313), .A2(new_n315), .A3(new_n319), .A4(new_n316), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n312), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n263), .A2(new_n270), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n273), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n262), .A2(new_n260), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT70), .B(KEYINPUT8), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n261), .B1(new_n326), .B2(G58), .ZN(new_n327));
  OAI211_X1 g0127(.A(KEYINPUT76), .B(new_n324), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n272), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT76), .B1(new_n263), .B2(new_n324), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n259), .A2(new_n222), .ZN(new_n332));
  OAI21_X1  g0132(.A(G20), .B1(new_n332), .B2(new_n201), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n267), .A2(G159), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n286), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n281), .A2(new_n282), .A3(new_n280), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT67), .B1(new_n285), .B2(new_n286), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n210), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n336), .B1(new_n343), .B2(new_n222), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n285), .A2(new_n210), .A3(new_n286), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n342), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n337), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n335), .B1(new_n349), .B2(G68), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n254), .B1(new_n350), .B2(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n331), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n281), .A2(new_n282), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G1698), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n356), .A3(G223), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G226), .A2(G1698), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n264), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n278), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n303), .A2(G232), .B1(new_n307), .B2(new_n302), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n362), .A2(G190), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n362), .B2(new_n363), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT17), .B1(new_n352), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(G20), .B1(new_n283), .B2(new_n287), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n337), .B1(new_n369), .B2(KEYINPUT7), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n335), .B1(new_n370), .B2(G68), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n351), .B1(new_n371), .B2(KEYINPUT16), .ZN(new_n372));
  INV_X1    g0172(.A(new_n272), .ZN(new_n373));
  INV_X1    g0173(.A(new_n260), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT70), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT8), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT70), .A2(KEYINPUT8), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n259), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n374), .B1(new_n379), .B2(new_n261), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n273), .B1(new_n380), .B2(new_n258), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n373), .B1(new_n381), .B2(KEYINPUT76), .ZN(new_n382));
  INV_X1    g0182(.A(new_n330), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n322), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n372), .A2(new_n384), .A3(new_n367), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n372), .A2(new_n384), .A3(new_n367), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n368), .B1(new_n389), .B2(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n372), .A2(new_n384), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n311), .B1(new_n362), .B2(new_n363), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n362), .A2(new_n363), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(G179), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n396), .B(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n390), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G13), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(G1), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT74), .A3(G20), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT74), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n270), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(new_n253), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(G77), .A3(new_n324), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n402), .A2(new_n404), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(G77), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT8), .B(G58), .ZN(new_n410));
  INV_X1    g0210(.A(new_n267), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n410), .A2(new_n411), .B1(new_n210), .B2(new_n224), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  INV_X1    g0213(.A(new_n265), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n253), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT73), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n409), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n223), .B1(new_n291), .B2(new_n293), .ZN(new_n419));
  INV_X1    g0219(.A(G232), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n296), .A2(new_n420), .B1(new_n206), .B2(new_n289), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n278), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n303), .A2(G244), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n307), .A2(new_n302), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n425), .B(KEYINPUT72), .Z(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G190), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n418), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n365), .B1(new_n422), .B2(new_n426), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n418), .B1(new_n427), .B2(new_n311), .ZN(new_n432));
  INV_X1    g0232(.A(G179), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n422), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n321), .A2(new_n399), .A3(new_n431), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n222), .A2(G20), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n437), .B1(new_n411), .B2(new_n202), .C1(new_n414), .C2(new_n224), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n253), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT11), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n406), .A2(G68), .A3(new_n324), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n401), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(KEYINPUT12), .A3(new_n437), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n405), .A2(new_n222), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(KEYINPUT12), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT14), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n303), .A2(G238), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n283), .A2(new_n287), .A3(G226), .A4(new_n295), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G97), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n283), .A2(new_n287), .A3(G232), .A4(G1698), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n305), .A2(new_n306), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n450), .B(new_n424), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT13), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n459), .A2(KEYINPUT13), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n449), .B(G169), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n450), .A2(new_n424), .ZN(new_n464));
  INV_X1    g0264(.A(new_n457), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n278), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT13), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G179), .A3(new_n460), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n460), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n449), .B1(new_n471), .B2(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n448), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n447), .B1(new_n471), .B2(new_n428), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n365), .B1(new_n468), .B2(new_n460), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n436), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT90), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT79), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G41), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n301), .A2(G1), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n300), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G264), .A3(new_n458), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT88), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT88), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n486), .A2(new_n489), .A3(new_n458), .A4(G264), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n285), .A2(new_n286), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n295), .ZN(new_n493));
  INV_X1    g0293(.A(G250), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(G257), .B(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n496));
  INV_X1    g0296(.A(G294), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n496), .B1(new_n264), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n278), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n486), .A2(new_n304), .A3(new_n278), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(G190), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n491), .A2(new_n499), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT89), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(new_n501), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n503), .B1(new_n508), .B2(new_n365), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n492), .A2(new_n210), .A3(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT22), .ZN(new_n511));
  OR3_X1    g0311(.A1(new_n360), .A2(KEYINPUT22), .A3(G20), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n288), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n514));
  XNOR2_X1  g0314(.A(new_n514), .B(KEYINPUT86), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(KEYINPUT87), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n515), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT87), .A4(new_n518), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n253), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n271), .A2(new_n206), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n527), .B(KEYINPUT25), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n209), .A2(G33), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n270), .A2(new_n529), .A3(new_n216), .A4(new_n252), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n206), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n480), .B1(new_n509), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT89), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT89), .B1(new_n491), .B2(new_n499), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n535), .A2(new_n536), .A3(new_n500), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n537), .A2(G200), .B1(G190), .B2(new_n502), .ZN(new_n538));
  INV_X1    g0338(.A(new_n532), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n525), .B2(new_n253), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(KEYINPUT90), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n502), .A2(G169), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n508), .B2(new_n433), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n533), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n492), .A2(new_n210), .A3(G68), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n210), .B1(new_n452), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G87), .B2(new_n207), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT80), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(new_n547), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n550), .B2(new_n547), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n546), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n253), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n402), .A2(new_n404), .A3(new_n413), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n557), .C1(new_n413), .C2(new_n530), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n492), .A2(G244), .A3(G1698), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G116), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n559), .B(new_n560), .C1(new_n493), .C2(new_n223), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n278), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n278), .A2(new_n494), .A3(new_n484), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n307), .B2(new_n484), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n433), .A3(new_n564), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n562), .A2(new_n564), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n558), .B(new_n565), .C1(new_n566), .C2(G169), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n530), .A2(new_n360), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n568), .B(new_n556), .C1(new_n554), .C2(new_n253), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(G190), .A3(new_n564), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n566), .C2(new_n365), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT4), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n225), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n283), .A2(new_n287), .A3(new_n295), .A4(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(G244), .B1(new_n281), .B2(new_n282), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n354), .A2(new_n356), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G283), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n288), .A2(new_n494), .A3(new_n292), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n278), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n486), .A2(new_n458), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n500), .B1(G257), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n311), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n582), .A2(new_n433), .A3(new_n584), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n271), .A2(KEYINPUT78), .A3(new_n205), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT78), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n270), .B2(G97), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n588), .B(new_n590), .C1(new_n205), .C2(new_n530), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n205), .A3(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n210), .B1(new_n224), .B2(new_n411), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n370), .B2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n592), .B1(new_n598), .B2(new_n254), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n586), .A2(new_n587), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n597), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n343), .B2(new_n206), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(new_n602), .B2(new_n253), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n585), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n428), .C2(new_n585), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n572), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n542), .A2(new_n545), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT83), .ZN(new_n609));
  AND2_X1   g0409(.A1(G264), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n281), .B2(new_n282), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT81), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n492), .A2(KEYINPUT81), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n288), .A2(G303), .ZN(new_n616));
  INV_X1    g0416(.A(G257), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n285), .B2(new_n286), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n295), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n288), .A2(G303), .B1(new_n295), .B2(new_n618), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT82), .A3(new_n615), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n458), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n500), .B1(G270), .B2(new_n583), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n609), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(KEYINPUT82), .A2(new_n615), .A3(new_n616), .A4(new_n619), .ZN(new_n629));
  AOI21_X1  g0429(.A(KEYINPUT82), .B1(new_n623), .B2(new_n615), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n278), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n631), .A2(KEYINPUT83), .A3(new_n626), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G200), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n579), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n635), .B(new_n253), .C1(new_n210), .C2(G116), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT20), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  INV_X1    g0439(.A(G116), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(new_n405), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n209), .B2(G33), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n406), .A2(KEYINPUT84), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT84), .B1(new_n406), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n628), .A2(G190), .A3(new_n632), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n634), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(G169), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n628), .B2(new_n632), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT21), .B1(new_n650), .B2(KEYINPUT85), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n645), .A2(G169), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n625), .A2(new_n609), .A3(new_n627), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT83), .B1(new_n631), .B2(new_n626), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT85), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT21), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n626), .A2(G179), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n645), .A2(new_n631), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n648), .A2(new_n651), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n608), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n479), .A2(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n435), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n471), .A2(G169), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT14), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n469), .A3(new_n463), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n477), .A2(new_n665), .B1(new_n668), .B2(new_n448), .ZN(new_n669));
  INV_X1    g0469(.A(new_n390), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n398), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n318), .A2(new_n320), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n312), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n436), .A2(new_n478), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n606), .B1(new_n534), .B2(new_n541), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n651), .A2(new_n658), .A3(new_n661), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n544), .A2(new_n533), .A3(KEYINPUT91), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT91), .B1(new_n544), .B2(new_n533), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n675), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n567), .A2(new_n571), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n600), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(new_n600), .A3(new_n681), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n567), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n673), .B1(new_n674), .B2(new_n690), .ZN(G369));
  OR3_X1    g0491(.A1(new_n443), .A2(KEYINPUT27), .A3(G20), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT27), .B1(new_n443), .B2(G20), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n676), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  OAI211_X1 g0499(.A(new_n542), .B(new_n545), .C1(new_n540), .C2(new_n697), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n537), .A2(G179), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n540), .B1(new_n701), .B2(new_n543), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n696), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n646), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n676), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n662), .B2(new_n706), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(G330), .A3(new_n704), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n679), .A2(new_n697), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n709), .A3(new_n710), .ZN(G399));
  INV_X1    g0511(.A(new_n213), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n220), .B2(new_n714), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n696), .B1(new_n680), .B2(new_n688), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n651), .A2(new_n658), .A3(new_n661), .A4(new_n545), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n675), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n681), .A2(KEYINPUT97), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n567), .B1(new_n683), .B2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT97), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n686), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n696), .B1(new_n723), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n506), .A2(new_n507), .A3(new_n566), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n631), .A2(new_n660), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n732), .B1(KEYINPUT94), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n631), .A2(new_n735), .A3(new_n660), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n585), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(KEYINPUT95), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT94), .B1(new_n625), .B2(new_n659), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n562), .A2(new_n564), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n535), .A2(new_n536), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n740), .A2(new_n736), .A3(new_n742), .A4(new_n738), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n739), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n585), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n740), .A2(new_n736), .A3(new_n742), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n585), .A2(new_n433), .A3(new_n741), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n537), .A2(new_n749), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n748), .A2(new_n737), .B1(new_n633), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n746), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(KEYINPUT96), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT96), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n746), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n753), .A2(new_n696), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT31), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n697), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n663), .A2(new_n697), .B1(new_n752), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n731), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n730), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n719), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR2_X1   g0563(.A1(new_n400), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n209), .B1(new_n764), .B2(G45), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n713), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n708), .B2(G330), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n708), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n216), .B1(G20), .B2(new_n311), .ZN(new_n770));
  OR2_X1    g0570(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(KEYINPUT98), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n210), .A2(new_n433), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n776), .A2(new_n428), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n776), .A2(new_n428), .A3(new_n365), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n778), .A2(new_n259), .B1(new_n780), .B2(new_n202), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n776), .A2(new_n365), .A3(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n775), .A2(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n783), .A2(new_n222), .B1(new_n785), .B2(new_n224), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n428), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n210), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n205), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n210), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n784), .ZN(new_n792));
  INV_X1    g0592(.A(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT32), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n790), .B(new_n796), .C1(G87), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n791), .A2(new_n428), .A3(G200), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT99), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G107), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n288), .B1(new_n795), .B2(new_n794), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n787), .A2(new_n799), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n785), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n779), .A2(G326), .B1(G311), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n789), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G294), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n806), .A2(new_n288), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n797), .B(KEYINPUT100), .Z(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G303), .B1(G283), .B2(new_n801), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n777), .A2(G322), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  INV_X1    g0613(.A(new_n792), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n782), .A2(new_n813), .B1(G329), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n809), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n774), .B1(new_n804), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G13), .A2(G33), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(G20), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n773), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n712), .A2(new_n492), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(G45), .B2(new_n220), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n250), .B2(G45), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n289), .A2(new_n213), .ZN(new_n825));
  INV_X1    g0625(.A(G355), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n825), .A2(new_n826), .B1(G116), .B2(new_n213), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n821), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n767), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n817), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n820), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n708), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n769), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NAND2_X1  g0634(.A1(new_n665), .A2(new_n697), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n429), .A2(new_n430), .B1(new_n418), .B2(new_n697), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n435), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n720), .A2(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n696), .B(new_n838), .C1(new_n680), .C2(new_n688), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n761), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n767), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n761), .A2(new_n840), .A3(new_n842), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n774), .A2(new_n819), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n767), .B1(new_n847), .B2(G77), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n780), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n783), .A2(new_n851), .B1(new_n785), .B2(new_n793), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n850), .B(new_n852), .C1(G143), .C2(new_n777), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT34), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n353), .B1(new_n814), .B2(G132), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n259), .C2(new_n789), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n801), .A2(G68), .ZN(new_n857));
  INV_X1    g0657(.A(new_n810), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n202), .B2(new_n858), .C1(new_n853), .C2(KEYINPUT34), .ZN(new_n859));
  OAI22_X1  g0659(.A1(new_n778), .A2(new_n497), .B1(new_n785), .B2(new_n640), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G311), .B2(new_n814), .ZN(new_n861));
  INV_X1    g0661(.A(new_n790), .ZN(new_n862));
  XNOR2_X1  g0662(.A(KEYINPUT101), .B(G283), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n864), .A2(new_n782), .B1(new_n779), .B2(G303), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n861), .A2(new_n288), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n801), .A2(G87), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n858), .B2(new_n206), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n856), .A2(new_n859), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n848), .B1(new_n869), .B2(new_n773), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n839), .B2(new_n819), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n846), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n764), .A2(new_n209), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n721), .A2(new_n729), .A3(new_n479), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n673), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n385), .B1(new_n352), .B2(new_n394), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n352), .A2(new_n694), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT37), .B1(new_n391), .B2(new_n395), .ZN(new_n882));
  INV_X1    g0682(.A(new_n694), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n391), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n882), .A2(new_n386), .A3(new_n388), .A4(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n881), .A2(new_n885), .A3(KEYINPUT102), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT102), .B1(new_n881), .B2(new_n885), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n390), .B2(new_n398), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n350), .A2(KEYINPUT16), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n892), .A2(new_n351), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n395), .B1(new_n893), .B2(new_n331), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n883), .B1(new_n893), .B2(new_n331), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n389), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n390), .B2(new_n398), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT38), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n878), .B1(new_n891), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n668), .A2(new_n448), .A3(new_n697), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT38), .B(new_n898), .C1(new_n399), .C2(new_n895), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT39), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n905), .A3(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n448), .B(new_n696), .C1(new_n668), .C2(new_n476), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n447), .A2(new_n697), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n473), .A2(new_n477), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n906), .A2(new_n907), .ZN(new_n915));
  INV_X1    g0715(.A(new_n835), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n915), .C1(new_n841), .C2(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n398), .A2(new_n883), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n909), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n877), .B(new_n919), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n889), .A2(new_n886), .A3(new_n887), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n907), .B1(new_n921), .B2(KEYINPUT38), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n838), .B1(new_n910), .B2(new_n913), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n746), .A2(new_n754), .A3(new_n751), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n754), .B1(new_n746), .B2(new_n751), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT31), .B1(new_n926), .B2(new_n696), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n753), .A2(new_n755), .A3(new_n759), .ZN(new_n928));
  INV_X1    g0728(.A(new_n662), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n702), .B(new_n606), .C1(new_n541), .C2(new_n534), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n929), .A2(new_n930), .A3(new_n697), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n922), .B(new_n923), .C1(new_n927), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT40), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n928), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n758), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT40), .B1(new_n906), .B2(new_n907), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n923), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n927), .A2(new_n932), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n940), .A2(new_n674), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n731), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n939), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n874), .B1(new_n920), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n920), .B2(new_n943), .ZN(new_n945));
  INV_X1    g0745(.A(new_n596), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n640), .B(new_n218), .C1(new_n946), .C2(KEYINPUT35), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT35), .B2(new_n946), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n220), .A2(new_n224), .A3(new_n332), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n222), .A2(G50), .ZN(new_n951));
  OAI211_X1 g0751(.A(G1), .B(new_n400), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n945), .A2(new_n949), .A3(new_n952), .ZN(G367));
  OAI211_X1 g0753(.A(new_n605), .B(new_n600), .C1(new_n603), .C2(new_n697), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n600), .A2(new_n697), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n699), .A2(new_n704), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT42), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n600), .B1(new_n954), .B2(new_n545), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n959), .A2(new_n960), .B1(new_n697), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n697), .A2(new_n569), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n687), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n682), .B2(new_n963), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT43), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT104), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n968), .A2(new_n969), .B1(new_n962), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(KEYINPUT104), .B1(new_n962), .B2(new_n967), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT105), .ZN(new_n974));
  INV_X1    g0774(.A(new_n956), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n709), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT105), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n977), .A3(new_n972), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n977), .B1(new_n971), .B2(new_n972), .ZN(new_n980));
  INV_X1    g0780(.A(new_n962), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n969), .A3(new_n966), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n962), .A2(new_n970), .ZN(new_n983));
  AND4_X1   g0783(.A1(new_n977), .A2(new_n982), .A3(new_n972), .A4(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n980), .A2(new_n984), .B1(new_n709), .B2(new_n975), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n713), .B(KEYINPUT41), .Z(new_n986));
  AOI21_X1  g0786(.A(new_n956), .B1(new_n705), .B2(new_n710), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n705), .A2(new_n710), .A3(new_n956), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n709), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n709), .ZN(new_n996));
  INV_X1    g0796(.A(new_n699), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n704), .B1(new_n708), .B2(G330), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n997), .B1(new_n996), .B2(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n990), .A2(new_n709), .A3(new_n993), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n995), .A2(new_n762), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n986), .B1(new_n1004), .B2(new_n762), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n979), .B(new_n985), .C1(new_n766), .C2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n821), .B1(new_n213), .B2(new_n413), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n242), .A2(new_n712), .A3(new_n492), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n767), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n492), .B1(new_n805), .B2(new_n864), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n205), .B2(new_n800), .C1(new_n206), .C2(new_n789), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n777), .A2(G303), .B1(new_n779), .B2(G311), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n782), .A2(G294), .B1(G317), .B2(new_n814), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n797), .B2(new_n640), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1014), .A2(new_n640), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1011), .B(new_n1016), .C1(new_n810), .C2(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n800), .A2(new_n224), .B1(new_n797), .B2(new_n259), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n789), .A2(new_n222), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n1019), .A2(new_n1020), .A3(new_n288), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n782), .A2(G159), .B1(G50), .B2(new_n805), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT108), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(KEYINPUT108), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n777), .A2(G150), .B1(G137), .B2(new_n814), .ZN(new_n1026));
  INV_X1    g0826(.A(G143), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n780), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1018), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1030), .A2(KEYINPUT47), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n774), .B1(new_n1030), .B2(KEYINPUT47), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1009), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n831), .B2(new_n965), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1006), .A2(new_n1034), .ZN(G387));
  NAND3_X1  g0835(.A1(new_n700), .A2(new_n703), .A3(new_n820), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n822), .B1(new_n239), .B2(new_n301), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n715), .B2(new_n825), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n410), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1039));
  OAI21_X1  g0839(.A(KEYINPUT50), .B1(new_n410), .B2(G50), .ZN(new_n1040));
  AOI21_X1  g0840(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1039), .A2(new_n715), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1038), .A2(new_n1042), .B1(new_n206), .B2(new_n712), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n821), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n767), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n492), .B1(new_n780), .B2(new_n793), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n797), .A2(new_n224), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n789), .A2(new_n413), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n263), .A2(new_n782), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n801), .A2(G97), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n785), .A2(new_n222), .B1(new_n792), .B2(new_n851), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G50), .B2(new_n777), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n789), .A2(new_n863), .B1(new_n797), .B2(new_n497), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n777), .A2(G317), .B1(new_n779), .B2(G322), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n782), .A2(G311), .B1(G303), .B2(new_n805), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT48), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n1059), .B2(new_n1058), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT49), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n492), .B1(new_n814), .B2(G326), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n640), .B2(new_n800), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1054), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1045), .B1(new_n1065), .B2(new_n773), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1002), .A2(new_n766), .B1(new_n1036), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n762), .A2(new_n999), .A3(new_n1000), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n762), .B1(new_n999), .B2(new_n1000), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT109), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n713), .B(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1002), .A2(KEYINPUT109), .A3(new_n762), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(G393));
  INV_X1    g0873(.A(new_n1003), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1068), .B1(new_n1074), .B2(new_n994), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1004), .A2(new_n1075), .A3(new_n713), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n247), .A2(new_n822), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n821), .B1(new_n205), .B2(new_n213), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n767), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n956), .A2(new_n831), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n777), .A2(G311), .B1(new_n779), .B2(G317), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1082));
  XNOR2_X1  g0882(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n807), .A2(G116), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n782), .A2(G303), .B1(G294), .B2(new_n805), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1083), .A2(new_n288), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(G322), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n797), .A2(new_n863), .B1(new_n792), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT111), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n802), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n777), .A2(G159), .B1(new_n779), .B2(G150), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n792), .A2(new_n1027), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n492), .B1(new_n785), .B2(new_n410), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(G50), .C2(new_n782), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n807), .A2(G77), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n798), .A2(G68), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1096), .A2(new_n867), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1086), .A2(new_n1091), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1079), .B(new_n1080), .C1(new_n773), .C2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1074), .A2(new_n994), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1102), .B2(new_n766), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1076), .A2(new_n1103), .ZN(G390));
  AOI21_X1  g0904(.A(new_n731), .B1(new_n935), .B2(new_n758), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n923), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n914), .B1(new_n841), .B2(new_n916), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1108), .A2(new_n904), .B1(new_n903), .B2(new_n908), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n922), .A2(new_n904), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n728), .A2(new_n837), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n835), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n914), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1107), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n916), .B1(new_n720), .B2(new_n839), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n914), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n904), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n903), .A2(new_n908), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1112), .A2(new_n914), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1110), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT112), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n761), .A2(new_n839), .A3(new_n914), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1114), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1117), .A2(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1123), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n766), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1118), .A2(new_n818), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n767), .B1(new_n847), .B2(new_n263), .ZN(new_n1132));
  INV_X1    g0932(.A(G283), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n778), .A2(new_n640), .B1(new_n780), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G97), .B2(new_n805), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n782), .A2(G107), .B1(G294), .B2(new_n814), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1135), .A2(new_n288), .A3(new_n1097), .A4(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n857), .B1(new_n858), .B2(new_n360), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n798), .A2(G150), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n814), .A2(G125), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1141), .B1(new_n785), .B2(new_n1142), .C1(new_n783), .C2(new_n849), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n779), .A2(G128), .ZN(new_n1144));
  INV_X1    g0944(.A(G132), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n289), .C1(new_n778), .C2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n789), .A2(new_n793), .B1(new_n800), .B2(new_n202), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1137), .A2(new_n1138), .B1(new_n1140), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1132), .B1(new_n1149), .B2(new_n773), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1131), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1112), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1124), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n914), .B1(new_n1105), .B2(new_n839), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n914), .B1(new_n761), .B2(new_n839), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT114), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n731), .B(new_n838), .C1(new_n758), .C2(new_n760), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT114), .B1(new_n1160), .B2(new_n914), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1161), .A3(new_n1106), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1115), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT113), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n940), .A2(new_n731), .A3(new_n674), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n876), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1105), .A2(new_n479), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1168), .A2(KEYINPUT113), .A3(new_n673), .A4(new_n875), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n713), .B1(new_n1171), .B2(new_n1129), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1106), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1160), .A2(KEYINPUT114), .A3(new_n914), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1163), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1156), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1170), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1119), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(KEYINPUT112), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1181), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1152), .B1(new_n1172), .B2(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1170), .B1(new_n1129), .B2(new_n1177), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n909), .A2(new_n917), .A3(new_n918), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n473), .A2(new_n477), .A3(new_n912), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n912), .B1(new_n473), .B2(new_n477), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n839), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n935), .B2(new_n758), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(new_n937), .B1(new_n933), .B2(KEYINPUT40), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1187), .B1(new_n1192), .B2(new_n731), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n939), .A2(G330), .A3(new_n919), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n277), .A2(new_n694), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT55), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n321), .B(new_n1196), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1198));
  XNOR2_X1  g0998(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1193), .A2(new_n1194), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1185), .B1(new_n1186), .B2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n939), .A2(G330), .A3(new_n919), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n919), .B1(new_n939), .B2(G330), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1199), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1193), .A2(new_n1194), .A3(new_n1200), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1185), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1178), .B1(new_n1182), .B2(new_n1164), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n714), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1204), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT119), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n765), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n767), .B1(new_n847), .B2(G50), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n353), .A2(new_n300), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n264), .A2(new_n300), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n202), .A3(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n778), .A2(new_n206), .B1(new_n413), .B2(new_n785), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n800), .A2(new_n259), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1219), .A2(new_n1020), .A3(new_n1047), .A4(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n779), .A2(G116), .B1(G283), .B2(new_n814), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1216), .B1(new_n782), .B2(G97), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1218), .B1(new_n1224), .B2(KEYINPUT58), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT115), .Z(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n777), .A2(G128), .B1(new_n779), .B2(G125), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1228), .B1(new_n851), .B2(new_n789), .C1(new_n797), .C2(new_n1142), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n782), .A2(G132), .B1(G137), .B2(new_n805), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT116), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1217), .B1(new_n814), .B2(G124), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT59), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1235), .B1(new_n793), .B2(new_n800), .C1(new_n1232), .C2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1226), .B(new_n1227), .C1(new_n1234), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1215), .B1(new_n1238), .B2(new_n773), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1199), .B2(new_n819), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT118), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1213), .B1(new_n1214), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n766), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(KEYINPUT119), .A3(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1212), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(G375));
  NAND3_X1  g1048(.A1(new_n1175), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(new_n1171), .A3(new_n986), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT120), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n767), .B1(new_n847), .B2(G68), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n914), .A2(new_n819), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n779), .A2(G132), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n778), .B2(new_n849), .C1(new_n783), .C2(new_n1142), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT121), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n492), .B1(new_n785), .B2(new_n851), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(G128), .B2(new_n814), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1220), .B1(G50), .B2(new_n807), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(new_n858), .C2(new_n793), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n778), .A2(new_n1133), .B1(new_n785), .B2(new_n206), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G303), .B2(new_n814), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1048), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n782), .A2(G116), .B1(new_n779), .B2(G294), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n288), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n801), .A2(G77), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n858), .B2(new_n205), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1257), .A2(new_n1261), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n1253), .B(new_n1254), .C1(new_n773), .C2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1177), .B2(new_n766), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1252), .A2(new_n1271), .ZN(G381));
  OAI211_X1 g1072(.A(new_n833), .B(new_n1067), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1273));
  OR3_X1    g1073(.A1(G390), .A2(G384), .A3(new_n1273), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(G381), .A2(G387), .A3(G378), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1247), .ZN(G407));
  NAND2_X1  g1076(.A1(new_n1130), .A2(new_n1151), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n714), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1171), .A2(new_n1129), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1247), .A2(new_n695), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(G393), .A2(G396), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G390), .A2(new_n1273), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1273), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1076), .A3(new_n1103), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G387), .A2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1006), .A2(new_n1284), .A3(new_n1286), .A4(new_n1034), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(G213), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1291), .A2(G343), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1212), .A2(new_n1246), .A3(G378), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1186), .A2(new_n1203), .A3(new_n986), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1244), .A2(new_n1241), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1280), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1292), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT122), .B1(new_n1249), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n714), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT122), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1164), .A2(new_n1301), .A3(KEYINPUT60), .A4(new_n1170), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1249), .A2(new_n1298), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1299), .A2(new_n1300), .A3(new_n1302), .A4(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1271), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OR2_X1    g1107(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1307), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1304), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1297), .A2(KEYINPUT62), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT62), .B1(new_n1297), .B2(new_n1312), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(new_n1313), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1297), .A2(new_n1312), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1315), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1292), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1292), .A2(G2897), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1304), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1308), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1310), .A2(new_n1311), .A3(new_n1323), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1322), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1319), .A2(new_n1330), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1290), .B1(new_n1316), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1288), .A2(new_n1333), .A3(new_n1289), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1317), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(KEYINPUT63), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1322), .A2(new_n1329), .A3(KEYINPUT124), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1317), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1322), .A2(new_n1329), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .A4(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1332), .A2(new_n1343), .ZN(G405));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1247), .B(new_n1280), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1312), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1345), .B(new_n1290), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1350), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1290), .A2(new_n1345), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1288), .A2(KEYINPUT126), .A3(new_n1289), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .A4(new_n1348), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1351), .A2(new_n1355), .ZN(G402));
endmodule


