

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  INV_X1 U323 ( .A(KEYINPUT94), .ZN(n366) );
  XNOR2_X1 U324 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U325 ( .A(n451), .B(KEYINPUT113), .ZN(n452) );
  NOR2_X1 U326 ( .A1(n475), .A2(n532), .ZN(n566) );
  XNOR2_X1 U327 ( .A(n378), .B(n377), .ZN(n380) );
  XNOR2_X1 U328 ( .A(n392), .B(n376), .ZN(n377) );
  XOR2_X1 U329 ( .A(KEYINPUT70), .B(G78GAT), .Z(n291) );
  INV_X1 U330 ( .A(KEYINPUT45), .ZN(n451) );
  XNOR2_X1 U331 ( .A(n457), .B(KEYINPUT112), .ZN(n458) );
  XNOR2_X1 U332 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U333 ( .A1(n461), .A2(n565), .ZN(n462) );
  XNOR2_X1 U334 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U335 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U336 ( .A(n417), .B(n368), .ZN(n372) );
  XNOR2_X1 U337 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U338 ( .A(n302), .B(n301), .ZN(n303) );
  OR2_X1 U339 ( .A1(n585), .A2(n414), .ZN(n415) );
  XNOR2_X1 U340 ( .A(n429), .B(n428), .ZN(n430) );
  NOR2_X1 U341 ( .A1(n549), .A2(n508), .ZN(n533) );
  NOR2_X1 U342 ( .A1(n412), .A2(n411), .ZN(n483) );
  AND2_X1 U343 ( .A1(n512), .A2(n467), .ZN(n572) );
  OR2_X1 U344 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U345 ( .A(n440), .B(n307), .ZN(n561) );
  XOR2_X1 U346 ( .A(KEYINPUT110), .B(n447), .Z(n530) );
  XNOR2_X1 U347 ( .A(n471), .B(G176GAT), .ZN(n472) );
  XNOR2_X1 U348 ( .A(n448), .B(G106GAT), .ZN(n449) );
  XNOR2_X1 U349 ( .A(n473), .B(n472), .ZN(G1349GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT7), .B(G50GAT), .Z(n293) );
  XNOR2_X1 U351 ( .A(KEYINPUT8), .B(G36GAT), .ZN(n292) );
  XNOR2_X1 U352 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U353 ( .A(G29GAT), .B(n294), .Z(n440) );
  XOR2_X1 U354 ( .A(G106GAT), .B(G218GAT), .Z(n296) );
  XOR2_X1 U355 ( .A(G162GAT), .B(KEYINPUT76), .Z(n397) );
  XOR2_X1 U356 ( .A(G134GAT), .B(G190GAT), .Z(n327) );
  XNOR2_X1 U357 ( .A(n397), .B(n327), .ZN(n295) );
  XNOR2_X1 U358 ( .A(n296), .B(n295), .ZN(n302) );
  XOR2_X1 U359 ( .A(KEYINPUT11), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U360 ( .A(G99GAT), .B(G92GAT), .ZN(n297) );
  XNOR2_X1 U361 ( .A(n298), .B(n297), .ZN(n300) );
  AND2_X1 U362 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U363 ( .A(n303), .B(KEYINPUT10), .Z(n306) );
  XNOR2_X1 U364 ( .A(G85GAT), .B(KEYINPUT71), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n304), .B(KEYINPUT72), .ZN(n431) );
  XNOR2_X1 U366 ( .A(n431), .B(KEYINPUT9), .ZN(n305) );
  XNOR2_X1 U367 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U368 ( .A(KEYINPUT36), .B(n561), .ZN(n585) );
  XOR2_X1 U369 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n309) );
  XNOR2_X1 U370 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n308) );
  XNOR2_X1 U371 ( .A(n309), .B(n308), .ZN(n317) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G78GAT), .Z(n311) );
  XNOR2_X1 U374 ( .A(G155GAT), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U375 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G211GAT), .Z(n312) );
  XNOR2_X1 U377 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n325) );
  XNOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT67), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n318), .B(KEYINPUT13), .ZN(n419) );
  XOR2_X1 U382 ( .A(G64GAT), .B(KEYINPUT77), .Z(n320) );
  XNOR2_X1 U383 ( .A(G71GAT), .B(G183GAT), .ZN(n319) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n419), .B(n321), .ZN(n323) );
  XOR2_X1 U386 ( .A(G1GAT), .B(G8GAT), .Z(n322) );
  XOR2_X1 U387 ( .A(KEYINPUT64), .B(n322), .Z(n439) );
  XOR2_X1 U388 ( .A(n323), .B(n439), .Z(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n565) );
  XNOR2_X1 U390 ( .A(G120GAT), .B(G99GAT), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n326), .B(G71GAT), .ZN(n416) );
  XOR2_X1 U392 ( .A(n327), .B(n416), .Z(n329) );
  NAND2_X1 U393 ( .A1(G227GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U395 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n331) );
  XNOR2_X1 U396 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n338) );
  XNOR2_X1 U399 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n334), .B(KEYINPUT0), .ZN(n355) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G15GAT), .Z(n336) );
  XNOR2_X1 U402 ( .A(G113GAT), .B(G43GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n437) );
  XNOR2_X1 U404 ( .A(n355), .B(n437), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U406 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n340) );
  XNOR2_X1 U407 ( .A(KEYINPUT18), .B(G176GAT), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U409 ( .A(G183GAT), .B(n341), .ZN(n379) );
  XNOR2_X1 U410 ( .A(n342), .B(n379), .ZN(n532) );
  XNOR2_X1 U411 ( .A(n532), .B(KEYINPUT84), .ZN(n400) );
  XOR2_X1 U412 ( .A(G155GAT), .B(KEYINPUT3), .Z(n344) );
  XNOR2_X1 U413 ( .A(KEYINPUT2), .B(KEYINPUT88), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n388) );
  XOR2_X1 U415 ( .A(n388), .B(KEYINPUT5), .Z(n346) );
  NAND2_X1 U416 ( .A1(G225GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U418 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n348) );
  XNOR2_X1 U419 ( .A(G57GAT), .B(G1GAT), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U421 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U422 ( .A(G120GAT), .B(G113GAT), .Z(n352) );
  XNOR2_X1 U423 ( .A(G141GAT), .B(G148GAT), .ZN(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n359) );
  XOR2_X1 U426 ( .A(G162GAT), .B(G85GAT), .Z(n357) );
  XNOR2_X1 U427 ( .A(G29GAT), .B(n355), .ZN(n356) );
  XNOR2_X1 U428 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U429 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U430 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n361) );
  XNOR2_X1 U431 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n362), .B(G134GAT), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n512) );
  XNOR2_X1 U435 ( .A(G92GAT), .B(G64GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n365), .B(G204GAT), .ZN(n417) );
  XNOR2_X1 U437 ( .A(G36GAT), .B(G190GAT), .ZN(n367) );
  XOR2_X1 U438 ( .A(KEYINPUT77), .B(KEYINPUT95), .Z(n370) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U441 ( .A(n372), .B(n371), .Z(n378) );
  XOR2_X1 U442 ( .A(KEYINPUT87), .B(G197GAT), .Z(n374) );
  XNOR2_X1 U443 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n373) );
  XNOR2_X1 U444 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U445 ( .A(G211GAT), .B(n375), .Z(n392) );
  XNOR2_X1 U446 ( .A(G8GAT), .B(G169GAT), .ZN(n376) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n516) );
  XNOR2_X1 U448 ( .A(KEYINPUT27), .B(n516), .ZN(n407) );
  NOR2_X1 U449 ( .A1(n512), .A2(n407), .ZN(n381) );
  XOR2_X1 U450 ( .A(KEYINPUT96), .B(n381), .Z(n549) );
  XOR2_X1 U451 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n383) );
  XNOR2_X1 U452 ( .A(G50GAT), .B(KEYINPUT22), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U454 ( .A(KEYINPUT85), .B(KEYINPUT89), .Z(n385) );
  XNOR2_X1 U455 ( .A(KEYINPUT86), .B(KEYINPUT90), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U457 ( .A(n387), .B(n386), .Z(n394) );
  XOR2_X1 U458 ( .A(n388), .B(G204GAT), .Z(n390) );
  NAND2_X1 U459 ( .A1(G228GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U460 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U462 ( .A(n394), .B(n393), .ZN(n396) );
  XNOR2_X1 U463 ( .A(G148GAT), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n291), .B(n395), .ZN(n418) );
  XOR2_X1 U465 ( .A(n396), .B(n418), .Z(n399) );
  XOR2_X1 U466 ( .A(G141GAT), .B(G22GAT), .Z(n444) );
  XNOR2_X1 U467 ( .A(n397), .B(n444), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n405) );
  XOR2_X1 U469 ( .A(n405), .B(KEYINPUT28), .Z(n521) );
  INV_X1 U470 ( .A(n521), .ZN(n508) );
  NAND2_X1 U471 ( .A1(n400), .A2(n533), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n401), .B(KEYINPUT97), .ZN(n412) );
  INV_X1 U473 ( .A(n512), .ZN(n525) );
  INV_X1 U474 ( .A(n532), .ZN(n529) );
  INV_X1 U475 ( .A(n516), .ZN(n527) );
  NAND2_X1 U476 ( .A1(n529), .A2(n527), .ZN(n402) );
  INV_X1 U477 ( .A(n405), .ZN(n468) );
  NAND2_X1 U478 ( .A1(n402), .A2(n468), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n403), .B(KEYINPUT25), .ZN(n404) );
  XNOR2_X1 U480 ( .A(n404), .B(KEYINPUT98), .ZN(n409) );
  NAND2_X1 U481 ( .A1(n532), .A2(n405), .ZN(n406) );
  XNOR2_X1 U482 ( .A(n406), .B(KEYINPUT26), .ZN(n550) );
  NOR2_X1 U483 ( .A1(n550), .A2(n407), .ZN(n408) );
  NOR2_X1 U484 ( .A1(n409), .A2(n408), .ZN(n410) );
  NOR2_X1 U485 ( .A1(n525), .A2(n410), .ZN(n411) );
  NOR2_X1 U486 ( .A1(n565), .A2(n483), .ZN(n413) );
  XNOR2_X1 U487 ( .A(n413), .B(KEYINPUT103), .ZN(n414) );
  XNOR2_X1 U488 ( .A(KEYINPUT37), .B(n415), .ZN(n498) );
  XOR2_X1 U489 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U490 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT74), .B(KEYINPUT68), .Z(n423) );
  XNOR2_X1 U493 ( .A(KEYINPUT69), .B(KEYINPUT73), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U495 ( .A(G176GAT), .B(KEYINPUT31), .Z(n424) );
  XNOR2_X1 U496 ( .A(n425), .B(n424), .ZN(n427) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XOR2_X1 U498 ( .A(n430), .B(KEYINPUT33), .Z(n433) );
  XNOR2_X1 U499 ( .A(n431), .B(KEYINPUT32), .ZN(n432) );
  XNOR2_X1 U500 ( .A(n433), .B(n432), .ZN(n578) );
  INV_X1 U501 ( .A(KEYINPUT41), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n578), .B(n434), .ZN(n554) );
  INV_X1 U503 ( .A(n554), .ZN(n538) );
  XOR2_X1 U504 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n436) );
  XNOR2_X1 U505 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n435) );
  XNOR2_X1 U506 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U507 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U508 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U509 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U510 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U511 ( .A1(G229GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n573) );
  AND2_X1 U513 ( .A1(n538), .A2(n573), .ZN(n511) );
  NAND2_X1 U514 ( .A1(n498), .A2(n511), .ZN(n447) );
  NAND2_X1 U515 ( .A1(n530), .A2(n508), .ZN(n450) );
  XOR2_X1 U516 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n448) );
  XNOR2_X1 U517 ( .A(n450), .B(n449), .ZN(G1339GAT) );
  XOR2_X1 U518 ( .A(n573), .B(KEYINPUT66), .Z(n563) );
  INV_X1 U519 ( .A(n565), .ZN(n581) );
  NOR2_X1 U520 ( .A1(n585), .A2(n581), .ZN(n453) );
  NAND2_X1 U521 ( .A1(n454), .A2(n578), .ZN(n455) );
  NOR2_X1 U522 ( .A1(n563), .A2(n455), .ZN(n456) );
  XNOR2_X1 U523 ( .A(KEYINPUT114), .B(n456), .ZN(n464) );
  NOR2_X1 U524 ( .A1(n573), .A2(n554), .ZN(n459) );
  INV_X1 U525 ( .A(KEYINPUT46), .ZN(n457) );
  NAND2_X1 U526 ( .A1(n460), .A2(n561), .ZN(n461) );
  XOR2_X1 U527 ( .A(KEYINPUT47), .B(n462), .Z(n463) );
  NOR2_X1 U528 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U529 ( .A(KEYINPUT48), .B(n465), .ZN(n548) );
  NOR2_X1 U530 ( .A1(n516), .A2(n548), .ZN(n466) );
  XNOR2_X1 U531 ( .A(KEYINPUT54), .B(n466), .ZN(n467) );
  NAND2_X1 U532 ( .A1(n572), .A2(n468), .ZN(n470) );
  XOR2_X1 U533 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n566), .A2(n538), .ZN(n473) );
  XOR2_X1 U536 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n471) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n477) );
  INV_X1 U539 ( .A(n561), .ZN(n543) );
  NAND2_X1 U540 ( .A1(n529), .A2(n543), .ZN(n474) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT79), .Z(n481) );
  NAND2_X1 U545 ( .A1(n565), .A2(n561), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  NOR2_X1 U547 ( .A1(n483), .A2(n482), .ZN(n510) );
  NAND2_X1 U548 ( .A1(n563), .A2(n578), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n484), .B(KEYINPUT75), .ZN(n499) );
  NAND2_X1 U550 ( .A1(n510), .A2(n499), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n485), .B(KEYINPUT99), .ZN(n494) );
  NAND2_X1 U552 ( .A1(n494), .A2(n525), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  XOR2_X1 U555 ( .A(G8GAT), .B(KEYINPUT101), .Z(n490) );
  NAND2_X1 U556 ( .A1(n494), .A2(n527), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n492) );
  NAND2_X1 U559 ( .A1(n494), .A2(n529), .ZN(n491) );
  XNOR2_X1 U560 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U562 ( .A1(n508), .A2(n494), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U566 ( .A(n497), .B(n496), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n501) );
  NAND2_X1 U568 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(n507) );
  NAND2_X1 U570 ( .A1(n525), .A2(n507), .ZN(n502) );
  XOR2_X1 U571 ( .A(n503), .B(n502), .Z(G1328GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n527), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U574 ( .A1(n529), .A2(n507), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U577 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n512), .A2(n520), .ZN(n514) );
  XNOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U583 ( .A(G57GAT), .B(n515), .ZN(G1332GAT) );
  NOR2_X1 U584 ( .A1(n516), .A2(n520), .ZN(n517) );
  XOR2_X1 U585 ( .A(KEYINPUT108), .B(n517), .Z(n518) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U587 ( .A1(n532), .A2(n520), .ZN(n519) );
  XOR2_X1 U588 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U589 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U590 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NAND2_X1 U593 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n526), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U599 ( .A1(n532), .A2(n548), .ZN(n534) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(KEYINPUT115), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n544), .A2(n563), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT116), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n544), .A2(n538), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U608 ( .A1(n544), .A2(n565), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U616 ( .A(n550), .ZN(n571) );
  NAND2_X1 U617 ( .A1(n551), .A2(n571), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n573), .A2(n560), .ZN(n552) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(n552), .Z(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U621 ( .A1(n560), .A2(n554), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n581), .A2(n560), .ZN(n559) );
  XOR2_X1 U627 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G183GAT), .B(KEYINPUT121), .Z(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n573), .A2(n584), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(n577), .B(n576), .Z(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n584), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(n582), .Z(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

