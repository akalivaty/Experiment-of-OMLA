//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1230, new_n1231,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1310, new_n1311;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G77), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n241), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n214), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(new_n251), .B2(new_n253), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n255), .B(new_n257), .C1(G1), .C2(new_n206), .ZN(new_n258));
  OR2_X1    g0058(.A1(new_n258), .A2(new_n242), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n251), .A2(new_n242), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n206), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n206), .B1(new_n201), .B2(new_n242), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n253), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(new_n260), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G223), .ZN(new_n278));
  OAI221_X1 g0078(.A(new_n276), .B1(new_n218), .B2(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(G274), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n288), .B1(G226), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n269), .B(new_n295), .C1(G179), .C2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n259), .A2(new_n260), .A3(new_n268), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n293), .A2(G200), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n269), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n281), .A2(new_n292), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n300), .A2(new_n306), .B1(new_n307), .B2(G190), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(KEYINPUT9), .A2(new_n298), .B1(new_n301), .B2(KEYINPUT70), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n311), .A2(new_n312), .A3(new_n308), .A4(new_n304), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n297), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n251), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n258), .B2(new_n315), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n272), .A2(new_n206), .A3(new_n273), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT7), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n273), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n244), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G58), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n244), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n325), .B2(new_n201), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n264), .A2(G159), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n318), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n253), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n322), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n319), .A2(new_n332), .A3(new_n320), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(G68), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n328), .A2(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n317), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n278), .A2(new_n275), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n338), .B1(G226), .B2(new_n275), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n286), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G232), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n287), .B1(new_n344), .B2(new_n290), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n346), .A2(new_n294), .ZN(new_n347));
  INV_X1    g0147(.A(G179), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n343), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT18), .B1(new_n337), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n334), .A2(new_n335), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(new_n253), .A3(new_n329), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n258), .A2(new_n315), .ZN(new_n355));
  INV_X1    g0155(.A(new_n316), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G190), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n346), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n343), .B2(new_n345), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n354), .A2(new_n366), .A3(new_n357), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n337), .A2(KEYINPUT17), .A3(new_n366), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n361), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n244), .A2(G20), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n373), .B1(new_n262), .B2(new_n218), .C1(new_n265), .C2(new_n242), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n253), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT11), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n378), .A2(new_n205), .A3(G13), .A4(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n253), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(G68), .C1(G1), .C2(new_n206), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G13), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(G1), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n385), .A2(KEYINPUT12), .A3(new_n373), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n377), .A2(new_n379), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n244), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(KEYINPUT12), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n274), .A2(G226), .A3(new_n275), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G33), .A2(G97), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n280), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n288), .B1(G238), .B2(new_n291), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g0201(.A(G200), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n404), .A2(G190), .A3(new_n399), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n391), .ZN(new_n408));
  OAI21_X1  g0208(.A(G169), .B1(new_n400), .B2(new_n401), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT14), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(G169), .C1(new_n400), .C2(new_n401), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n404), .A2(G179), .A3(new_n399), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n416));
  INV_X1    g0216(.A(G107), .ZN(new_n417));
  INV_X1    g0217(.A(G238), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n416), .B1(new_n417), .B2(new_n274), .C1(new_n277), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n280), .ZN(new_n420));
  INV_X1    g0220(.A(new_n217), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n288), .B1(new_n421), .B2(new_n291), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n348), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n387), .A2(G77), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n315), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT15), .B(G87), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n429), .B1(new_n206), .B2(new_n218), .C1(new_n262), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n426), .B1(new_n431), .B2(new_n253), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n380), .B(G77), .C1(G1), .C2(new_n206), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n423), .A2(new_n294), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n425), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n432), .B(new_n433), .C1(new_n423), .C2(new_n362), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n424), .A2(new_n364), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n314), .A2(new_n372), .A3(new_n415), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G116), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n205), .B2(G33), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n380), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT74), .A2(G116), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT74), .A2(G116), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n388), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(G20), .B1(G33), .B2(G283), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n271), .A2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g0252(.A(KEYINPUT74), .B(G116), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n253), .C1(new_n453), .C2(new_n206), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT20), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n448), .A2(G20), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n450), .A2(new_n451), .B1(new_n252), .B2(new_n214), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT20), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n445), .B(new_n449), .C1(new_n456), .C2(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n275), .A2(G264), .ZN(new_n461));
  NOR2_X1   g0261(.A1(G257), .A2(G1698), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n461), .A2(new_n462), .B1(new_n339), .B2(new_n340), .ZN(new_n463));
  INV_X1    g0263(.A(G303), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n272), .A2(new_n464), .A3(new_n273), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n280), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n283), .A2(G1), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(G274), .A3(new_n286), .A4(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G270), .A3(new_n286), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n466), .A2(new_n469), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n460), .A2(KEYINPUT21), .A3(G169), .A4(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n348), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n460), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(G169), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT21), .B1(new_n480), .B2(new_n460), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT76), .ZN(new_n483));
  INV_X1    g0283(.A(new_n460), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT75), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n474), .A2(G200), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n466), .A2(new_n469), .A3(new_n473), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G190), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n454), .A2(new_n455), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n457), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n388), .A2(new_n448), .B1(new_n380), .B2(new_n444), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n492), .B(new_n493), .C1(new_n362), .C2(new_n474), .ZN(new_n494));
  INV_X1    g0294(.A(new_n486), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT75), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n482), .A2(new_n483), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n483), .B1(new_n482), .B2(new_n497), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n472), .A2(G257), .A3(new_n286), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n469), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI211_X1 g0303(.A(G244), .B(new_n275), .C1(new_n339), .C2(new_n340), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G283), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n271), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G250), .A2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(KEYINPUT4), .A2(G244), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(G1698), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n274), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n286), .B1(new_n506), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT72), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI211_X1 g0315(.A(KEYINPUT72), .B(new_n286), .C1(new_n506), .C2(new_n512), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n348), .B(new_n503), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n506), .A2(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n280), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n503), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n294), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT6), .ZN(new_n522));
  INV_X1    g0322(.A(G97), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n522), .A2(new_n523), .A3(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(G97), .B(G107), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(new_n206), .B1(new_n218), .B2(new_n265), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n417), .B1(new_n321), .B2(new_n322), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n253), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n250), .A2(G97), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n253), .B(new_n251), .C1(new_n205), .C2(G33), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(G97), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n517), .A2(new_n521), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n418), .A2(new_n275), .ZN(new_n535));
  INV_X1    g0335(.A(G244), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G1698), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n537), .C1(new_n339), .C2(new_n340), .ZN(new_n538));
  OAI21_X1  g0338(.A(G33), .B1(new_n446), .B2(new_n447), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n280), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT73), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n283), .B2(G1), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n205), .A2(KEYINPUT73), .A3(G45), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n286), .A2(new_n543), .A3(G250), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n286), .A2(G274), .A3(new_n468), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n541), .A2(new_n547), .A3(G190), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT19), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n206), .B1(new_n394), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G87), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n551), .A2(new_n523), .A3(new_n417), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n206), .B(G68), .C1(new_n339), .C2(new_n340), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n549), .B1(new_n262), .B2(new_n523), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n253), .B1(new_n388), .B2(new_n430), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n531), .A2(G87), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n286), .B1(new_n538), .B2(new_n539), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n545), .A2(new_n546), .ZN(new_n560));
  OAI21_X1  g0360(.A(G200), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n548), .A2(new_n557), .A3(new_n558), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n556), .A2(new_n253), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n388), .A2(new_n430), .ZN(new_n564));
  INV_X1    g0364(.A(new_n430), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n254), .B(new_n565), .C1(G1), .C2(new_n271), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n294), .B1(new_n559), .B2(new_n560), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n541), .A2(new_n547), .A3(new_n348), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n513), .B(new_n514), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n364), .B1(new_n572), .B2(new_n503), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n519), .A2(new_n503), .A3(G190), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n529), .A3(new_n532), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n534), .B(new_n571), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n472), .A2(G264), .A3(new_n286), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G250), .A2(G1698), .ZN(new_n578));
  INV_X1    g0378(.A(G257), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n579), .B2(G1698), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n580), .A2(new_n274), .B1(G33), .B2(G294), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n469), .B(new_n577), .C1(new_n581), .C2(new_n286), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n364), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT78), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n581), .B2(new_n286), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n577), .A2(new_n469), .ZN(new_n586));
  OR2_X1    g0386(.A1(G250), .A2(G1698), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n579), .A2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n587), .B(new_n588), .C1(new_n339), .C2(new_n340), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G33), .A2(G294), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(KEYINPUT78), .A3(new_n280), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n583), .B1(new_n593), .B2(G190), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n206), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n595));
  NAND2_X1  g0395(.A1(KEYINPUT77), .A2(KEYINPUT22), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n274), .A2(new_n206), .A3(G87), .A4(new_n596), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  INV_X1    g0401(.A(new_n447), .ZN(new_n602));
  NAND2_X1  g0402(.A1(KEYINPUT74), .A2(G116), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n271), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n206), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n417), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n604), .A2(new_n206), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n600), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n601), .B1(new_n600), .B2(new_n608), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n253), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n254), .B1(G1), .B2(new_n271), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n417), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n251), .A2(new_n417), .ZN(new_n614));
  XNOR2_X1  g0414(.A(new_n614), .B(KEYINPUT25), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n594), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n600), .A2(new_n608), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT24), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n600), .A2(new_n608), .A3(new_n601), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n330), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n616), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n582), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n593), .A2(G169), .B1(new_n624), .B2(G179), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n617), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n576), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n442), .A2(new_n500), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(new_n570), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n594), .A2(new_n611), .A3(new_n616), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n593), .A2(G169), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(G179), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n621), .B2(new_n622), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n630), .B1(new_n482), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n576), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n629), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n529), .A2(new_n532), .B1(new_n520), .B2(new_n294), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n571), .A2(KEYINPUT26), .A3(new_n517), .A4(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT79), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n534), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n643), .A2(KEYINPUT79), .A3(KEYINPUT26), .A4(new_n571), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n562), .A2(new_n570), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n534), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n644), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n442), .B1(new_n638), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n414), .A2(new_n408), .B1(new_n437), .B2(new_n406), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n351), .B(new_n360), .C1(new_n651), .C2(new_n371), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n310), .A2(new_n313), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n297), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n650), .A2(new_n654), .ZN(G369));
  OR3_X1    g0455(.A1(new_n385), .A2(KEYINPUT27), .A3(G20), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT27), .B1(new_n385), .B2(G20), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(G213), .A3(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G343), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n460), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n500), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n662), .B1(new_n482), .B2(new_n661), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n625), .B1(new_n611), .B2(new_n616), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(new_n630), .ZN(new_n666));
  INV_X1    g0466(.A(new_n660), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n623), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n634), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n482), .A2(new_n660), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n666), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n670), .B(new_n672), .C1(new_n634), .C2(new_n660), .ZN(G399));
  INV_X1    g0473(.A(new_n209), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n552), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n212), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n647), .A2(new_n640), .ZN(new_n681));
  INV_X1    g0481(.A(new_n481), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n477), .A3(new_n475), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n617), .B1(new_n683), .B2(new_n665), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n681), .B(new_n570), .C1(new_n684), .C2(new_n576), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT82), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(new_n667), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n685), .B2(new_n667), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT29), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n660), .B1(new_n637), .B2(new_n648), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT29), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT81), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT80), .ZN(new_n695));
  INV_X1    g0495(.A(new_n214), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n467), .A2(new_n468), .B1(new_n696), .B2(new_n285), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n280), .A2(new_n591), .B1(new_n697), .B2(G264), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n559), .A2(new_n560), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n487), .A2(new_n698), .A3(new_n699), .A4(G179), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n519), .A2(new_n503), .A3(KEYINPUT30), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n695), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT30), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n513), .A2(new_n502), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n703), .A2(new_n705), .A3(KEYINPUT80), .A4(new_n476), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n541), .A2(new_n547), .ZN(new_n708));
  AND4_X1   g0508(.A1(new_n348), .A2(new_n708), .A3(new_n582), .A4(new_n474), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n503), .B1(new_n515), .B2(new_n516), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n704), .B1(new_n700), .B2(new_n520), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n694), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n702), .A2(new_n706), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT81), .A3(new_n712), .A4(new_n711), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n714), .A2(new_n660), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n627), .B(new_n667), .C1(new_n498), .C2(new_n499), .ZN(new_n720));
  OAI211_X1 g0520(.A(KEYINPUT31), .B(new_n660), .C1(new_n707), .C2(new_n713), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n693), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n680), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(new_n383), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n205), .B1(new_n727), .B2(G45), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n676), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n663), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n214), .B1(G20), .B2(new_n294), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT84), .Z(new_n737));
  INV_X1    g0537(.A(new_n274), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n209), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT83), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n213), .A2(new_n283), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n740), .B(new_n741), .C1(new_n283), .C2(new_n248), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n674), .A2(new_n738), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n743), .A2(G355), .B1(new_n443), .B2(new_n674), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n737), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n362), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n206), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G97), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n206), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n362), .A3(G200), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(new_n362), .A3(new_n364), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT87), .B(G159), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n749), .B1(new_n417), .B2(new_n751), .C1(KEYINPUT32), .C2(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n738), .B(new_n757), .C1(KEYINPUT32), .C2(new_n756), .ZN(new_n758));
  NAND2_X1  g0558(.A1(G20), .A2(G179), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT85), .Z(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n364), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n362), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n364), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n242), .A2(new_n763), .B1(new_n766), .B2(new_n244), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n764), .A2(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT88), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n769), .A2(new_n218), .B1(new_n551), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n761), .A2(G200), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT86), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n758), .B(new_n776), .C1(new_n324), .C2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI22_X1  g0580(.A1(G322), .A2(new_n777), .B1(new_n765), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT89), .B(G326), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n769), .C1(new_n763), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G329), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n751), .A2(new_n507), .B1(new_n752), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT90), .Z(new_n787));
  AOI21_X1  g0587(.A(new_n274), .B1(new_n748), .B2(G294), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n788), .C1(new_n464), .C2(new_n774), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n779), .B1(new_n784), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n745), .B1(new_n790), .B2(new_n735), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n729), .B1(new_n734), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n664), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n663), .A2(G330), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n792), .B1(new_n729), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT91), .Z(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  INV_X1    g0598(.A(new_n729), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n434), .A2(new_n660), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n438), .B2(new_n439), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n436), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n437), .A2(new_n667), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n691), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n799), .B1(new_n806), .B2(new_n723), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n723), .B2(new_n806), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n738), .B1(new_n753), .B2(G132), .ZN(new_n809));
  INV_X1    g0609(.A(new_n751), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(new_n324), .C2(new_n747), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n762), .B1(new_n768), .B2(new_n755), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n813), .B1(new_n263), .B2(new_n766), .C1(new_n778), .C2(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT34), .Z(new_n816));
  INV_X1    g0616(.A(new_n774), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n812), .B(new_n816), .C1(G50), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(G107), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n810), .A2(G87), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n274), .B1(new_n753), .B2(G311), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n819), .A2(new_n749), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G303), .A2(new_n762), .B1(new_n768), .B2(new_n453), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  INV_X1    g0624(.A(new_n777), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n765), .A2(KEYINPUT93), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT94), .B(G283), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n822), .B(new_n826), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n735), .B1(new_n818), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n735), .A2(new_n730), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n729), .B1(new_n218), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT92), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(new_n731), .C2(new_n805), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n808), .A2(new_n838), .ZN(G384));
  NOR2_X1   g0639(.A1(new_n727), .A2(new_n205), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n660), .A4(new_n716), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n719), .A2(new_n720), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n414), .A2(new_n408), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n408), .A2(new_n660), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n406), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n408), .B(new_n660), .C1(new_n407), .C2(new_n414), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n804), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(new_n328), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n322), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n333), .A2(G68), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n318), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n317), .B1(new_n854), .B2(new_n336), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n367), .B1(new_n855), .B2(new_n658), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n350), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n352), .A2(new_n358), .ZN(new_n859));
  INV_X1    g0659(.A(new_n658), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n358), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n859), .A2(new_n861), .A3(new_n862), .A4(new_n367), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n858), .A2(KEYINPUT95), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n855), .A2(new_n658), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n361), .B2(new_n371), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT95), .B1(new_n858), .B2(new_n863), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n849), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n858), .A2(new_n863), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT95), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n866), .A4(new_n864), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n848), .A2(KEYINPUT97), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT97), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n842), .A2(new_n847), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT40), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n859), .A2(new_n861), .A3(new_n367), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n863), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n372), .B2(new_n861), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n849), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n873), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n842), .A2(new_n847), .A3(KEYINPUT40), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n877), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n442), .A2(new_n842), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT98), .ZN(new_n888));
  OAI21_X1  g0688(.A(G330), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT99), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n886), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n890), .B2(new_n889), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n691), .A2(new_n802), .B1(new_n437), .B2(new_n667), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n845), .A2(new_n846), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n869), .A2(new_n873), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n899), .A2(new_n900), .B1(new_n361), .B2(new_n658), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n883), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n414), .A2(new_n408), .A3(new_n667), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT96), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n690), .A2(new_n442), .A3(new_n692), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n654), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n840), .B1(new_n895), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n911), .B2(new_n895), .ZN(new_n913));
  INV_X1    g0713(.A(new_n526), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n914), .A2(KEYINPUT35), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(KEYINPUT35), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n915), .A2(G116), .A3(new_n215), .A4(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT36), .ZN(new_n918));
  OAI21_X1  g0718(.A(G77), .B1(new_n324), .B2(new_n244), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n243), .B1(new_n212), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(G1), .A3(new_n383), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(new_n918), .A3(new_n921), .ZN(G367));
  INV_X1    g0722(.A(new_n737), .ZN(new_n923));
  INV_X1    g0723(.A(new_n740), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n923), .B1(new_n209), .B2(new_n430), .C1(new_n924), .C2(new_n233), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n799), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT104), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n557), .A2(new_n558), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n660), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n571), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n570), .B2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n733), .B2(new_n931), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n814), .A2(new_n763), .B1(new_n825), .B2(new_n263), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G58), .B2(new_n817), .ZN(new_n934));
  XNOR2_X1  g0734(.A(KEYINPUT106), .B(G137), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n738), .B1(new_n753), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n748), .A2(G68), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n810), .A2(G77), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G50), .B2(new_n768), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n934), .B(new_n940), .C1(new_n829), .C2(new_n754), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT46), .B1(new_n817), .B2(new_n453), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n810), .A2(G97), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n274), .B1(new_n753), .B2(G317), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n942), .B(new_n946), .C1(G311), .C2(new_n762), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n947), .B1(new_n824), .B2(new_n829), .C1(new_n464), .C2(new_n778), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n768), .A2(new_n832), .B1(G107), .B2(new_n748), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT105), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n941), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n932), .B1(new_n952), .B2(new_n735), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT107), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n710), .A2(G200), .ZN(new_n955));
  INV_X1    g0755(.A(new_n533), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n956), .A3(new_n574), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n957), .A2(new_n534), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n533), .A2(new_n660), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n958), .A2(new_n959), .B1(new_n643), .B2(new_n660), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT100), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n534), .B1(new_n961), .B2(new_n634), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n667), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(new_n672), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT42), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(new_n965), .B1(KEYINPUT43), .B2(new_n931), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n670), .A2(new_n961), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n728), .B(KEYINPUT103), .Z(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n672), .B1(new_n634), .B2(new_n660), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(new_n960), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n960), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT101), .B(KEYINPUT44), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n669), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n672), .B1(new_n669), .B2(new_n671), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n664), .B(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n725), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n725), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n675), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n972), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n954), .B1(new_n970), .B2(new_n988), .ZN(G387));
  INV_X1    g0789(.A(new_n677), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n743), .A2(new_n990), .B1(new_n417), .B2(new_n674), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n237), .A2(new_n283), .ZN(new_n992));
  AOI21_X1  g0792(.A(G45), .B1(G68), .B2(G77), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n315), .A2(KEYINPUT50), .A3(new_n242), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT50), .B1(new_n315), .B2(new_n242), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n677), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n740), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n991), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n729), .B1(new_n998), .B2(new_n923), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n669), .B2(new_n733), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G77), .A2(new_n817), .B1(new_n762), .B2(G159), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G50), .A2(new_n777), .B1(new_n768), .B2(G68), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n944), .B(new_n274), .C1(new_n263), .C2(new_n752), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n565), .B2(new_n748), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n765), .A2(new_n315), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(G303), .A2(new_n768), .B1(new_n762), .B2(G322), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(new_n778), .B2(new_n1008), .C1(new_n782), .C2(new_n829), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT108), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n817), .A2(G294), .B1(new_n748), .B2(new_n832), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n738), .B1(new_n752), .B2(new_n783), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n453), .B2(new_n810), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1006), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n1022), .B2(new_n735), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n983), .B2(new_n972), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n984), .A2(new_n675), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n983), .A2(new_n725), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(G393));
  OR2_X1    g0827(.A1(new_n981), .A2(new_n984), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n984), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n664), .A2(KEYINPUT109), .A3(new_n669), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n979), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT109), .B1(new_n664), .B2(new_n669), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1028), .B(new_n675), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n740), .A2(new_n241), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n923), .B1(new_n523), .B2(new_n209), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G311), .A2(new_n777), .B1(new_n762), .B2(G317), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  NOR2_X1   g0838(.A1(new_n774), .A2(new_n831), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n274), .B1(new_n753), .B2(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n417), .B2(new_n751), .C1(new_n448), .C2(new_n747), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(G294), .C2(new_n768), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1038), .B(new_n1042), .C1(new_n464), .C2(new_n829), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G150), .A2(new_n762), .B1(new_n777), .B2(G159), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT51), .Z(new_n1045));
  AOI21_X1  g0845(.A(new_n738), .B1(new_n753), .B2(G143), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n748), .A2(G77), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n820), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n774), .A2(new_n244), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n1048), .B(new_n1049), .C1(new_n315), .C2(new_n768), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1045), .B(new_n1050), .C1(new_n242), .C2(new_n829), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n735), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n799), .B1(new_n1035), .B2(new_n1036), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n961), .B2(new_n732), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1033), .B2(new_n972), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1034), .A2(new_n1056), .ZN(G390));
  INV_X1    g0857(.A(new_n905), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n896), .B2(new_n898), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n906), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT39), .B1(new_n882), .B2(new_n873), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n685), .A2(new_n667), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(KEYINPUT82), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1064), .A2(new_n687), .A3(new_n803), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT110), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n897), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n845), .A2(KEYINPUT110), .A3(new_n846), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1069), .A3(new_n802), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n905), .B1(new_n882), .B2(new_n873), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n722), .A2(G330), .A3(new_n805), .A4(new_n897), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1062), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n903), .A2(new_n906), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1075), .A2(new_n1059), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n842), .A2(G330), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n847), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1074), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT112), .B1(new_n1080), .B2(new_n971), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1062), .A2(new_n1072), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n847), .A3(new_n1078), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT112), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1083), .A2(new_n1084), .A3(new_n972), .A4(new_n1074), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n443), .A2(new_n825), .B1(new_n763), .B2(new_n507), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G97), .B2(new_n768), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n274), .B1(new_n753), .B2(G294), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n1047), .A3(new_n811), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G87), .B2(new_n817), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1091), .C1(new_n829), .C2(new_n417), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n830), .A2(new_n935), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n774), .A2(new_n263), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT53), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n738), .B1(new_n753), .B2(G125), .ZN(new_n1096));
  INV_X1    g0896(.A(G159), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1096), .B1(new_n242), .B2(new_n751), .C1(new_n1097), .C2(new_n747), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(KEYINPUT54), .B(G143), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n768), .B2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G128), .A2(new_n762), .B1(new_n777), .B2(G132), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1093), .A2(new_n1095), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1053), .B1(new_n1092), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n729), .B1(new_n261), .B2(new_n835), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(new_n1075), .C2(new_n730), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1086), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT113), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1086), .A2(KEYINPUT113), .A3(new_n1108), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1068), .B(new_n1067), .C1(new_n1077), .C2(new_n804), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1065), .A2(new_n802), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n1073), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n898), .B1(new_n723), .B2(new_n804), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1079), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1117), .B2(new_n896), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1078), .A2(new_n442), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n910), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1083), .A2(new_n1118), .A3(new_n1074), .A4(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1115), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n896), .B1(new_n1079), .B2(new_n1116), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1080), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1125), .A3(new_n675), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT111), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1121), .A2(new_n1125), .A3(KEYINPUT111), .A4(new_n675), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1111), .A2(new_n1112), .A3(new_n1128), .A4(new_n1129), .ZN(G378));
  INV_X1    g0930(.A(new_n908), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n883), .ZN(new_n1132));
  OAI21_X1  g0932(.A(G330), .B1(new_n1132), .B2(new_n884), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n298), .A2(new_n658), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n314), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n314), .A2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n314), .A2(new_n1137), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n314), .A2(new_n1137), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n1134), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n877), .A2(new_n1133), .A3(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n848), .A2(KEYINPUT97), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n900), .A3(new_n876), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT40), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G330), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n885), .B2(new_n883), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1146), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1131), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1144), .B1(new_n877), .B2(new_n1133), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1150), .A2(new_n1152), .A3(new_n1146), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n1156), .A3(new_n908), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n972), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n753), .C2(G124), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n762), .B1(new_n777), .B2(G128), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n263), .B2(new_n747), .C1(new_n774), .C2(new_n1099), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n768), .A2(G137), .ZN(new_n1163));
  INV_X1    g0963(.A(G132), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n766), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT115), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(KEYINPUT115), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1162), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT59), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1160), .B1(new_n751), .B2(new_n754), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1169), .B2(new_n1168), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n274), .A2(G41), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n242), .B1(G33), .B2(G41), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n443), .A2(new_n763), .B1(new_n769), .B2(new_n430), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G97), .B2(new_n765), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n777), .A2(G107), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT114), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n751), .A2(new_n324), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n937), .B(new_n1172), .C1(new_n507), .C2(new_n752), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G77), .C2(new_n817), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT58), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1174), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n1183), .B2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n735), .B1(new_n1171), .B2(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT116), .Z(new_n1187));
  AOI211_X1 g0987(.A(new_n729), .B(new_n1187), .C1(new_n242), .C2(new_n835), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1146), .A2(new_n730), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1159), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1120), .B1(new_n1124), .B2(new_n1080), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1158), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n676), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT117), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1157), .A2(new_n1196), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(KEYINPUT57), .B(new_n1192), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1191), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G375));
  OR2_X1    g1002(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(new_n987), .A3(new_n1124), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1118), .A2(new_n972), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n729), .B1(new_n244), .B2(new_n835), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n274), .B1(new_n753), .B2(G303), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n938), .C1(new_n430), .C2(new_n747), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G107), .A2(new_n768), .B1(new_n762), .B2(G294), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n507), .B2(new_n825), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G97), .C2(new_n817), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n830), .A2(new_n453), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1164), .A2(new_n763), .B1(new_n769), .B2(new_n263), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n738), .B(new_n1179), .C1(G128), .C2(new_n753), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n242), .B2(new_n747), .C1(new_n1097), .C2(new_n774), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n778), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1213), .B(new_n1215), .C1(new_n1216), .C2(new_n935), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n830), .A2(new_n1100), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1211), .A2(new_n1212), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1206), .B1(new_n1053), .B2(new_n1219), .C1(new_n1069), .C2(new_n731), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1205), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1204), .A2(new_n1221), .ZN(G381));
  INV_X1    g1022(.A(G390), .ZN(new_n1223));
  INV_X1    g1023(.A(G384), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(G396), .A2(G393), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1225), .A2(G387), .A3(G381), .A4(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1111), .A2(new_n1112), .A3(new_n1126), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n1201), .A3(new_n1228), .ZN(G407));
  NAND2_X1  g1029(.A1(new_n659), .A2(G213), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT118), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1201), .A3(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(G407), .A2(new_n1232), .A3(G213), .ZN(G409));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT119), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1155), .A2(new_n1156), .A3(new_n908), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n908), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1237));
  OAI21_X1  g1037(.A(KEYINPUT117), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n971), .B1(new_n1238), .B2(new_n1198), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1235), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n972), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(KEYINPUT119), .A3(new_n1190), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1193), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n987), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1246), .A2(new_n1228), .B1(G378), .B2(new_n1201), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1124), .A2(new_n675), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT120), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1203), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1203), .A2(new_n1249), .A3(KEYINPUT60), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1248), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1221), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1224), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1252), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n1250), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G384), .B(new_n1221), .C1(new_n1257), .C2(new_n1248), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1247), .A2(new_n1231), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1234), .B1(new_n1260), .B2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1231), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1259), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1111), .A2(new_n1112), .A3(new_n1126), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1238), .A2(new_n1198), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1240), .B1(new_n1266), .B2(new_n972), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n1267), .A2(KEYINPUT119), .B1(new_n987), .B2(new_n1244), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1265), .B1(new_n1268), .B2(new_n1241), .ZN(new_n1269));
  AND2_X1   g1069(.A1(G378), .A2(new_n1201), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1263), .B(new_n1264), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1262), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1247), .A2(new_n1231), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1274), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1264), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(KEYINPUT125), .A3(new_n1272), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1261), .A2(new_n1273), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1231), .A2(G2897), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1259), .B(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT127), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G390), .B(new_n954), .C1(new_n988), .C2(new_n970), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1284), .A2(KEYINPUT123), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G396), .B(G393), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(KEYINPUT123), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1223), .A2(G387), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1284), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(KEYINPUT122), .B2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(KEYINPUT122), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1277), .A2(new_n1294), .A3(new_n1281), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT124), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n1293), .B2(KEYINPUT61), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT61), .ZN(new_n1299));
  OAI211_X1 g1099(.A(KEYINPUT124), .B(new_n1299), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT121), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1280), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1280), .A2(new_n1302), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1278), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1306));
  OR2_X1    g1106(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1301), .A2(new_n1305), .A3(new_n1306), .A4(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1296), .A2(new_n1308), .ZN(G405));
  AOI21_X1  g1109(.A(new_n1270), .B1(G375), .B2(new_n1228), .ZN(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1259), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1311), .B(new_n1293), .ZN(G402));
endmodule


