//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(KEYINPUT16), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n193), .ZN(new_n197));
  OAI211_X1 g011(.A(G146), .B(new_n189), .C1(new_n197), .C2(new_n187), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT71), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n196), .A2(new_n200), .ZN(new_n201));
  NOR3_X1   g015(.A1(new_n195), .A2(new_n199), .A3(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g017(.A(G119), .B(G128), .Z(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT24), .B(G110), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n207), .B2(G128), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n211), .B2(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G110), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n203), .A2(new_n206), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(new_n205), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n212), .B2(G110), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n194), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n198), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  INV_X1    g037(.A(G221), .ZN(new_n224));
  INV_X1    g038(.A(G234), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n224), .A2(new_n225), .A3(G953), .ZN(new_n226));
  XOR2_X1   g040(.A(new_n223), .B(new_n226), .Z(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n214), .A2(new_n221), .A3(new_n227), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G217), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(G234), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT73), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n233), .A3(new_n230), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT25), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n229), .A2(new_n240), .A3(new_n233), .A4(new_n230), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n234), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n231), .A2(new_n243), .A3(new_n235), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n237), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT9), .B(G234), .Z(new_n246));
  AOI21_X1  g060(.A(new_n224), .B1(new_n246), .B2(new_n233), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G134), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g067(.A(G137), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(G137), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n249), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT65), .B(G134), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT11), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G131), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n258), .A2(new_n259), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n249), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n252), .A2(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n250), .A2(G134), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n255), .B1(new_n267), .B2(G137), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n263), .B(new_n264), .C1(new_n249), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n261), .A2(KEYINPUT66), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n271), .B(G131), .C1(new_n257), .C2(new_n260), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G107), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(G104), .ZN(new_n275));
  INV_X1    g089(.A(G104), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G107), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(KEYINPUT74), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n274), .A2(KEYINPUT75), .A3(G104), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT74), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT3), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n279), .B2(new_n280), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G101), .ZN(new_n285));
  INV_X1    g099(.A(G101), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(new_n278), .C1(new_n282), .C2(new_n283), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(KEYINPUT4), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G143), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT64), .B1(new_n289), .B2(G146), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT64), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n217), .A3(G143), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n289), .A2(G146), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT0), .B(G128), .Z(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n217), .A2(G143), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n293), .A3(KEYINPUT0), .A4(G128), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(new_n301), .A3(new_n298), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n284), .A2(new_n304), .A3(G101), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n288), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n289), .A2(G146), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n308));
  OAI21_X1  g122(.A(G128), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n294), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n297), .A2(new_n293), .A3(new_n308), .A4(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(KEYINPUT10), .ZN(new_n313));
  OAI21_X1  g127(.A(G101), .B1(new_n277), .B2(new_n275), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n287), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n297), .A2(new_n293), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n311), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n287), .A2(new_n318), .A3(new_n314), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n320));
  AOI22_X1  g134(.A1(new_n313), .A2(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n273), .A2(new_n306), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n273), .A2(new_n306), .A3(new_n321), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n306), .A2(new_n321), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n273), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n306), .A2(new_n321), .A3(KEYINPUT79), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G110), .B(G140), .ZN(new_n334));
  INV_X1    g148(.A(G227), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(G953), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n334), .B(new_n336), .Z(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n323), .B2(new_n325), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n287), .A2(new_n314), .ZN(new_n341));
  INV_X1    g155(.A(new_n312), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n343), .B1(new_n341), .B2(new_n342), .ZN(new_n346));
  INV_X1    g160(.A(new_n319), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n340), .B1(new_n348), .B2(new_n273), .ZN(new_n349));
  INV_X1    g163(.A(new_n346), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n319), .A3(new_n344), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(KEYINPUT12), .A3(new_n330), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n333), .A2(new_n338), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G469), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NOR4_X1   g172(.A1(new_n354), .A2(G902), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n339), .A2(new_n332), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n349), .A2(new_n352), .B1(new_n323), .B2(new_n325), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(new_n337), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n355), .B1(new_n362), .B2(new_n233), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n245), .B(new_n248), .C1(new_n359), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G478), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(KEYINPUT15), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n246), .A2(G217), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G122), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT87), .B1(new_n372), .B2(G116), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT87), .ZN(new_n374));
  INV_X1    g188(.A(G116), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(G122), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n373), .A2(new_n376), .B1(G116), .B2(new_n372), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G107), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n377), .A2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n380));
  INV_X1    g194(.A(G128), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(G143), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n289), .A2(KEYINPUT88), .A3(G128), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n289), .A2(G128), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n267), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT13), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n382), .A2(KEYINPUT13), .A3(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT89), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n392), .A2(new_n393), .A3(G134), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n392), .B2(G134), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n378), .B(new_n388), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT90), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n382), .A2(KEYINPUT13), .A3(new_n383), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT13), .B1(new_n382), .B2(new_n383), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n398), .A2(new_n399), .A3(new_n385), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT89), .B1(new_n400), .B2(new_n252), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n392), .A2(new_n393), .A3(G134), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n378), .A4(new_n388), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n384), .A2(new_n386), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n258), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n387), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT91), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n372), .A2(G116), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n274), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n377), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n414), .A3(new_n387), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n410), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n371), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n416), .ZN(new_n418));
  AOI211_X1 g232(.A(new_n418), .B(new_n370), .C1(new_n397), .C2(new_n405), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n233), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT92), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n233), .C1(new_n417), .C2(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n368), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n367), .B1(new_n420), .B2(KEYINPUT92), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G214), .B1(G237), .B2(G902), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n312), .A2(G125), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n299), .B2(G125), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n431), .B(new_n433), .C1(new_n430), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G224), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT2), .B(G113), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G119), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n288), .A2(new_n305), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n375), .A2(KEYINPUT5), .A3(G119), .ZN(new_n448));
  INV_X1    g262(.A(G113), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n447), .A2(new_n450), .B1(new_n441), .B2(new_n442), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n315), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(G110), .B(G122), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n447), .A2(KEYINPUT82), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n450), .B1(new_n447), .B2(KEYINPUT82), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n444), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n315), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n341), .A2(new_n451), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n453), .B(KEYINPUT8), .Z(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n435), .A2(new_n430), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n438), .A2(new_n432), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(new_n431), .A3(new_n464), .A4(new_n433), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n439), .A2(new_n455), .A3(new_n462), .A4(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(new_n233), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n431), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(new_n438), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n446), .A2(new_n452), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n453), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n453), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(new_n475), .A3(new_n477), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n429), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n369), .A2(G952), .ZN(new_n482));
  INV_X1    g296(.A(G237), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n482), .B1(new_n225), .B2(new_n483), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n233), .B(new_n369), .C1(G234), .C2(G237), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT21), .B(G898), .Z(new_n487));
  OAI21_X1  g301(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n276), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n197), .A2(G146), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n218), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(G237), .A2(G953), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n289), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(G143), .A3(G214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n264), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(G131), .ZN(new_n501));
  OAI221_X1 g315(.A(new_n493), .B1(new_n498), .B2(new_n500), .C1(new_n501), .C2(new_n499), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT17), .ZN(new_n503));
  OAI22_X1  g317(.A1(new_n201), .A2(new_n202), .B1(new_n503), .B2(new_n501), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(new_n264), .A3(new_n497), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT85), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT85), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(new_n508), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n491), .B(new_n502), .C1(new_n504), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n501), .A2(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n194), .B1(KEYINPUT84), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n194), .B2(new_n515), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n512), .B(new_n198), .C1(G146), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n502), .ZN(new_n518));
  INV_X1    g332(.A(new_n491), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G475), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n233), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT20), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n522), .A4(new_n233), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n504), .A2(new_n510), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n491), .B1(new_n527), .B2(new_n502), .ZN(new_n528));
  INV_X1    g342(.A(new_n511), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n233), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT86), .B(G475), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n524), .A2(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n427), .A2(new_n489), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n299), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n270), .A2(new_n272), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n262), .B1(G134), .B2(new_n259), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G131), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n269), .A2(new_n312), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n270), .A2(new_n272), .A3(new_n303), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT30), .A3(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n445), .A3(new_n544), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n494), .A2(G210), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n445), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n552), .A3(new_n539), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n545), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT69), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n543), .A2(new_n552), .A3(new_n539), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n552), .B1(new_n536), .B2(new_n539), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n556), .B(KEYINPUT28), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n540), .A2(new_n445), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n553), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n553), .A2(new_n560), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT69), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n559), .B(new_n550), .C1(new_n562), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n545), .A2(new_n566), .A3(new_n551), .A4(new_n553), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n555), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT32), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n559), .B(new_n551), .C1(new_n562), .C2(new_n564), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n545), .A2(new_n550), .A3(new_n553), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT29), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n552), .B1(new_n543), .B2(new_n539), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n557), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n563), .B1(new_n577), .B2(new_n560), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n551), .A2(KEYINPUT29), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n233), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G472), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT70), .B1(new_n572), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n568), .A2(new_n569), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT32), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n569), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(KEYINPUT70), .A3(new_n586), .A4(new_n581), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n365), .B(new_n534), .C1(new_n582), .C2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n568), .A2(new_n233), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n583), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n591), .B1(new_n594), .B2(new_n364), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n592), .A2(G472), .B1(new_n568), .B2(new_n569), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n333), .A2(new_n338), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n339), .A2(new_n353), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n356), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(new_n233), .A3(new_n600), .A4(new_n357), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n353), .A2(new_n326), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(new_n338), .B1(new_n339), .B2(new_n332), .ZN(new_n603));
  OAI21_X1  g417(.A(G469), .B1(new_n603), .B2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n247), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n596), .A2(new_n605), .A3(KEYINPUT93), .A4(new_n245), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n406), .A2(new_n416), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n370), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n406), .A2(new_n416), .A3(new_n371), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(KEYINPUT33), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n611), .B1(new_n417), .B2(new_n419), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n366), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n366), .B(new_n233), .C1(new_n417), .C2(new_n419), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n366), .A2(new_n233), .ZN(new_n616));
  NOR4_X1   g430(.A1(new_n613), .A2(new_n532), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n489), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n595), .A2(new_n606), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT94), .B(KEYINPUT95), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n489), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n524), .A2(new_n627), .A3(new_n526), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n530), .A2(new_n531), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n523), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n625), .A2(new_n427), .A3(new_n626), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n481), .A2(new_n488), .A3(new_n631), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT97), .B1(new_n633), .B2(new_n426), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n595), .A3(new_n606), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  INV_X1    g452(.A(new_n605), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n222), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n235), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n242), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n534), .A3(new_n596), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  OAI21_X1  g462(.A(new_n484), .B1(new_n486), .B2(G900), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n608), .A2(new_n609), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n422), .B1(new_n651), .B2(new_n233), .ZN(new_n652));
  INV_X1    g466(.A(new_n423), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n367), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n425), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n605), .A2(new_n656), .A3(new_n481), .A4(new_n643), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n657), .B1(new_n582), .B2(new_n588), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n585), .A2(new_n586), .A3(new_n581), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT70), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n587), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT98), .A3(new_n657), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n660), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  NAND2_X1  g481(.A1(new_n585), .A2(new_n586), .ZN(new_n668));
  INV_X1    g482(.A(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n545), .A2(new_n553), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n551), .ZN(new_n671));
  AOI21_X1  g485(.A(G902), .B1(new_n577), .B2(new_n550), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n649), .B(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n639), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n675), .B1(KEYINPUT40), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n479), .A2(new_n480), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n682), .B(new_n683), .Z(new_n684));
  NAND2_X1  g498(.A1(new_n427), .A2(new_n533), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n685), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n643), .A2(new_n429), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n681), .A2(new_n684), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NAND3_X1  g504(.A1(new_n605), .A2(new_n481), .A3(new_n643), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n663), .B2(new_n587), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n617), .A2(new_n649), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  AOI21_X1  g509(.A(new_n355), .B1(new_n599), .B2(new_n233), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n359), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n248), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n664), .A2(new_n245), .A3(new_n619), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n635), .A2(new_n664), .A3(new_n245), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NAND4_X1  g518(.A1(new_n697), .A2(new_n248), .A3(new_n481), .A4(new_n643), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n427), .A2(new_n533), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n664), .A2(new_n706), .A3(new_n488), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  XNOR2_X1  g523(.A(new_n245), .B(KEYINPUT101), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n578), .A2(new_n550), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n555), .A3(new_n567), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n569), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n593), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n685), .A2(new_n698), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n625), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT102), .B(G122), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G24));
  NAND4_X1  g533(.A1(new_n617), .A2(new_n593), .A3(new_n649), .A4(new_n713), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n705), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n192), .ZN(G27));
  NOR2_X1   g536(.A1(new_n582), .A2(new_n588), .ZN(new_n723));
  INV_X1    g537(.A(new_n245), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n682), .A2(new_n429), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n605), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n727), .A2(new_n693), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n710), .A2(new_n661), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n725), .A2(new_n728), .B1(KEYINPUT42), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  AND4_X1   g546(.A1(new_n245), .A2(new_n664), .A3(new_n656), .A4(new_n727), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n252), .ZN(G36));
  NOR2_X1   g548(.A1(new_n613), .A2(new_n616), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n614), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n533), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT43), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n644), .B1(new_n738), .B2(KEYINPUT103), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n739), .B(new_n594), .C1(KEYINPUT103), .C2(new_n738), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT44), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n362), .B(KEYINPUT45), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND2_X1  g557(.A1(G469), .A2(G902), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(new_n745), .B(KEYINPUT46), .Z(new_n746));
  OAI21_X1  g560(.A(new_n248), .B1(new_n746), .B2(new_n359), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n678), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n741), .A2(new_n726), .A3(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  XNOR2_X1  g564(.A(new_n747), .B(KEYINPUT47), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n664), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n724), .A3(new_n693), .A4(new_n726), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G140), .ZN(G42));
  NAND4_X1  g568(.A1(new_n710), .A2(new_n248), .A3(new_n428), .A4(new_n737), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT104), .Z(new_n756));
  XOR2_X1   g570(.A(new_n697), .B(KEYINPUT49), .Z(new_n757));
  OR4_X1    g571(.A1(new_n684), .A2(new_n756), .A3(new_n674), .A4(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n699), .A2(new_n726), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT112), .Z(new_n760));
  INV_X1    g574(.A(new_n484), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n738), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT113), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n643), .A3(new_n714), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n247), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n751), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n738), .A2(new_n761), .A3(new_n715), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n768), .A2(new_n726), .A3(new_n769), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n684), .A2(new_n698), .A3(new_n428), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n769), .ZN(new_n773));
  XOR2_X1   g587(.A(new_n773), .B(KEYINPUT50), .Z(new_n774));
  AND3_X1   g588(.A1(new_n764), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n760), .A2(new_n245), .A3(new_n761), .A4(new_n675), .ZN(new_n776));
  INV_X1    g590(.A(new_n736), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n776), .A2(new_n533), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n770), .A2(KEYINPUT114), .A3(new_n774), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n780), .A4(new_n778), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n782), .A2(new_n482), .A3(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n721), .B1(new_n692), .B2(new_n693), .ZN(new_n786));
  INV_X1    g600(.A(new_n481), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n685), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n605), .A2(new_n644), .A3(new_n649), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n674), .B(new_n788), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n664), .A2(KEYINPUT98), .A3(new_n657), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT98), .B1(new_n664), .B2(new_n657), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n786), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT52), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n666), .A2(new_n798), .A3(new_n786), .A4(new_n793), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n703), .A2(new_n708), .A3(new_n700), .A4(new_n717), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(new_n731), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT105), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n654), .B2(new_n655), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n424), .A2(KEYINPUT105), .A3(new_n425), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n532), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n618), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n625), .A3(new_n595), .A4(new_n606), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n589), .A3(new_n646), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n808), .A2(new_n589), .A3(KEYINPUT106), .A4(new_n646), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n645), .ZN(new_n814));
  INV_X1    g628(.A(new_n650), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n654), .A2(new_n803), .A3(new_n655), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT105), .B1(new_n424), .B2(new_n425), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n664), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n814), .B1(new_n820), .B2(new_n720), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n733), .B1(new_n821), .B2(new_n726), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n813), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n785), .B1(new_n802), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT108), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n802), .A2(new_n785), .A3(new_n823), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n769), .A2(new_n481), .A3(new_n699), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n650), .B(new_n818), .C1(new_n663), .C2(new_n587), .ZN(new_n832));
  INV_X1    g646(.A(new_n720), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n645), .B(new_n726), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n733), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n811), .B2(new_n812), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n799), .A2(new_n731), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n813), .A2(new_n838), .A3(new_n822), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n800), .B1(new_n796), .B2(KEYINPUT52), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n824), .B(new_n829), .C1(new_n839), .C2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n784), .A2(new_n830), .A3(new_n831), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n776), .A2(new_n618), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n763), .A2(new_n729), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT115), .Z(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT48), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(G952), .A2(G953), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n758), .B1(new_n850), .B2(new_n851), .ZN(G75));
  OAI21_X1  g666(.A(new_n824), .B1(new_n839), .B2(new_n843), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(G210), .A3(G902), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n853), .A2(new_n857), .A3(G210), .A4(G902), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n474), .A2(new_n472), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(new_n469), .Z(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(KEYINPUT117), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT117), .B1(new_n859), .B2(new_n862), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n867));
  INV_X1    g681(.A(new_n862), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n854), .A2(new_n856), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n369), .A2(G952), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n866), .A2(new_n867), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n869), .B(new_n871), .C1(new_n864), .C2(new_n865), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(G51));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n844), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n853), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n744), .B(KEYINPUT57), .Z(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT120), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n879), .A2(new_n884), .A3(new_n880), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n876), .B1(new_n886), .B2(new_n599), .ZN(new_n887));
  AOI211_X1 g701(.A(KEYINPUT121), .B(new_n354), .C1(new_n883), .C2(new_n885), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n853), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n233), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n743), .B(KEYINPUT122), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n870), .B1(new_n889), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(new_n521), .Z(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n870), .ZN(G60));
  NAND2_X1  g711(.A1(new_n610), .A2(new_n612), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n830), .A2(new_n844), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n616), .B(KEYINPUT59), .Z(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n899), .A2(new_n879), .A3(new_n880), .A4(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n870), .A3(new_n903), .ZN(G63));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n905));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n890), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n870), .B1(new_n908), .B2(new_n641), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n231), .B2(new_n908), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n911), .B(new_n912), .Z(G66));
  INV_X1    g727(.A(new_n487), .ZN(new_n914));
  OAI21_X1  g728(.A(G953), .B1(new_n914), .B2(new_n437), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n800), .B1(new_n811), .B2(new_n812), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n860), .B1(G898), .B2(new_n369), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  NAND2_X1  g733(.A1(new_n542), .A2(new_n544), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n516), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n369), .A2(G900), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT126), .ZN(new_n925));
  INV_X1    g739(.A(new_n731), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n741), .A2(new_n726), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n729), .A2(new_n788), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(new_n748), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n666), .A2(new_n786), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n835), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n930), .A2(new_n753), .A3(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n923), .B(new_n925), .C1(new_n934), .C2(G953), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n689), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT62), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n723), .A2(new_n724), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n938), .A2(new_n677), .A3(new_n727), .A4(new_n807), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n749), .A2(new_n937), .A3(new_n753), .A4(new_n939), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n940), .A2(G953), .A3(new_n923), .ZN(new_n941));
  INV_X1    g755(.A(G900), .ZN(new_n942));
  OAI21_X1  g756(.A(G953), .B1(new_n335), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n935), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(G72));
  NAND2_X1  g761(.A1(new_n934), .A2(new_n916), .ZN(new_n948));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  AOI21_X1  g764(.A(new_n574), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n940), .A2(new_n916), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n671), .B1(new_n952), .B2(new_n950), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n671), .A2(new_n574), .A3(new_n950), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n828), .A2(new_n954), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n951), .A2(new_n953), .A3(new_n870), .A4(new_n955), .ZN(G57));
endmodule


