//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n542, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g037(.A1(new_n459), .A2(KEYINPUT66), .A3(G101), .A4(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n459), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n459), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n475), .A2(new_n459), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n459), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n475), .A2(new_n493), .A3(G138), .A4(new_n459), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT67), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n503), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n498), .A2(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(KEYINPUT68), .B1(G89), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n507), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n520), .A3(new_n524), .ZN(G286));
  INV_X1    g100(.A(G286), .ZN(G168));
  AOI22_X1  g101(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n502), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n507), .A2(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n510), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G171));
  XOR2_X1   g107(.A(KEYINPUT69), .B(G81), .Z(new_n533));
  AOI22_X1  g108(.A1(new_n517), .A2(new_n533), .B1(new_n507), .B2(G43), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n502), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n534), .B(KEYINPUT70), .C1(new_n502), .C2(new_n535), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G188));
  NAND2_X1  g121(.A1(new_n509), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT9), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n507), .A2(new_n550), .A3(G53), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  AND3_X1   g128(.A1(KEYINPUT67), .A2(KEYINPUT5), .A3(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(G543), .B1(KEYINPUT67), .B2(KEYINPUT5), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(G91), .B2(new_n517), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n552), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  NAND2_X1  g136(.A1(new_n517), .A2(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n507), .A2(G49), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  NAND3_X1  g140(.A1(new_n507), .A2(KEYINPUT71), .A3(G48), .ZN(new_n566));
  INV_X1    g141(.A(new_n506), .ZN(new_n567));
  NOR2_X1   g142(.A1(KEYINPUT6), .A2(G651), .ZN(new_n568));
  OAI211_X1 g143(.A(G48), .B(G543), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT71), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n556), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n517), .A2(G86), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n502), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n510), .A2(new_n581), .B1(new_n547), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  INV_X1    g162(.A(G92), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n510), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n589), .A2(new_n590), .B1(G54), .B2(new_n507), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n556), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT72), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n596), .B(new_n592), .C1(new_n556), .C2(new_n593), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(G651), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n586), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n586), .B1(new_n600), .B2(G868), .ZN(G321));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g178(.A(G297), .B(KEYINPUT73), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n600), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n480), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(G2100), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n613), .B2(new_n612), .ZN(new_n616));
  OR3_X1    g191(.A1(new_n616), .A2(new_n614), .A3(G2100), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n614), .B2(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n480), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n459), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(G156));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2427), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n626), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n629), .B2(new_n628), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G14), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n636), .A2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(G401));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT75), .Z(new_n644));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n644), .B(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n642), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n647), .B(new_n648), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n642), .A2(new_n648), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT78), .B(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n662), .A2(new_n665), .A3(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1986), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT79), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G27), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n492), .A2(new_n494), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n486), .A2(new_n489), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n682), .B1(new_n685), .B2(G29), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2078), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(G35), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G162), .B2(new_n680), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT29), .Z(new_n690));
  INV_X1    g265(.A(G2090), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n680), .A2(G33), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT25), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n475), .A2(G127), .ZN(new_n696));
  NAND2_X1  g271(.A1(G115), .A2(G2104), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n459), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g273(.A(new_n695), .B(new_n698), .C1(G139), .C2(new_n480), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n693), .B1(new_n699), .B2(new_n680), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT88), .B(G2072), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n680), .A2(G32), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n465), .A2(G2105), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n480), .A2(G141), .B1(G105), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT26), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n477), .B2(G129), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n704), .B1(new_n711), .B2(new_n680), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n703), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G34), .ZN(new_n716));
  AOI21_X1  g291(.A(G29), .B1(new_n716), .B2(KEYINPUT24), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(KEYINPUT24), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G160), .B2(G29), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n712), .A2(new_n714), .B1(G2084), .B2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT30), .B(G28), .ZN(new_n722));
  OR2_X1    g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  NAND2_X1  g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n722), .A2(new_n680), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(new_n623), .B2(new_n680), .ZN(new_n726));
  INV_X1    g301(.A(new_n720), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  NOR4_X1   g305(.A1(new_n692), .A2(new_n702), .A3(new_n715), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT89), .B(G1966), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NOR2_X1   g313(.A1(G171), .A2(new_n732), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G5), .B2(new_n732), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n738), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n734), .A2(new_n736), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT90), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n731), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n732), .A2(G19), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n540), .B2(new_n732), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT84), .B(G1341), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT83), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n599), .B2(new_n732), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1348), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n690), .A2(new_n691), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT92), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n680), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(G104), .A2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT85), .Z(new_n763));
  INV_X1    g338(.A(G128), .ZN(new_n764));
  INV_X1    g339(.A(G140), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n764), .A2(new_n476), .B1(new_n479), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT86), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n760), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2067), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n732), .A2(G20), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT23), .Z(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n755), .A2(new_n757), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n732), .A2(G22), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n732), .ZN(new_n777));
  INV_X1    g352(.A(G1971), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G6), .A2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G305), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n780), .B1(new_n781), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n786));
  OR2_X1    g361(.A1(G288), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(G288), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G16), .B2(G23), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n792), .A2(new_n794), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n785), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT34), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n785), .B(new_n799), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n477), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n480), .A2(G131), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n459), .A2(G107), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n807), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G24), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n584), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1986), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n800), .A2(new_n801), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n801), .B1(new_n800), .B2(new_n814), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n798), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n818), .A2(KEYINPUT82), .A3(KEYINPUT36), .ZN(new_n819));
  NAND2_X1  g394(.A1(KEYINPUT82), .A2(KEYINPUT36), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n798), .B(new_n820), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n775), .B1(new_n819), .B2(new_n821), .ZN(G311));
  XNOR2_X1  g397(.A(G311), .B(KEYINPUT93), .ZN(G150));
  AOI22_X1  g398(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n502), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n507), .A2(G55), .ZN(new_n826));
  INV_X1    g401(.A(G93), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n510), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT37), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n599), .A2(new_n605), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n538), .B2(new_n539), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n536), .A2(new_n825), .A3(new_n828), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n835), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n830), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n832), .B1(new_n841), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n768), .B(new_n685), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n806), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n699), .B(new_n710), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n477), .A2(G130), .B1(new_n480), .B2(G142), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT95), .B1(new_n459), .B2(G118), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n459), .A2(KEYINPUT95), .A3(G118), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n612), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n846), .B(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n845), .B(new_n857), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n623), .B(new_n484), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(G160), .Z(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n858), .A2(KEYINPUT97), .A3(new_n860), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n845), .B(new_n857), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n861), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g443(.A1(new_n584), .A2(KEYINPUT98), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n584), .A2(KEYINPUT98), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n790), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n789), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n781), .B(G303), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(KEYINPUT99), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(new_n876), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n838), .B(new_n607), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n599), .A2(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n599), .A2(G299), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(KEYINPUT41), .A3(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n881), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G868), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(G868), .B2(new_n829), .ZN(G295));
  OAI21_X1  g470(.A(new_n894), .B1(G868), .B2(new_n829), .ZN(G331));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  INV_X1    g472(.A(new_n880), .ZN(new_n898));
  NAND2_X1  g473(.A1(G171), .A2(KEYINPUT100), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n528), .B2(new_n531), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(G286), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(G286), .A3(new_n901), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n838), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n906), .A2(new_n902), .B1(new_n836), .B2(new_n837), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n838), .A3(KEYINPUT102), .A4(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n886), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n905), .A2(new_n907), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(KEYINPUT101), .A3(new_n889), .A4(new_n890), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT101), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n905), .A2(new_n907), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n916), .B2(new_n891), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n898), .A2(new_n912), .A3(new_n914), .A4(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI22_X1  g495(.A1(new_n911), .A2(new_n891), .B1(new_n885), .B2(new_n913), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n880), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n917), .A2(new_n914), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n923), .A2(KEYINPUT103), .A3(new_n898), .A4(new_n912), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT104), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n920), .A2(new_n924), .A3(new_n927), .A4(new_n922), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n897), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n923), .A2(new_n912), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n920), .B(new_n924), .C1(new_n930), .C2(new_n898), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(new_n897), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT44), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(KEYINPUT43), .B2(new_n925), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n937), .ZN(G397));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(G164), .B2(G1384), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n471), .A2(new_n472), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G2105), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(G40), .A3(new_n469), .A4(new_n464), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n768), .B(G2067), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n710), .ZN(new_n946));
  INV_X1    g521(.A(new_n944), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(G1996), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT46), .Z(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n945), .A2(new_n944), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(G1996), .A3(new_n710), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n806), .A2(new_n809), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n806), .A2(new_n809), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n944), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n948), .A2(new_n711), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT105), .Z(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n947), .A2(G1986), .A3(G290), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT126), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT48), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n952), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n958), .A3(new_n961), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n768), .A2(G2067), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n947), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n971));
  INV_X1    g546(.A(G1956), .ZN(new_n972));
  INV_X1    g547(.A(G40), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n470), .A2(new_n473), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n683), .B2(new_n684), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n558), .A2(G651), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n517), .A2(G91), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n981), .A2(KEYINPUT112), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(G299), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n552), .B(new_n559), .C1(KEYINPUT112), .C2(KEYINPUT57), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n685), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT56), .B(G2072), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n940), .A2(new_n988), .A3(new_n974), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n979), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n979), .A2(new_n986), .A3(new_n993), .A4(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n979), .A2(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(new_n986), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT61), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT114), .B(G1996), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n940), .A2(new_n988), .A3(new_n974), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n975), .A2(new_n974), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT58), .B(G1341), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n540), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT59), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT59), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1008), .A3(new_n540), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n991), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n971), .B1(new_n999), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT61), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n996), .B2(new_n997), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n991), .A2(new_n1015), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n992), .A2(new_n994), .B1(new_n997), .B2(new_n996), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1016), .B(KEYINPUT115), .C1(KEYINPUT61), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1002), .A2(G2067), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n685), .A2(new_n987), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n943), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  NOR4_X1   g596(.A1(G164), .A2(KEYINPUT107), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1023), .B1(new_n975), .B2(new_n976), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1019), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT60), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n600), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n599), .B1(new_n1027), .B2(KEYINPUT60), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1029), .A2(new_n1030), .B1(KEYINPUT60), .B2(new_n1027), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1013), .A2(new_n1018), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n998), .B1(new_n1027), .B2(new_n599), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n995), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(KEYINPUT116), .A3(new_n1034), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1021), .B(new_n728), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n940), .A2(new_n988), .A3(new_n974), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n735), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G286), .A2(G8), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT119), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1039), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT120), .B(new_n1039), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1044), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1044), .B2(new_n1053), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1049), .A2(new_n1050), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1045), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT117), .Z(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n503), .B2(new_n512), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1042), .A2(new_n778), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n975), .A2(new_n976), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n691), .A4(new_n974), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(G8), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1025), .B2(G2090), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(G8), .A3(new_n1062), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(KEYINPUT111), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n977), .A2(new_n978), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1072), .A2(new_n691), .B1(new_n1042), .B2(new_n778), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT111), .B(new_n1061), .C1(new_n1073), .C2(new_n1040), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n787), .A2(G1976), .A3(new_n788), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT108), .B1(new_n1002), .B2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT108), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1077), .B(new_n1040), .C1(new_n975), .C2(new_n974), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n943), .A2(G164), .A3(G1384), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1077), .B1(new_n1080), .B2(new_n1040), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1002), .A2(KEYINPUT108), .A3(G8), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n575), .A2(G651), .B1(G86), .B2(new_n517), .ZN(new_n1084));
  INV_X1    g659(.A(G1981), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n572), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1084), .B2(new_n572), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT49), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G305), .A2(G1981), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1084), .A2(new_n1085), .A3(new_n572), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g668(.A1(KEYINPUT52), .A2(new_n1079), .B1(new_n1083), .B2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT109), .B(G1976), .Z(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT52), .B1(G288), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1083), .A2(new_n1075), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1074), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1071), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n940), .A2(new_n988), .A3(new_n1101), .A4(new_n974), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1025), .A2(new_n738), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1104), .A2(new_n1106), .A3(G171), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1100), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1103), .B(new_n1105), .C1(KEYINPUT123), .C2(G301), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(KEYINPUT54), .ZN(new_n1113));
  AND4_X1   g688(.A1(new_n1059), .A2(new_n1099), .A3(new_n1109), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1037), .A2(new_n1038), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT110), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1079), .A2(KEYINPUT52), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1083), .A2(new_n1093), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1097), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(new_n1070), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G288), .A2(G1976), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1086), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1083), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  OAI221_X1 g700(.A(KEYINPUT110), .B1(new_n1122), .B2(new_n1123), .C1(new_n1070), .C2(new_n1119), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1044), .A2(G168), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n1099), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1070), .A2(KEYINPUT63), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1062), .B1(new_n1069), .B2(G8), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1044), .A2(G168), .ZN(new_n1132));
  NOR4_X1   g707(.A1(new_n1130), .A2(new_n1119), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1059), .B2(KEYINPUT62), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1115), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n584), .B(G1986), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n944), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n956), .A2(new_n1141), .A3(new_n959), .A4(new_n961), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT124), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT124), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1145), .B(new_n1142), .C1(new_n1115), .C2(new_n1138), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n970), .B1(new_n1144), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g722(.A(G319), .B1(new_n639), .B2(new_n640), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G227), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g724(.A(new_n1150), .B(KEYINPUT127), .ZN(new_n1151));
  NOR2_X1   g725(.A1(G229), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g726(.A1(new_n1152), .A2(new_n867), .A3(new_n935), .ZN(G225));
  INV_X1    g727(.A(G225), .ZN(G308));
endmodule


