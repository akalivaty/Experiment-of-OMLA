//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G113), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  AOI22_X1  g010(.A1(new_n192), .A2(new_n195), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT3), .A3(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT81), .B1(new_n201), .B2(G104), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n199), .A3(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n204), .A3(new_n205), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT83), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n199), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n201), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND3_X1   g026(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n208), .B2(new_n212), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n197), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G110), .B(G122), .ZN(new_n216));
  INV_X1    g030(.A(new_n193), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT2), .B(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n196), .A2(new_n193), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  INV_X1    g036(.A(new_n203), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n205), .A2(new_n207), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n222), .B(G101), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n205), .A2(new_n207), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n204), .B1(new_n227), .B2(new_n203), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n221), .B(new_n225), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n215), .A2(new_n216), .A3(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G953), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G224), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT7), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n234), .A2(G146), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  OAI21_X1  g050(.A(G128), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G143), .ZN(new_n240));
  AOI21_X1  g054(.A(G146), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G143), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n234), .A2(KEYINPUT65), .A3(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n237), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n235), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n240), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n248), .B(new_n250), .C1(new_n251), .C2(new_n243), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G125), .ZN(new_n254));
  INV_X1    g068(.A(G125), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n241), .B2(new_n246), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n248), .C1(new_n251), .C2(new_n243), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n233), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT64), .B(G143), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n244), .B(new_n245), .C1(new_n264), .C2(G146), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n235), .B1(new_n264), .B2(G146), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n265), .A2(new_n237), .B1(new_n266), .B2(new_n250), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n255), .ZN(new_n268));
  INV_X1    g082(.A(new_n262), .ZN(new_n269));
  INV_X1    g083(.A(new_n233), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n230), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n216), .B(KEYINPUT8), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n192), .B1(new_n275), .B2(new_n217), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n220), .B(new_n276), .C1(new_n213), .C2(new_n214), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n189), .A2(new_n191), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(G113), .A3(new_n195), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n220), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n208), .A2(new_n212), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n274), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n187), .B1(new_n272), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n216), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n281), .A2(KEYINPUT83), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n280), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n226), .A2(new_n228), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n225), .A2(new_n221), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n288), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT6), .A3(new_n230), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n254), .A2(new_n262), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n232), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT6), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n288), .C1(new_n291), .C2(new_n294), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT85), .B(new_n187), .C1(new_n272), .C2(new_n283), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n286), .A2(new_n287), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT86), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n301), .A2(new_n302), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(KEYINPUT86), .A3(new_n287), .A4(new_n286), .ZN(new_n307));
  INV_X1    g121(.A(new_n287), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n277), .A2(new_n282), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n273), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n263), .A2(new_n271), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n230), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT85), .B1(new_n313), .B2(new_n187), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n305), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G140), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT79), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT80), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n231), .A2(G227), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT82), .B1(new_n241), .B2(new_n236), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(KEYINPUT1), .C1(new_n264), .C2(G146), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(G128), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n266), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n252), .ZN(new_n331));
  INV_X1    g145(.A(new_n281), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT10), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT10), .B(new_n253), .C1(new_n213), .C2(new_n214), .ZN(new_n334));
  OAI21_X1  g148(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n260), .A2(new_n261), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(new_n225), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT11), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g156(.A(G134), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(G137), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(G137), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT11), .ZN(new_n349));
  INV_X1    g163(.A(G137), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G134), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G131), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(G134), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n342), .B2(new_n344), .ZN(new_n355));
  INV_X1    g169(.A(G131), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n348), .A2(KEYINPUT11), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n349), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n353), .A2(KEYINPUT68), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT68), .B1(new_n353), .B2(new_n359), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n333), .A2(new_n340), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n289), .A2(new_n290), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n267), .A2(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n225), .A2(new_n261), .A3(new_n260), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n365), .A2(new_n367), .B1(new_n368), .B2(new_n336), .ZN(new_n369));
  INV_X1    g183(.A(new_n252), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n370), .B1(new_n328), .B2(new_n329), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n371), .B2(new_n281), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n362), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n324), .B1(new_n364), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(new_n362), .A3(new_n372), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n289), .A2(new_n267), .A3(new_n290), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n371), .B2(new_n281), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT12), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n353), .A2(new_n359), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT12), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n331), .A2(new_n332), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(new_n376), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n375), .B(new_n323), .C1(new_n378), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n374), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n187), .ZN(new_n386));
  NAND2_X1  g200(.A1(G469), .A2(G902), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n378), .A2(new_n382), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n324), .B1(new_n388), .B2(new_n364), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n375), .A2(new_n323), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n363), .B1(new_n333), .B2(new_n340), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n392), .A3(G469), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n264), .A2(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n249), .A2(G143), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(KEYINPUT13), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT13), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n264), .A2(new_n398), .A3(G128), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(G134), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n343), .A3(new_n396), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G116), .B(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n201), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n395), .A2(KEYINPUT90), .A3(new_n343), .A4(new_n396), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n400), .A2(new_n403), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G122), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G116), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n201), .B1(new_n409), .B2(KEYINPUT14), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n404), .ZN(new_n411));
  INV_X1    g225(.A(new_n401), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n343), .B1(new_n395), .B2(new_n396), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT9), .B(G234), .ZN(new_n415));
  INV_X1    g229(.A(G217), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(G953), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n407), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n417), .B1(new_n407), .B2(new_n414), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n187), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G478), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT15), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n187), .B1(KEYINPUT15), .B2(new_n421), .C1(new_n418), .C2(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(G234), .A2(G237), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n425), .A2(G952), .A3(new_n231), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G902), .A3(G953), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT91), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(G898), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n423), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G237), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n231), .A3(G214), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n238), .A3(new_n240), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n433), .A2(new_n231), .A3(G143), .A4(G214), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n356), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n436), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(G131), .ZN(new_n441));
  AOI211_X1 g255(.A(KEYINPUT87), .B(new_n356), .C1(new_n435), .C2(new_n436), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n437), .B(new_n438), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(G131), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT87), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n439), .A3(G131), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G140), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n255), .A2(G140), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT16), .ZN(new_n451));
  OR3_X1    g265(.A1(new_n255), .A2(KEYINPUT16), .A3(G140), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n243), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(G146), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n443), .A2(new_n447), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n199), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n440), .A2(KEYINPUT18), .A3(G131), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT18), .A2(G131), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n435), .A2(new_n436), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G125), .B(G140), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n243), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n458), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n460), .B1(new_n458), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n187), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G475), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT88), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(new_n437), .C1(new_n441), .C2(new_n442), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT89), .A2(KEYINPUT19), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n464), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n455), .B1(new_n480), .B2(G146), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n474), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n460), .B1(new_n483), .B2(new_n466), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n471), .B(new_n472), .C1(new_n484), .C2(new_n467), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n458), .A2(new_n460), .A3(new_n466), .ZN(new_n487));
  INV_X1    g301(.A(new_n466), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n481), .B1(new_n473), .B2(KEYINPUT88), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n489), .B2(new_n476), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n487), .B1(new_n490), .B2(new_n460), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n471), .B1(new_n491), .B2(new_n472), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n432), .B(new_n470), .C1(new_n486), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n415), .B2(G902), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n394), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n318), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n338), .B1(new_n360), .B2(new_n361), .ZN(new_n498));
  INV_X1    g312(.A(new_n221), .ZN(new_n499));
  OAI21_X1  g313(.A(G131), .B1(new_n344), .B2(new_n354), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n253), .A2(new_n359), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n433), .A2(new_n231), .A3(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT27), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G101), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT29), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n359), .A2(new_n500), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT69), .B1(new_n267), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n253), .A2(new_n514), .A3(new_n359), .A4(new_n500), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT68), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n346), .A2(new_n352), .A3(G131), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n356), .B1(new_n355), .B2(new_n358), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n353), .A2(KEYINPUT68), .A3(new_n359), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n337), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n221), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n498), .A2(new_n499), .A3(new_n513), .A4(new_n515), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT72), .B1(new_n525), .B2(KEYINPUT28), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n504), .B(new_n511), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT30), .B1(new_n516), .B2(new_n522), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n257), .A2(new_n258), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n244), .A2(new_n245), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n239), .A2(G143), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n234), .A2(KEYINPUT64), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n243), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n532), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n256), .B(new_n235), .C1(new_n264), .C2(G146), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n260), .A2(KEYINPUT66), .A3(new_n261), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n379), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n501), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n499), .B1(new_n530), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n516), .A2(new_n522), .A3(new_n221), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n509), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n501), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n221), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n548), .A2(new_n524), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n504), .B1(new_n549), .B2(new_n503), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n508), .B(KEYINPUT71), .Z(new_n551));
  OAI211_X1 g365(.A(new_n546), .B(new_n510), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n529), .A2(new_n552), .A3(new_n187), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G472), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n524), .A2(new_n508), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n530), .A2(new_n543), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n221), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT31), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n550), .A2(new_n551), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n545), .A2(new_n509), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n541), .A2(new_n542), .A3(new_n501), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n498), .A2(new_n513), .A3(new_n515), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n562), .B1(KEYINPUT30), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT70), .B(new_n561), .C1(new_n564), .C2(new_n499), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n544), .B2(new_n556), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT31), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(G472), .A2(G902), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n555), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  AOI211_X1 g386(.A(KEYINPUT32), .B(new_n572), .C1(new_n560), .C2(new_n568), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n554), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n231), .A2(G221), .A3(G234), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT76), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n249), .A2(G119), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n190), .A2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT24), .B(G110), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n249), .A2(G119), .B1(KEYINPUT74), .B2(KEYINPUT23), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT74), .B(KEYINPUT23), .Z(new_n586));
  XNOR2_X1  g400(.A(G119), .B(G128), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n583), .B1(new_n588), .B2(G110), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n464), .A2(new_n243), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n455), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n584), .B1(new_n581), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n595));
  OAI21_X1  g409(.A(G110), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI211_X1 g410(.A(KEYINPUT75), .B(new_n584), .C1(new_n581), .C2(new_n593), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT73), .B1(new_n581), .B2(new_n582), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT24), .B(G110), .Z(new_n600));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n587), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n455), .ZN(new_n603));
  AOI21_X1  g417(.A(G146), .B1(new_n451), .B2(new_n452), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n599), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n592), .B1(new_n598), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n578), .B1(new_n606), .B2(KEYINPUT77), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(KEYINPUT77), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n602), .A2(new_n599), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n609), .B(new_n456), .C1(new_n596), .C2(new_n597), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT77), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n592), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n607), .B1(new_n613), .B2(new_n578), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n416), .B1(G234), .B2(new_n187), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G902), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT78), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n610), .A2(new_n611), .A3(new_n592), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n611), .B1(new_n610), .B2(new_n592), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n578), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n607), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n187), .A3(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n620), .B1(new_n629), .B2(new_n616), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n497), .A2(new_n574), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  NAND2_X1  g446(.A1(new_n394), .A2(new_n495), .ZN(new_n633));
  INV_X1    g447(.A(new_n630), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n572), .B1(new_n560), .B2(new_n568), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n565), .A2(new_n567), .A3(KEYINPUT31), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n558), .A2(new_n559), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n503), .B1(new_n548), .B2(new_n524), .ZN(new_n639));
  INV_X1    g453(.A(new_n504), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n551), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n187), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n636), .B1(new_n643), .B2(G472), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n635), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n317), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n315), .B2(new_n303), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n470), .B1(new_n486), .B2(new_n492), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n407), .A2(new_n414), .A3(new_n417), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT92), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(KEYINPUT33), .C1(new_n418), .C2(new_n419), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n407), .A2(new_n414), .ZN(new_n652));
  INV_X1    g466(.A(new_n417), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n654), .B(new_n649), .C1(KEYINPUT92), .C2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(G478), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n421), .A2(new_n187), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n654), .B2(new_n649), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n659), .B2(new_n421), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n648), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n430), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n645), .A2(new_n647), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  NAND2_X1  g480(.A1(new_n423), .A2(new_n424), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n667), .B(new_n470), .C1(new_n486), .C2(new_n492), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n430), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n645), .A2(new_n647), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G107), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  AOI21_X1  g487(.A(KEYINPUT25), .B1(new_n614), .B2(new_n187), .ZN(new_n674));
  INV_X1    g488(.A(new_n628), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n616), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n606), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n618), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n497), .A2(new_n644), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT37), .B(G110), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT94), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G12));
  INV_X1    g498(.A(G900), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n426), .B1(new_n428), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n423), .B2(new_n424), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n470), .B(new_n687), .C1(new_n486), .C2(new_n492), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n647), .A2(new_n689), .A3(new_n680), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n633), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n574), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT95), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n574), .A2(new_n691), .A3(KEYINPUT95), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  INV_X1    g511(.A(new_n633), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n686), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  XOR2_X1   g516(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n316), .B(new_n703), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n570), .B1(new_n637), .B2(new_n642), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT32), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n636), .A2(new_n555), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n565), .A2(new_n567), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n525), .A2(new_n551), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n187), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G472), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n648), .A2(new_n667), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n680), .A3(new_n646), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n702), .A2(new_n704), .A3(new_n713), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n251), .ZN(G45));
  INV_X1    g531(.A(new_n679), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n629), .B2(new_n616), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n708), .B2(new_n554), .ZN(new_n720));
  INV_X1    g534(.A(new_n686), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n648), .A2(new_n661), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(KEYINPUT98), .A3(new_n647), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT98), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n315), .A2(new_n303), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n317), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n725), .B1(new_n727), .B2(new_n722), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n633), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n720), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  INV_X1    g545(.A(KEYINPUT99), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n706), .A2(new_n707), .B1(G472), .B2(new_n553), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n385), .B1(new_n384), .B2(new_n187), .ZN(new_n734));
  AOI211_X1 g548(.A(G469), .B(G902), .C1(new_n374), .C2(new_n383), .ZN(new_n735));
  INV_X1    g549(.A(new_n495), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n663), .A2(new_n737), .A3(new_n630), .A4(new_n647), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n732), .B1(new_n733), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n657), .A2(new_n660), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n472), .B1(new_n484), .B2(new_n467), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT20), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n485), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n740), .B1(new_n743), .B2(new_n470), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n647), .A2(new_n744), .A3(new_n431), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n378), .A2(new_n382), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n391), .A2(new_n375), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n746), .A2(new_n390), .B1(new_n747), .B2(new_n324), .ZN(new_n748));
  OAI21_X1  g562(.A(G469), .B1(new_n748), .B2(G902), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n630), .A2(new_n749), .A3(new_n495), .A4(new_n386), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n574), .A2(new_n751), .A3(KEYINPUT99), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n739), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND2_X1  g569(.A1(new_n669), .A2(new_n647), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n750), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n574), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g572(.A(KEYINPUT100), .B(G116), .Z(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G18));
  NAND3_X1  g574(.A1(new_n749), .A2(new_n495), .A3(new_n386), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n727), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n719), .A2(new_n493), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n574), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G119), .ZN(G21));
  NAND2_X1  g579(.A1(new_n525), .A2(KEYINPUT28), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT72), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n640), .B1(new_n768), .B2(new_n526), .ZN(new_n769));
  INV_X1    g583(.A(new_n551), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n568), .B(new_n638), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI22_X1  g585(.A1(G472), .A2(new_n643), .B1(new_n771), .B2(new_n570), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT101), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n630), .A2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n616), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n627), .B2(new_n628), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT101), .B1(new_n776), .B2(new_n620), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n727), .A2(new_n714), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n761), .A2(new_n430), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n772), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  XNOR2_X1  g596(.A(new_n722), .B(KEYINPUT102), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n680), .A3(new_n762), .A4(new_n772), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  INV_X1    g599(.A(new_n778), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n733), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n286), .A2(new_n301), .A3(new_n302), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n646), .B1(new_n788), .B2(new_n308), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n305), .A3(new_n307), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n633), .A2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n783), .A2(KEYINPUT42), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n783), .A2(new_n574), .A3(new_n630), .A4(new_n791), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n787), .A2(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n356), .ZN(G33));
  NAND4_X1  g610(.A1(new_n574), .A2(new_n630), .A3(new_n689), .A4(new_n791), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NAND3_X1  g612(.A1(new_n743), .A2(new_n661), .A3(new_n470), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT43), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT103), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT104), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n644), .B2(new_n719), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n644), .A2(new_n802), .A3(new_n719), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT44), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n790), .ZN(new_n808));
  AOI21_X1  g622(.A(KEYINPUT45), .B1(new_n389), .B2(new_n392), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n385), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT46), .B1(new_n812), .B2(new_n387), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n735), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(KEYINPUT46), .A3(new_n387), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n736), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n700), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n805), .A2(new_n806), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n807), .A2(new_n808), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  XNOR2_X1  g634(.A(new_n816), .B(KEYINPUT47), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n790), .A2(new_n630), .A3(new_n722), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n733), .A3(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  AND3_X1   g638(.A1(new_n574), .A2(new_n751), .A3(KEYINPUT99), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT99), .B1(new_n574), .B2(new_n751), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT107), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n764), .A2(new_n758), .A3(new_n781), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n737), .A2(new_n630), .A3(new_n669), .A4(new_n647), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n737), .A2(new_n763), .A3(new_n647), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n708), .A2(new_n554), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n772), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT107), .B1(new_n835), .B2(new_n753), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n318), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n430), .B1(new_n662), .B2(new_n668), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n635), .A3(new_n644), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n631), .A2(new_n681), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n783), .A2(new_n680), .A3(new_n772), .A4(new_n791), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n648), .A2(new_n667), .A3(new_n686), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n574), .A2(new_n680), .A3(new_n791), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n797), .A3(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n795), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n837), .A2(KEYINPUT108), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n647), .A2(new_n648), .A3(new_n667), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n719), .A2(new_n721), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n849), .A2(new_n633), .A3(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n720), .A2(new_n729), .B1(new_n713), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n696), .A2(new_n852), .A3(new_n853), .A4(new_n784), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n574), .A2(new_n691), .A3(KEYINPUT95), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT95), .B1(new_n574), .B2(new_n691), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n784), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT109), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n784), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n852), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n855), .B1(new_n862), .B2(KEYINPUT52), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n835), .A2(new_n753), .A3(KEYINPUT107), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n846), .A2(new_n841), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n792), .A2(new_n787), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n793), .A2(new_n794), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT108), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n848), .A2(new_n863), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(KEYINPUT110), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n713), .A2(new_n851), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n724), .A2(new_n728), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n698), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n574), .A2(new_n680), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT52), .B1(new_n858), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n837), .A2(new_n854), .A3(new_n847), .A4(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(KEYINPUT111), .B(KEYINPUT53), .Z(new_n883));
  OAI21_X1  g697(.A(new_n875), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT110), .B1(new_n873), .B2(new_n874), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n881), .A2(new_n854), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n883), .B1(new_n870), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT112), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT112), .B(new_n883), .C1(new_n870), .C2(new_n887), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n846), .ZN(new_n895));
  INV_X1    g709(.A(new_n841), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n835), .A2(new_n753), .A3(KEYINPUT53), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n795), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n894), .B1(new_n863), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n886), .A2(KEYINPUT54), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n772), .A2(new_n778), .ZN(new_n902));
  INV_X1    g716(.A(new_n426), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n800), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n762), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(G952), .A3(new_n231), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT48), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n790), .A2(new_n761), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n787), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n713), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n630), .A3(new_n426), .A4(new_n910), .ZN(new_n915));
  OAI221_X1 g729(.A(new_n913), .B1(new_n909), .B2(new_n912), .C1(new_n662), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n821), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT114), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n734), .A2(new_n735), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n736), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(KEYINPUT114), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n808), .A3(new_n906), .ZN(new_n923));
  NOR4_X1   g737(.A1(new_n905), .A2(new_n317), .A3(new_n704), .A4(new_n761), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT50), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n680), .A3(new_n772), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n743), .A2(new_n470), .A3(new_n740), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n926), .C1(new_n915), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT115), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT51), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n923), .B(new_n929), .C1(new_n928), .C2(new_n931), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n790), .B(new_n905), .C1(new_n917), .C2(new_n920), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT51), .B1(new_n928), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n916), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n901), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(G952), .B2(G953), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n786), .A2(new_n646), .A3(new_n736), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n939), .A2(KEYINPUT105), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(KEYINPUT105), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n940), .A2(new_n941), .A3(new_n799), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(KEYINPUT106), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n919), .B(KEYINPUT49), .Z(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n713), .A3(new_n704), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n937), .A2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n863), .A2(new_n899), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT112), .B1(new_n882), .B2(new_n883), .ZN(new_n952));
  INV_X1    g766(.A(new_n891), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(G902), .ZN(new_n955));
  INV_X1    g769(.A(G210), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n296), .A2(new_n300), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(new_n298), .Z(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n957), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n957), .A2(new_n961), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n231), .A2(G952), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(G51));
  NOR2_X1   g779(.A1(new_n955), .A2(new_n812), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n954), .A2(KEYINPUT119), .A3(new_n894), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT119), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n969), .A2(new_n854), .A3(new_n899), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n890), .B2(new_n891), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n968), .B1(new_n971), .B2(new_n893), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT118), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n892), .A2(new_n973), .A3(new_n900), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(new_n892), .B2(new_n900), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n967), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n387), .B(KEYINPUT57), .Z(new_n978));
  AOI21_X1  g792(.A(new_n748), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT120), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n966), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n892), .A2(new_n900), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT118), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n893), .B1(new_n892), .B2(new_n951), .ZN(new_n985));
  AOI22_X1  g799(.A1(new_n984), .A2(new_n974), .B1(new_n985), .B2(KEYINPUT119), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n982), .B1(new_n986), .B2(new_n972), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT120), .B1(new_n987), .B2(new_n748), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n964), .B1(new_n981), .B2(new_n988), .ZN(G54));
  NAND4_X1  g803(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n990));
  INV_X1    g804(.A(new_n491), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n964), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n991), .B2(new_n990), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT121), .ZN(G60));
  AND2_X1   g808(.A1(new_n651), .A2(new_n656), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n658), .B(KEYINPUT59), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n901), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n995), .A2(new_n996), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n964), .B1(new_n977), .B2(new_n998), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n997), .A2(new_n999), .ZN(G63));
  XNOR2_X1  g814(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G217), .A2(G902), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n971), .A2(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1004), .A2(new_n678), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT61), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n1005), .A2(new_n1006), .A3(new_n964), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n615), .B1(new_n971), .B2(new_n1003), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1009), .A2(KEYINPUT123), .A3(new_n964), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT123), .ZN(new_n1014));
  INV_X1    g828(.A(new_n964), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1014), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1013), .A2(new_n1016), .A3(new_n1005), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n1017), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g832(.A(new_n429), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n231), .B1(new_n1019), .B2(G224), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n837), .A2(new_n896), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(new_n231), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n958), .B1(G898), .B2(new_n231), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT126), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT125), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1022), .B(new_n1025), .ZN(G69));
  XNOR2_X1  g840(.A(new_n564), .B(new_n480), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n819), .A2(new_n823), .ZN(new_n1028));
  INV_X1    g842(.A(new_n701), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n790), .B1(new_n662), .B2(new_n668), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1029), .A2(new_n574), .A3(new_n630), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n859), .A2(new_n730), .A3(new_n861), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n716), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1032), .B1(KEYINPUT62), .B2(new_n1034), .ZN(new_n1035));
  OR2_X1    g849(.A1(new_n1034), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1027), .B1(new_n1037), .B2(new_n231), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n817), .A2(new_n779), .A3(new_n787), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1039), .A2(new_n869), .A3(new_n797), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n1028), .A2(new_n1033), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n1041), .A2(G953), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1027), .B1(new_n685), .B2(new_n231), .ZN(new_n1043));
  NOR2_X1   g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(KEYINPUT127), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT127), .ZN(new_n1046));
  AOI21_X1  g860(.A(G953), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1047));
  OAI221_X1 g861(.A(new_n1046), .B1(new_n1042), .B2(new_n1043), .C1(new_n1047), .C2(new_n1027), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n231), .B1(G227), .B2(G900), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1045), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1049), .ZN(new_n1051));
  OAI211_X1 g865(.A(KEYINPUT127), .B(new_n1051), .C1(new_n1038), .C2(new_n1044), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1050), .A2(new_n1052), .ZN(G72));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  OAI21_X1  g869(.A(new_n1055), .B1(new_n1037), .B2(new_n1021), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n544), .A2(new_n545), .ZN(new_n1057));
  INV_X1    g871(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1056), .A2(new_n508), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1055), .B1(new_n1041), .B2(new_n1021), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n1058), .A2(new_n508), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n964), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n565), .A2(new_n567), .A3(new_n546), .ZN(new_n1064));
  AND2_X1   g878(.A1(new_n1064), .A2(new_n1055), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1063), .B1(new_n886), .B2(new_n1065), .ZN(G57));
endmodule


