//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT15), .Z(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT94), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n208), .B(KEYINPUT14), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT94), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n203), .A2(new_n207), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(KEYINPUT15), .B(new_n202), .C1(new_n212), .C2(new_n206), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n216), .B(KEYINPUT17), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n223), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n216), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT95), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(KEYINPUT18), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(new_n223), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n226), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n229), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n224), .A2(new_n226), .A3(new_n229), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G113gat), .B(G141gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G169gat), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT12), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n239), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n230), .A2(new_n235), .A3(new_n238), .A4(new_n247), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n246), .A2(KEYINPUT96), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT96), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n253), .B(G22gat), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G155gat), .A2(G162gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G155gat), .A2(G162gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G141gat), .B(G148gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(G155gat), .B2(G162gat), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G141gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G148gat), .ZN(new_n264));
  INV_X1    g063(.A(G148gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G141gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268));
  INV_X1    g067(.A(G155gat), .ZN(new_n269));
  INV_X1    g068(.A(G162gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT2), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT86), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279));
  INV_X1    g078(.A(G211gat), .ZN(new_n280));
  INV_X1    g079(.A(G218gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(G211gat), .B(G218gat), .Z(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT79), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT78), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n283), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n284), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT3), .B1(new_n291), .B2(new_n275), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n262), .A2(new_n272), .ZN(new_n293));
  OAI22_X1  g092(.A1(new_n277), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G228gat), .ZN(new_n295));
  INV_X1    g094(.A(G233gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n283), .A2(new_n284), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT85), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT29), .B1(new_n287), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n273), .B1(new_n300), .B2(KEYINPUT3), .ZN(new_n301));
  INV_X1    g100(.A(new_n291), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n276), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n294), .B(new_n297), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OAI22_X1  g105(.A1(new_n304), .A2(KEYINPUT84), .B1(new_n295), .B2(new_n296), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT31), .B(G50gat), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n306), .B2(new_n307), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n255), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n306), .A2(new_n307), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n308), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(new_n254), .A3(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT27), .B(G183gat), .Z(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT27), .B(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(KEYINPUT67), .B(G190gat), .Z(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT28), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(KEYINPUT69), .A2(KEYINPUT28), .ZN(new_n329));
  AOI211_X1 g128(.A(new_n328), .B(new_n329), .C1(new_n324), .C2(new_n320), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n332), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT71), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n325), .A2(new_n331), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT72), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  INV_X1    g143(.A(new_n324), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n319), .B2(new_n322), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n330), .B1(new_n346), .B2(KEYINPUT28), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n341), .A2(new_n338), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(KEYINPUT67), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n350), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n332), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n360), .A2(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT24), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT65), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT65), .ZN(new_n369));
  OAI22_X1  g168(.A1(new_n357), .A2(new_n369), .B1(G183gat), .B2(G190gat), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT66), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n366), .B2(KEYINPUT65), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n369), .B1(new_n356), .B2(new_n357), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n376), .A3(new_n363), .ZN(new_n377));
  XOR2_X1   g176(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n378));
  AOI221_X4 g177(.A(KEYINPUT68), .B1(new_n359), .B2(new_n363), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n363), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n343), .B(new_n349), .C1(new_n379), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G226gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n377), .A2(new_n378), .B1(new_n363), .B2(new_n359), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n275), .B1(new_n342), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n302), .B1(new_n389), .B2(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT80), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n386), .A2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n384), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n342), .A2(new_n388), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(new_n302), .C1(new_n385), .C2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n387), .A2(new_n397), .A3(new_n390), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT81), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G8gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(new_n205), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n392), .A2(new_n396), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n407));
  INV_X1    g206(.A(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n404), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G127gat), .B(G134gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415));
  INV_X1    g214(.A(G120gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(G113gat), .ZN(new_n417));
  INV_X1    g216(.A(G113gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G120gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n415), .B1(new_n420), .B2(KEYINPUT73), .ZN(new_n421));
  XNOR2_X1  g220(.A(G113gat), .B(G120gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n414), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT74), .B1(new_n418), .B2(G120gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT74), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(new_n416), .A3(G113gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n428), .A3(new_n419), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(new_n415), .A3(new_n413), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n293), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT4), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT1), .B1(new_n422), .B2(new_n423), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(KEYINPUT73), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n413), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n429), .A2(new_n415), .A3(new_n413), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n293), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n430), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n274), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(KEYINPUT5), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n440), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n445), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n438), .B1(new_n437), .B2(new_n293), .ZN(new_n450));
  AND4_X1   g249(.A1(new_n438), .A2(new_n425), .A3(new_n293), .A4(new_n430), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n449), .B(new_n443), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n273), .B1(new_n435), .B2(new_n436), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n431), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n456), .B2(new_n445), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n453), .B1(new_n452), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n448), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT0), .B(G57gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(G1gat), .B(G29gat), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n462), .B(new_n463), .Z(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n464), .B(new_n448), .C1(new_n458), .C2(new_n459), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n467), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n468), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n317), .B1(new_n412), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT77), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT36), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(KEYINPUT77), .A2(KEYINPUT36), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n388), .B(new_n380), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(new_n441), .A3(new_n343), .A4(new_n349), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n384), .A2(new_n437), .ZN(new_n480));
  INV_X1    g279(.A(G227gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n481), .A2(new_n296), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n483), .B1(KEYINPUT32), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT75), .B(G15gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(G71gat), .B(G99gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n489), .B2(KEYINPUT33), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n483), .A2(KEYINPUT76), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT76), .B1(new_n483), .B2(new_n492), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n482), .B1(new_n479), .B2(new_n480), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT34), .B(new_n482), .C1(new_n479), .C2(new_n480), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n495), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n493), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n505), .B2(new_n490), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n476), .B(new_n477), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n496), .A2(new_n502), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(new_n501), .A3(new_n490), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n474), .A4(new_n475), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n473), .A2(new_n507), .A3(KEYINPUT87), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n473), .A2(new_n507), .A3(new_n510), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n460), .A2(new_n515), .A3(new_n465), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n460), .B2(new_n465), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n471), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n468), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n403), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n522));
  NOR2_X1   g321(.A1(new_n402), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n407), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n394), .B1(new_n385), .B2(new_n395), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n291), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n384), .A2(new_n386), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n389), .A2(new_n385), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n302), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(KEYINPUT37), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n524), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n392), .A2(new_n396), .A3(KEYINPUT37), .A4(new_n398), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n402), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n522), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n317), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n452), .A2(new_n457), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT83), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n452), .A2(new_n453), .A3(new_n457), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n447), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT90), .B1(new_n543), .B2(new_n464), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n516), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n274), .A2(new_n441), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n442), .A2(new_n546), .B1(new_n432), .B2(new_n439), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT88), .B1(new_n547), .B2(new_n444), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n440), .A2(new_n443), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(new_n445), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT39), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT89), .B1(new_n456), .B2(new_n445), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n456), .A2(KEYINPUT89), .A3(new_n445), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n553), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n548), .A2(new_n551), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n464), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT40), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT40), .A4(new_n464), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n412), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT92), .B1(new_n539), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n470), .B1(new_n544), .B2(new_n516), .ZN(new_n567));
  INV_X1    g366(.A(new_n403), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n567), .A2(new_n468), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n387), .A2(new_n397), .A3(new_n390), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n397), .B1(new_n387), .B2(new_n390), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n342), .A2(new_n388), .A3(new_n385), .ZN(new_n572));
  AOI211_X1 g371(.A(new_n291), .B(new_n572), .C1(new_n384), .C2(new_n393), .ZN(new_n573));
  NOR3_X1   g372(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n532), .B1(new_n574), .B2(KEYINPUT37), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n523), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n569), .B(new_n576), .C1(new_n536), .C2(new_n537), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n312), .A2(new_n316), .ZN(new_n578));
  AND4_X1   g377(.A1(KEYINPUT92), .A2(new_n577), .A3(new_n578), .A4(new_n565), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n511), .B(new_n514), .C1(new_n566), .C2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n468), .B1(new_n545), .B2(new_n471), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(new_n409), .A3(new_n406), .A4(new_n411), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n578), .A2(new_n508), .A3(new_n509), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n412), .A2(new_n472), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n503), .A2(new_n506), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n587), .A2(KEYINPUT35), .A3(new_n588), .A4(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n252), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  INV_X1    g392(.A(G64gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n593), .B1(new_n594), .B2(G57gat), .ZN(new_n595));
  INV_X1    g394(.A(G57gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT97), .A3(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  OR2_X1    g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(KEYINPUT98), .A3(new_n599), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G57gat), .B(G64gat), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n603), .B(new_n604), .C1(new_n609), .C2(new_n605), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n608), .A2(KEYINPUT99), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT99), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n225), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G183gat), .ZN(new_n616));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT102), .B(G211gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n618), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT101), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n631));
  NAND2_X1  g430(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n631), .A2(G85gat), .A3(G92gat), .A4(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(G85gat), .ZN(new_n634));
  INV_X1    g433(.A(G92gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n637), .A2(new_n638), .B1(new_n639), .B2(KEYINPUT8), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n633), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G99gat), .B(G106gat), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n633), .A2(new_n640), .A3(new_n636), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n642), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT104), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n217), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g450(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n216), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n352), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n352), .B1(new_n651), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n281), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(G218gat), .A3(new_n655), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(KEYINPUT105), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT105), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OR3_X1    g465(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  INV_X1    g470(.A(new_n648), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n608), .A2(new_n610), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT99), .ZN(new_n674));
  INV_X1    g473(.A(new_n612), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n648), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n653), .A2(KEYINPUT10), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n613), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n614), .A2(KEYINPUT106), .A3(KEYINPUT10), .A4(new_n653), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n678), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(G230gat), .A2(G233gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n676), .A2(new_n677), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G176gat), .B(G204gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT107), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G120gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(new_n265), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n687), .B(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n630), .A2(new_n670), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n592), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n472), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g495(.A1(new_n694), .A2(new_n412), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n699), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n222), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n701), .B1(new_n699), .B2(KEYINPUT42), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT108), .B1(new_n699), .B2(KEYINPUT42), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(G1325gat));
  AND2_X1   g503(.A1(new_n694), .A2(new_n588), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(G15gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n507), .A2(new_n510), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n694), .A2(G15gat), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT110), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n317), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n630), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n692), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n592), .A2(new_n670), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n204), .A3(new_n472), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n580), .A2(new_n591), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n669), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT92), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n576), .A2(new_n582), .A3(new_n403), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n536), .A2(new_n537), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n578), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n565), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n577), .A2(KEYINPUT92), .A3(new_n565), .A4(new_n578), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n512), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n590), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n721), .B1(new_n733), .B2(new_n669), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n246), .A2(new_n248), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n723), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT111), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n723), .A2(new_n734), .A3(new_n737), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n472), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n719), .B1(new_n743), .B2(new_n204), .ZN(G1328gat));
  NAND3_X1  g543(.A1(new_n717), .A2(new_n205), .A3(new_n412), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT46), .Z(new_n746));
  INV_X1    g545(.A(new_n412), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n739), .B2(new_n741), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n205), .B2(new_n748), .ZN(G1329gat));
  INV_X1    g548(.A(new_n708), .ZN(new_n750));
  OAI21_X1  g549(.A(G43gat), .B1(new_n738), .B2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(G43gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n717), .A2(new_n752), .A3(new_n588), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n753), .A3(KEYINPUT47), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n750), .B1(new_n739), .B2(new_n741), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(new_n752), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT47), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n754), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g562(.A(KEYINPUT113), .B(new_n754), .C1(new_n759), .C2(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1330gat));
  OAI21_X1  g564(.A(G50gat), .B1(new_n738), .B2(new_n578), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n578), .A2(G50gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n717), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(KEYINPUT48), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n742), .A2(new_n317), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n770), .A2(G50gat), .B1(new_n717), .B2(new_n767), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g571(.A1(new_n733), .A2(new_n735), .ZN(new_n773));
  INV_X1    g572(.A(new_n692), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n630), .A2(new_n670), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n472), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g578(.A1(new_n776), .A2(new_n747), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  AND2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(new_n780), .B2(new_n781), .ZN(G1333gat));
  INV_X1    g583(.A(G71gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n777), .A2(new_n785), .A3(new_n588), .ZN(new_n786));
  OAI21_X1  g585(.A(G71gat), .B1(new_n776), .B2(new_n750), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g588(.A1(new_n777), .A2(new_n317), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(G78gat), .ZN(G1335gat));
  INV_X1    g590(.A(new_n733), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n715), .A2(new_n735), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n670), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n774), .ZN(new_n796));
  AOI21_X1  g595(.A(G85gat), .B1(new_n796), .B2(new_n472), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n723), .A2(new_n734), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n692), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n800), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n634), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n797), .B1(new_n807), .B2(new_n472), .ZN(G1336gat));
  NOR2_X1   g607(.A1(new_n747), .A2(G92gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n796), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  OAI21_X1  g610(.A(G92gat), .B1(new_n801), .B2(new_n747), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n635), .B1(new_n805), .B2(new_n412), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n796), .B2(new_n809), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n815), .B2(new_n811), .ZN(G1337gat));
  OAI21_X1  g615(.A(G99gat), .B1(new_n806), .B2(new_n750), .ZN(new_n817));
  INV_X1    g616(.A(G99gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n796), .A2(new_n818), .A3(new_n588), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1338gat));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(G106gat), .C1(new_n806), .C2(new_n578), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n578), .A2(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n796), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n578), .B1(new_n802), .B2(new_n804), .ZN(new_n825));
  INV_X1    g624(.A(G106gat), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT116), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n822), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n798), .A2(new_n800), .A3(new_n317), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n832), .B2(G106gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n796), .A2(KEYINPUT117), .A3(new_n823), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n829), .A2(new_n835), .ZN(G1339gat));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  INV_X1    g637(.A(new_n684), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n678), .A2(new_n682), .A3(new_n681), .A4(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n840), .B2(KEYINPUT118), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n685), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n691), .B1(new_n685), .B2(KEYINPUT54), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT119), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n687), .A2(new_n691), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n840), .ZN(new_n849));
  INV_X1    g648(.A(new_n841), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(KEYINPUT55), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n838), .C1(new_n844), .C2(new_n845), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n847), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n847), .A2(new_n852), .A3(KEYINPUT120), .A4(new_n854), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n227), .A2(new_n229), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n233), .A2(new_n234), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n244), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n248), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n670), .A2(new_n857), .A3(new_n858), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n857), .A2(new_n735), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n692), .A2(new_n862), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n837), .B(new_n863), .C1(new_n866), .C2(new_n670), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n670), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  INV_X1    g667(.A(new_n863), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT121), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n630), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n735), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n693), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n585), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n747), .A2(new_n472), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n252), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n418), .A3(new_n735), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1340gat));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n692), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g681(.A1(new_n876), .A2(new_n715), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g683(.A1(new_n876), .A2(new_n670), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(G134gat), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT56), .B1(new_n885), .B2(G134gat), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G1343gat));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n578), .B1(new_n871), .B2(new_n873), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n750), .A2(new_n875), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n891), .A2(new_n263), .A3(new_n251), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n871), .A2(new_n873), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n317), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT57), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n251), .A2(new_n852), .A3(new_n846), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n865), .B(KEYINPUT122), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n669), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n863), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n630), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n578), .B1(new_n902), .B2(new_n873), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n893), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n897), .A2(new_n252), .A3(new_n905), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n890), .B(new_n894), .C1(new_n906), .C2(new_n263), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n894), .A2(new_n908), .ZN(new_n909));
  AOI211_X1 g708(.A(G141gat), .B(new_n578), .C1(new_n871), .C2(new_n873), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n251), .A4(new_n893), .ZN(new_n911));
  AOI211_X1 g710(.A(new_n872), .B(new_n905), .C1(new_n891), .C2(new_n904), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n909), .B(new_n911), .C1(new_n912), .C2(new_n263), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT58), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n913), .B2(KEYINPUT58), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G1344gat));
  NAND4_X1  g716(.A1(new_n891), .A2(new_n265), .A3(new_n692), .A4(new_n893), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n670), .A2(new_n862), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n900), .B1(new_n855), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n630), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n693), .A2(new_n252), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT57), .B(new_n578), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n692), .A3(new_n893), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n265), .B1(new_n926), .B2(KEYINPUT125), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n925), .A2(new_n928), .A3(new_n692), .A4(new_n893), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n897), .A2(new_n905), .ZN(new_n931));
  AOI211_X1 g730(.A(KEYINPUT59), .B(new_n265), .C1(new_n931), .C2(new_n692), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n918), .B1(new_n930), .B2(new_n932), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n931), .A2(G155gat), .A3(new_n715), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n891), .A2(new_n893), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n269), .B1(new_n935), .B2(new_n630), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n934), .A2(new_n936), .ZN(G1346gat));
  NAND3_X1  g736(.A1(new_n931), .A2(G162gat), .A3(new_n670), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n270), .B1(new_n935), .B2(new_n669), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n938), .A2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n747), .A2(new_n472), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n874), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n943), .A2(G169gat), .A3(new_n872), .ZN(new_n944));
  OAI21_X1  g743(.A(G169gat), .B1(new_n943), .B2(new_n252), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1348gat));
  NAND2_X1  g745(.A1(new_n942), .A2(new_n692), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n323), .A3(new_n715), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n943), .A2(new_n630), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n351), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n943), .B2(new_n669), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n943), .A2(new_n669), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n955), .B1(new_n956), .B2(new_n324), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n953), .B2(new_n957), .ZN(G1351gat));
  INV_X1    g757(.A(new_n924), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n750), .A2(new_n941), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n959), .B(new_n961), .C1(new_n891), .C2(new_n904), .ZN(new_n962));
  OAI21_X1  g761(.A(G197gat), .B1(new_n962), .B2(new_n252), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n896), .A2(new_n960), .ZN(new_n964));
  INV_X1    g763(.A(G197gat), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n965), .A3(new_n735), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1352gat));
  NOR4_X1   g766(.A1(new_n896), .A2(G204gat), .A3(new_n774), .A4(new_n960), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n925), .A2(new_n692), .A3(new_n961), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(G204gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n964), .A2(new_n280), .A3(new_n715), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n925), .A2(KEYINPUT126), .A3(new_n715), .A4(new_n961), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n962), .B2(new_n630), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n974), .A2(G211gat), .A3(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n973), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  XOR2_X1   g780(.A(new_n962), .B(KEYINPUT127), .Z(new_n982));
  OAI21_X1  g781(.A(G218gat), .B1(new_n982), .B2(new_n669), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n964), .A2(new_n281), .A3(new_n670), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n983), .A2(new_n984), .ZN(G1355gat));
endmodule


