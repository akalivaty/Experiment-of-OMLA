//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n209), .A2(G13), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT0), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n203), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n222), .A2(new_n223), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n223), .B2(new_n222), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n220), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  NAND2_X1  g0042(.A1(new_n211), .A2(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n250), .A2(new_n252), .A3(G223), .A4(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G87), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n250), .A2(new_n252), .A3(G1698), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n212), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G190), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n258), .A2(new_n263), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(G232), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n259), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT77), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT77), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n259), .A2(new_n269), .A3(new_n266), .A4(new_n260), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n259), .A2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT16), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT75), .B1(new_n201), .B2(new_n202), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT75), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G58), .A3(G68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n278), .A3(new_n203), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G20), .ZN(new_n280));
  INV_X1    g0080(.A(G159), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT7), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT3), .B(G33), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n285), .B1(new_n286), .B2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n250), .A2(new_n252), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT7), .A3(new_n227), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n202), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n275), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n286), .A2(new_n285), .A3(G20), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT7), .B1(new_n288), .B2(new_n227), .ZN(new_n293));
  OAI21_X1  g0093(.A(G68), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n279), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(KEYINPUT16), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n226), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n291), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(KEYINPUT67), .B1(new_n201), .B2(KEYINPUT8), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT8), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(G58), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(G58), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G1), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n306), .B2(G20), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(G13), .A3(G20), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n299), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT17), .B1(new_n274), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n297), .A2(new_n226), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n294), .A2(new_n295), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n314), .B1(new_n315), .B2(new_n275), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n310), .B1(new_n316), .B2(new_n296), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT17), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n259), .A2(new_n323), .A3(new_n266), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT76), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT76), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n259), .A2(new_n326), .A3(new_n266), .A4(new_n323), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n271), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n322), .B1(new_n317), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n325), .A2(new_n327), .A3(new_n329), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT18), .A3(new_n312), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n321), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT78), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n307), .A2(G77), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G77), .B2(new_n309), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n303), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n342), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n249), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(KEYINPUT15), .B(G87), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n339), .B1(new_n347), .B2(new_n298), .ZN(new_n348));
  OAI211_X1 g0148(.A(G1), .B(G13), .C1(new_n249), .C2(new_n261), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT65), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n256), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n286), .A2(KEYINPUT65), .A3(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(G238), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n250), .A2(new_n252), .A3(G232), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n253), .B1(G107), .B2(new_n288), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n349), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n263), .A2(G274), .ZN(new_n357));
  INV_X1    g0157(.A(new_n265), .ZN(new_n358));
  INV_X1    g0158(.A(G244), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n348), .B1(new_n361), .B2(new_n272), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT69), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n348), .B(KEYINPUT69), .C1(new_n361), .C2(new_n272), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(G190), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n348), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n361), .A2(new_n323), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n328), .B1(new_n356), .B2(new_n360), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n337), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT73), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n250), .A2(new_n252), .A3(G232), .A4(G1698), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n250), .A2(new_n252), .A3(G226), .A4(new_n253), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n258), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n306), .B1(G41), .B2(G45), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n349), .A2(G238), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT70), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n380), .A2(new_n381), .A3(new_n357), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n380), .B2(new_n357), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n357), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT70), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n381), .A3(new_n357), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n378), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n391), .A3(G179), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n328), .B1(new_n385), .B2(new_n391), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT14), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI211_X1 g0195(.A(KEYINPUT14), .B(new_n328), .C1(new_n385), .C2(new_n391), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n373), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n384), .A2(KEYINPUT13), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n390), .B1(new_n389), .B2(new_n378), .ZN(new_n399));
  OAI21_X1  g0199(.A(G169), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n393), .A2(new_n394), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n401), .A2(KEYINPUT73), .A3(new_n402), .A4(new_n392), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n309), .A2(G68), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT12), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT71), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n407), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n307), .A2(G68), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n344), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n211), .B2(new_n283), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT11), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n413), .A2(new_n414), .A3(new_n298), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n414), .B1(new_n413), .B2(new_n298), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n410), .B(new_n411), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n417), .B(KEYINPUT74), .Z(new_n418));
  NAND3_X1  g0218(.A1(new_n397), .A2(new_n403), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n417), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n385), .A2(new_n391), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(new_n260), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(G200), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT72), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n398), .A2(new_n399), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n417), .B1(new_n426), .B2(G190), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT72), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(new_n428), .A3(new_n423), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n264), .B1(new_n265), .B2(G226), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n205), .B1(new_n250), .B2(new_n252), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n288), .A2(G1698), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(G222), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n351), .A2(new_n352), .A3(G223), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT66), .B(new_n432), .C1(new_n437), .C2(new_n349), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT66), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n349), .B1(new_n435), .B2(new_n436), .ZN(new_n440));
  INV_X1    g0240(.A(new_n432), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n438), .A2(G200), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n211), .B1(new_n306), .B2(G20), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT68), .ZN(new_n445));
  INV_X1    g0245(.A(new_n309), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n298), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n445), .A2(new_n447), .B1(new_n211), .B2(new_n446), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n345), .B1(new_n302), .B2(new_n304), .ZN(new_n449));
  INV_X1    g0249(.A(G150), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n204), .A2(new_n227), .B1(new_n283), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n298), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n448), .A2(new_n452), .A3(KEYINPUT9), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT9), .B1(new_n448), .B2(new_n452), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n443), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n260), .B1(new_n438), .B2(new_n442), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT10), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n438), .A2(new_n442), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G190), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT10), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n443), .A4(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n448), .A2(new_n452), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n459), .B2(new_n323), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G169), .B2(new_n459), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n463), .B(new_n466), .C1(new_n335), .C2(new_n336), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n372), .A2(new_n431), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT19), .ZN(new_n470));
  INV_X1    g0270(.A(G97), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G97), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n470), .B1(new_n475), .B2(new_n345), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n227), .B1(new_n376), .B2(new_n470), .ZN(new_n477));
  XNOR2_X1  g0277(.A(KEYINPUT79), .B(G97), .ZN(new_n478));
  INV_X1    g0278(.A(G107), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n213), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n286), .A2(new_n227), .A3(G68), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n476), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n298), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n346), .B(KEYINPUT83), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n306), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n309), .A2(new_n486), .A3(new_n226), .A4(new_n297), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n346), .A2(new_n446), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n484), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(G1698), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n250), .A2(new_n252), .A3(G238), .A4(new_n253), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G116), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n258), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n262), .A2(G1), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n214), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n498), .A2(new_n349), .B1(G274), .B2(new_n497), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n328), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n323), .A3(new_n499), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n491), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n490), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n487), .A2(new_n213), .ZN(new_n505));
  AOI211_X1 g0305(.A(new_n504), .B(new_n505), .C1(new_n483), .C2(new_n298), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(G190), .A3(new_n499), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n500), .A2(G200), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(new_n253), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  INV_X1    g0311(.A(G257), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n510), .B(new_n511), .C1(new_n256), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n258), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n261), .A3(KEYINPUT5), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(KEYINPUT81), .B2(G41), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n518), .A3(new_n497), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n519), .A2(new_n349), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G264), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n516), .A2(new_n518), .A3(new_n497), .A4(G274), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n514), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n514), .A2(new_n521), .A3(G190), .A4(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n446), .A2(KEYINPUT25), .A3(new_n479), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n309), .B2(G107), .ZN(new_n529));
  AOI22_X1  g0329(.A1(G107), .A2(new_n488), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n479), .A2(KEYINPUT23), .A3(G20), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT23), .B1(new_n479), .B2(G20), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(G20), .B2(new_n494), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n250), .A2(new_n252), .A3(new_n227), .A4(G87), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT22), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n286), .A2(new_n536), .A3(new_n227), .A4(G87), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n298), .B1(new_n538), .B2(KEYINPUT24), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n530), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n503), .B(new_n509), .C1(new_n526), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n523), .A2(new_n328), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n514), .A2(new_n521), .A3(new_n323), .A4(new_n522), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n286), .A2(G264), .A3(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n288), .A2(G303), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n286), .A2(new_n253), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n550), .C2(new_n512), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n258), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n519), .A2(G270), .A3(new_n349), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n522), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G169), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n488), .A2(G116), .ZN(new_n558));
  INV_X1    g0358(.A(G116), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n446), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n227), .B(new_n562), .C1(new_n475), .C2(G33), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n298), .B1(new_n227), .B2(G116), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT20), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n227), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n478), .B2(new_n249), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n567), .B1(new_n569), .B2(new_n564), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n561), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n547), .B1(new_n557), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n554), .B1(new_n258), .B2(new_n551), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n574), .B(new_n571), .C1(new_n272), .C2(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n566), .A2(new_n570), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n576), .A2(new_n558), .A3(new_n560), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n577), .A2(KEYINPUT21), .A3(G169), .A4(new_n556), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(G179), .A3(new_n573), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n572), .A2(new_n575), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n250), .A2(new_n252), .A3(G250), .A4(G1698), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n250), .A2(new_n252), .A3(G244), .A4(new_n253), .ZN(new_n582));
  NOR2_X1   g0382(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n562), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  XNOR2_X1  g0384(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n258), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n520), .A2(G257), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n522), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n591), .A2(G107), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n472), .A3(new_n474), .ZN(new_n593));
  AND2_X1   g0393(.A1(G97), .A2(G107), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G97), .A2(G107), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G20), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n282), .A2(G77), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n479), .B1(new_n287), .B2(new_n289), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n298), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n309), .A2(G97), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n603), .B1(new_n488), .B2(G97), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n587), .A2(G190), .A3(new_n522), .A4(new_n588), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n590), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n589), .A2(new_n328), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n604), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n587), .A2(new_n323), .A3(new_n522), .A4(new_n588), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n606), .A2(new_n610), .A3(KEYINPUT82), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT82), .B1(new_n606), .B2(new_n610), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n546), .B(new_n580), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n469), .A2(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n371), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n430), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n419), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n617), .A2(new_n321), .ZN(new_n618));
  INV_X1    g0418(.A(new_n334), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n463), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT85), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n328), .A2(new_n589), .B1(new_n602), .B2(new_n604), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n622), .A2(new_n609), .A3(new_n503), .A4(new_n509), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n509), .A2(new_n503), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n610), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(KEYINPUT84), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n629), .B(new_n624), .C1(new_n626), .C2(new_n610), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n503), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n621), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n623), .A2(new_n624), .ZN(new_n634));
  INV_X1    g0434(.A(new_n630), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n629), .B1(new_n623), .B2(new_n624), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(KEYINPUT85), .A3(new_n503), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n541), .A2(new_n543), .A3(new_n544), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n606), .A2(new_n610), .ZN(new_n642));
  INV_X1    g0442(.A(new_n542), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n633), .A2(new_n638), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n468), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n620), .A2(new_n466), .A3(new_n646), .ZN(G369));
  AND2_X1   g0447(.A1(new_n227), .A2(G13), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(new_n306), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(KEYINPUT27), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(G213), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n571), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n578), .A2(new_n579), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n572), .A3(new_n575), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n658), .B2(KEYINPUT86), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT86), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n580), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n657), .A2(new_n572), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n656), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n526), .A2(new_n541), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n541), .A2(new_n654), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n545), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n640), .A2(new_n654), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(G330), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n639), .A2(new_n654), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n221), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n478), .A2(G116), .A3(new_n480), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n224), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(new_n644), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n628), .A2(new_n630), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n632), .B1(new_n683), .B2(new_n634), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(KEYINPUT85), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n654), .B1(new_n685), .B2(new_n633), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n556), .A2(new_n323), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n587), .A2(new_n588), .ZN(new_n691));
  AND4_X1   g0491(.A1(new_n496), .A2(new_n514), .A3(new_n521), .A4(new_n499), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(G179), .B1(new_n496), .B2(new_n499), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n589), .A2(new_n556), .A3(new_n523), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n691), .A4(new_n692), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n689), .B1(new_n699), .B2(new_n654), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n613), .B2(new_n654), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(new_n689), .A3(new_n654), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G330), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n634), .A2(new_n627), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n644), .A2(new_n503), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n655), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n688), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n681), .B1(new_n709), .B2(G1), .ZN(G364));
  AOI21_X1  g0510(.A(new_n306), .B1(new_n648), .B2(G45), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n676), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n659), .A2(new_n661), .B1(new_n663), .B2(new_n656), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n716), .B2(new_n715), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n226), .B1(G20), .B2(new_n328), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n272), .A2(G179), .ZN(new_n721));
  NAND2_X1  g0521(.A1(G20), .A2(G190), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G303), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n288), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n722), .A2(new_n323), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G322), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n323), .A2(new_n272), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n726), .B(new_n730), .C1(G326), .C2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n227), .A2(G190), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n323), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(G311), .A2(new_n741), .B1(new_n744), .B2(G329), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n734), .A2(new_n738), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n735), .A2(new_n721), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT87), .ZN(new_n749));
  INV_X1    g0549(.A(G294), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n227), .B1(new_n742), .B2(G190), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT88), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT88), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n746), .B1(new_n747), .B2(new_n749), .C1(new_n750), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n744), .A2(G159), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n286), .B1(new_n211), .B2(new_n732), .C1(new_n756), .C2(KEYINPUT32), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(KEYINPUT32), .B2(new_n756), .ZN(new_n758));
  INV_X1    g0558(.A(new_n754), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G97), .ZN(new_n760));
  INV_X1    g0560(.A(new_n749), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n724), .A2(new_n213), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n731), .A2(new_n735), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n764), .A2(new_n202), .B1(new_n740), .B2(new_n205), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n763), .B(new_n765), .C1(G58), .C2(new_n727), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n758), .A2(new_n760), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n720), .B1(new_n755), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n719), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n286), .A2(G355), .A3(new_n221), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n247), .A2(new_n262), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n675), .A2(new_n286), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(G45), .B2(new_n224), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n773), .B1(G116), .B2(new_n221), .C1(new_n774), .C2(new_n776), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n714), .B(new_n768), .C1(new_n772), .C2(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT89), .Z(new_n779));
  NAND2_X1  g0579(.A1(new_n715), .A2(new_n771), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n718), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  NAND2_X1  g0582(.A1(new_n368), .A2(new_n654), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n615), .B1(new_n367), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n371), .A2(new_n654), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT94), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT94), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n362), .A2(new_n363), .B1(G190), .B2(new_n361), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(new_n365), .B1(new_n368), .B2(new_n654), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n787), .B(new_n788), .C1(new_n790), .C2(new_n615), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n786), .A2(KEYINPUT95), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT95), .B1(new_n786), .B2(new_n791), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n645), .A2(new_n655), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT96), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT96), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n786), .A2(new_n791), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n645), .A2(new_n655), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n797), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n713), .B1(new_n802), .B2(new_n703), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n703), .B2(new_n802), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n719), .A2(new_n769), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n714), .B1(new_n205), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n733), .A2(G303), .B1(new_n741), .B2(G116), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n736), .A2(KEYINPUT90), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT90), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n764), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n807), .B1(new_n812), .B2(new_n747), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT91), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n761), .A2(G87), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n288), .B1(new_n724), .B2(new_n479), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT92), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n744), .A2(G311), .B1(G294), .B2(new_n727), .ZN(new_n818));
  AND4_X1   g0618(.A1(new_n760), .A2(new_n815), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n286), .B1(new_n743), .B2(new_n820), .C1(new_n211), .C2(new_n724), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n749), .A2(new_n202), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(G58), .C2(new_n759), .ZN(new_n823));
  XNOR2_X1  g0623(.A(KEYINPUT93), .B(G143), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n736), .A2(G150), .B1(new_n727), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n826), .B2(new_n732), .C1(new_n281), .C2(new_n740), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT34), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n814), .A2(new_n819), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n806), .B1(new_n720), .B2(new_n829), .C1(new_n800), .C2(new_n770), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n804), .A2(new_n830), .ZN(G384));
  OAI211_X1 g0631(.A(G116), .B(new_n228), .C1(new_n597), .C2(KEYINPUT35), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(KEYINPUT35), .B2(new_n597), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT36), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n225), .A2(G77), .A3(new_n278), .A4(new_n276), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n306), .B(G13), .C1(new_n835), .C2(new_n243), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n317), .A2(new_n652), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n335), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n274), .A2(new_n312), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n330), .A2(new_n652), .B1(new_n299), .B2(new_n311), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n652), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n312), .B1(new_n332), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n317), .A2(new_n319), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(KEYINPUT37), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n839), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  INV_X1    g0650(.A(new_n838), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n321), .B2(new_n334), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n843), .A2(new_n847), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n419), .A2(new_n654), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n856), .A2(new_n857), .B1(new_n619), .B2(new_n652), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n418), .A2(new_n654), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n419), .B2(new_n430), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n419), .A2(new_n430), .A3(new_n859), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n801), .B2(new_n788), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n855), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n469), .B1(new_n688), .B2(new_n707), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n620), .A2(new_n466), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n867), .B(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n839), .B2(new_n848), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n852), .A2(new_n853), .A3(new_n850), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n419), .A2(new_n430), .A3(new_n859), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n873), .A2(new_n874), .B1(new_n875), .B2(new_n860), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n701), .A2(new_n702), .A3(new_n786), .A4(new_n791), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND4_X1   g0678(.A1(new_n701), .A2(new_n702), .A3(new_n786), .A4(new_n791), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n879), .A2(new_n863), .A3(KEYINPUT40), .A4(new_n855), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n468), .A2(new_n701), .A3(new_n702), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n878), .A2(G330), .A3(new_n880), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n469), .A2(new_n703), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n881), .A2(new_n882), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n871), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n306), .B2(new_n648), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n871), .A2(new_n886), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n837), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT97), .ZN(G367));
  INV_X1    g0691(.A(new_n775), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n772), .B1(new_n221), .B2(new_n346), .C1(new_n238), .C2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(KEYINPUT103), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n894), .A2(new_n895), .A3(new_n714), .ZN(new_n896));
  INV_X1    g0696(.A(new_n771), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n655), .A2(new_n506), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n632), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n626), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n759), .A2(G68), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n450), .B2(new_n728), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT104), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n286), .B1(new_n743), .B2(new_n826), .ZN(new_n904));
  INV_X1    g0704(.A(new_n724), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n733), .A2(new_n824), .B1(new_n905), .B2(G58), .ZN(new_n906));
  OAI221_X1 g0706(.A(new_n906), .B1(new_n211), .B2(new_n740), .C1(new_n205), .C2(new_n748), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n904), .B(new_n907), .C1(G159), .C2(new_n811), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT105), .Z(new_n910));
  AOI21_X1  g0710(.A(new_n286), .B1(new_n733), .B2(G311), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n905), .A2(KEYINPUT46), .A3(G116), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT46), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n724), .B2(new_n559), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n744), .A2(G317), .B1(G303), .B2(new_n727), .ZN(new_n916));
  INV_X1    g0716(.A(new_n748), .ZN(new_n917));
  AOI22_X1  g0717(.A1(G283), .A2(new_n741), .B1(new_n917), .B2(new_n478), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n916), .B(new_n918), .C1(new_n812), .C2(new_n750), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n915), .B(new_n919), .C1(G107), .C2(new_n759), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n910), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT47), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n720), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n896), .B1(new_n897), .B2(new_n900), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n900), .A2(KEYINPUT98), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n900), .A2(KEYINPUT98), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n928), .A2(new_n929), .A3(KEYINPUT43), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(KEYINPUT43), .B2(new_n900), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n608), .A2(new_n654), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n642), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n622), .A2(new_n609), .A3(new_n654), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT99), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n610), .B1(new_n936), .B2(new_n640), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n655), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT42), .ZN(new_n939));
  AND4_X1   g0739(.A1(new_n642), .A2(new_n670), .A3(new_n641), .A4(new_n672), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n939), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n941), .A2(KEYINPUT100), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(KEYINPUT100), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n938), .B1(new_n939), .B2(new_n940), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n930), .B(new_n931), .S(new_n944), .Z(new_n945));
  INV_X1    g0745(.A(new_n671), .ZN(new_n946));
  INV_X1    g0746(.A(new_n936), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n945), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n670), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n663), .A2(new_n655), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT102), .B1(new_n670), .B2(new_n672), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n955), .A2(new_n715), .A3(new_n716), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n665), .B2(G330), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n955), .B1(new_n715), .B2(new_n716), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n665), .A2(G330), .A3(new_n954), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n958), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n708), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n673), .B2(new_n935), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n951), .A2(new_n668), .B1(new_n640), .B2(new_n654), .ZN(new_n966));
  INV_X1    g0766(.A(new_n935), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT45), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n671), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(KEYINPUT101), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n969), .A2(new_n973), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n946), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT101), .B1(new_n977), .B2(new_n974), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n963), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n709), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n676), .B(KEYINPUT41), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n712), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n927), .B1(new_n949), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT106), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(G387));
  NAND2_X1  g0785(.A1(new_n962), .A2(new_n708), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n958), .A2(new_n961), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n987), .A2(new_n703), .A3(new_n707), .A4(new_n688), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(new_n988), .A3(new_n676), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n775), .B1(new_n235), .B2(new_n262), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n286), .A2(new_n221), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n678), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n341), .A2(G50), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g0794(.A(G45), .B1(G68), .B2(G77), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n678), .A3(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n992), .A2(new_n996), .B1(new_n479), .B2(new_n675), .ZN(new_n997));
  INV_X1    g0797(.A(new_n772), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n713), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n727), .A2(G317), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n740), .B2(new_n725), .C1(new_n729), .C2(new_n732), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n811), .B2(G311), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT48), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n759), .A2(G283), .B1(G294), .B2(new_n905), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(KEYINPUT48), .B2(new_n1002), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT49), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n748), .A2(new_n559), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n286), .B(new_n1011), .C1(G326), .C2(new_n744), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n761), .A2(G97), .B1(new_n305), .B2(new_n736), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n728), .A2(new_n211), .B1(new_n740), .B2(new_n202), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n286), .B1(new_n743), .B2(new_n450), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n732), .A2(new_n281), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n724), .A2(new_n205), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n485), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1014), .B(new_n1019), .C1(new_n1020), .C2(new_n754), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n720), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n999), .B(new_n1022), .C1(new_n950), .C2(new_n771), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n712), .B2(new_n987), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n989), .A2(new_n1024), .ZN(G393));
  NOR2_X1   g0825(.A1(new_n242), .A2(new_n892), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n998), .B1(new_n675), .B2(new_n478), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n714), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n288), .B1(new_n743), .B2(new_n729), .C1(new_n747), .C2(new_n724), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n761), .B2(G107), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT109), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n812), .A2(new_n725), .B1(new_n750), .B2(new_n740), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G116), .B2(new_n759), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n733), .A2(G317), .B1(G311), .B2(new_n727), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT52), .Z(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT110), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n811), .A2(G50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n288), .B1(new_n342), .B2(new_n741), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G68), .A2(new_n905), .B1(new_n744), .B2(new_n824), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n815), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n728), .A2(new_n281), .B1(new_n732), .B2(new_n450), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n759), .A2(G77), .ZN(new_n1046));
  AND4_X1   g0846(.A1(new_n1039), .A2(new_n1042), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1038), .A2(new_n1047), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1048), .A2(KEYINPUT111), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n719), .B1(new_n1048), .B2(KEYINPUT111), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1029), .B1(new_n947), .B2(new_n897), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n976), .B(new_n946), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n711), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n978), .A2(new_n975), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n677), .B1(new_n1054), .B2(new_n963), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT113), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT112), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n988), .A2(new_n1057), .A3(new_n1052), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n977), .A2(new_n974), .ZN(new_n1059));
  OAI21_X1  g0859(.A(KEYINPUT112), .B1(new_n963), .B2(new_n1059), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1060), .A2(new_n979), .A3(new_n676), .A4(new_n1058), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT113), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1053), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  OAI21_X1  g0865(.A(new_n788), .B1(new_n706), .B2(new_n799), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT114), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1066), .B(new_n1067), .ZN(new_n1068));
  OAI211_X1 g0868(.A(KEYINPUT116), .B(new_n864), .C1(new_n794), .C2(new_n703), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n792), .A2(new_n793), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n703), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n863), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT116), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n703), .A2(new_n799), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n863), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1068), .B(new_n1069), .C1(new_n1072), .C2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n785), .B1(new_n686), .B2(new_n800), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n864), .B1(new_n703), .B2(new_n799), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(new_n863), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1076), .A2(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n868), .A2(new_n869), .A3(new_n884), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n857), .ZN(new_n1086));
  OAI211_X1 g0886(.A(KEYINPUT115), .B(new_n1086), .C1(new_n1077), .C2(new_n864), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT115), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n865), .B2(new_n857), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n856), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n855), .B(new_n1086), .C1(new_n1068), .C2(new_n864), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1091), .A2(new_n1080), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1080), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1085), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1080), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1080), .A3(new_n1092), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1077), .B1(new_n1080), .B2(new_n1079), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1072), .A2(KEYINPUT116), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n864), .B1(new_n794), .B2(new_n703), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1097), .B2(new_n1073), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1100), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n870), .A2(new_n885), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1098), .A2(new_n1099), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1095), .A2(new_n1109), .A3(new_n676), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1098), .A2(new_n712), .A3(new_n1099), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n288), .B1(new_n744), .B2(G125), .ZN(new_n1112));
  OR3_X1    g0912(.A1(new_n724), .A2(KEYINPUT53), .A3(new_n450), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT53), .B1(new_n724), .B2(new_n450), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  XOR2_X1   g0915(.A(KEYINPUT54), .B(G143), .Z(new_n1116));
  AOI22_X1  g0916(.A1(new_n733), .A2(G128), .B1(new_n741), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n917), .A2(G50), .B1(new_n727), .B2(G132), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(new_n812), .C2(new_n826), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1115), .B(new_n1119), .C1(G159), .C2(new_n759), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n822), .B1(G107), .B2(new_n811), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n728), .A2(new_n559), .B1(new_n740), .B2(new_n475), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n732), .A2(new_n747), .B1(new_n743), .B2(new_n750), .ZN(new_n1123));
  NOR4_X1   g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n286), .A4(new_n763), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1121), .A2(new_n1046), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n719), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n805), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n713), .B1(new_n1127), .B2(new_n305), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT117), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1126), .B(new_n1129), .C1(new_n856), .C2(new_n770), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1110), .A2(new_n1111), .A3(new_n1130), .ZN(G378));
  XNOR2_X1  g0931(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n463), .A2(KEYINPUT55), .A3(new_n466), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT55), .B1(new_n463), .B2(new_n466), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n464), .A2(new_n652), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n463), .A2(new_n466), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT55), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1139), .B1(new_n1142), .B2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1133), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1137), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1139), .A3(new_n1134), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n1146), .A3(new_n1132), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n883), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1150), .A2(G330), .A3(new_n878), .A4(new_n880), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n867), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1149), .A2(new_n1151), .A3(new_n866), .A4(new_n858), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(KEYINPUT121), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT121), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1152), .A2(new_n1156), .A3(new_n867), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n712), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G58), .A2(new_n917), .B1(new_n744), .B2(G283), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n479), .B2(new_n728), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n288), .A2(new_n261), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n732), .A2(new_n559), .B1(new_n764), .B2(new_n471), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1161), .A2(new_n1018), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1164), .B(new_n901), .C1(new_n1020), .C2(new_n740), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(G33), .A2(G41), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(G50), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1165), .A2(new_n1166), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(G128), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n728), .A2(new_n1170), .B1(new_n740), .B2(new_n826), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G125), .B2(new_n733), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n905), .A2(new_n1116), .B1(new_n736), .B2(G132), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n450), .C2(new_n754), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT118), .B(G124), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1167), .B1(new_n743), .B2(new_n1177), .C1(new_n281), .C2(new_n748), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT119), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1169), .B1(new_n1166), .B2(new_n1165), .C1(new_n1175), .C2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n719), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n714), .B1(new_n211), .B2(new_n805), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(new_n1150), .C2(new_n770), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1159), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1186), .A2(KEYINPUT57), .ZN(new_n1187));
  NOR3_X1   g0987(.A1(new_n1093), .A2(new_n1094), .A3(new_n1085), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1084), .B(KEYINPUT122), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n676), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1189), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1109), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT57), .B1(new_n1193), .B2(new_n1158), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1191), .B2(new_n1194), .ZN(G375));
  AOI21_X1  g0995(.A(new_n711), .B1(new_n1076), .B2(new_n1082), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n728), .A2(new_n826), .B1(new_n724), .B2(new_n281), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n288), .B(new_n1197), .C1(G58), .C2(new_n917), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n759), .A2(G50), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n811), .A2(new_n1116), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n740), .A2(new_n450), .B1(new_n743), .B2(new_n1170), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G132), .B2(new_n733), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n728), .A2(new_n747), .B1(new_n743), .B2(new_n725), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n740), .A2(new_n479), .B1(new_n724), .B2(new_n471), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n288), .B1(new_n732), .B2(new_n750), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n205), .B2(new_n749), .C1(new_n812), .C2(new_n559), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1020), .A2(new_n754), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n719), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n714), .B1(new_n202), .B2(new_n805), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n863), .C2(new_n770), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT123), .B1(new_n1196), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT123), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1216), .B(new_n1213), .C1(new_n1106), .C2(new_n711), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(new_n1085), .A3(new_n981), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(G381));
  INV_X1    g1021(.A(G384), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(G393), .A2(G396), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1111), .A2(new_n1130), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n677), .B1(new_n1227), .B2(new_n1085), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1226), .B1(new_n1228), .B2(new_n1109), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G375), .A2(KEYINPUT124), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1225), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(G407));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  INV_X1    g1034(.A(new_n983), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1053), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n781), .B1(new_n989), .B2(new_n1024), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n984), .B1(new_n1223), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1223), .A2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1064), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1235), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1064), .A2(new_n1239), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n983), .C1(new_n1064), .C2(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1185), .B(G378), .C1(new_n1191), .C2(new_n1194), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1186), .A2(new_n712), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1184), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1109), .B2(new_n1192), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1249), .B1(new_n1251), .B2(new_n981), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT125), .B1(new_n1252), .B2(G378), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n981), .B(new_n1158), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1249), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1229), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1247), .A2(new_n1253), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n653), .A2(G213), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n653), .A2(G213), .A3(G2897), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n677), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1218), .A2(new_n1268), .A3(G384), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1218), .B2(new_n1268), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1263), .B1(new_n1271), .B2(KEYINPUT126), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1273), .B(new_n1262), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1272), .A2(new_n1274), .B1(KEYINPUT126), .B2(new_n1271), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1261), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1259), .A2(new_n1271), .A3(new_n1260), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT62), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(KEYINPUT62), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT61), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1246), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1271), .A2(KEYINPUT126), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1218), .A2(new_n1268), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1222), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1218), .A2(new_n1268), .A3(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1262), .B1(new_n1287), .B2(new_n1273), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1274), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1260), .B2(new_n1259), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1277), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT63), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1243), .A2(new_n1280), .A3(new_n1245), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT127), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1243), .A2(KEYINPUT127), .A3(new_n1245), .A4(new_n1280), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1277), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1282), .A2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1229), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1247), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1271), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1246), .ZN(G402));
endmodule


