//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G104), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n188), .A2(new_n193), .A3(new_n189), .A4(G104), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n191), .A2(new_n192), .A3(new_n194), .A4(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT82), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n190), .A2(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n199), .A2(new_n200), .A3(new_n192), .A4(new_n194), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n192), .B1(new_n199), .B2(new_n194), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT2), .B(G113), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(G116), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  INV_X1    g023(.A(G116), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G119), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n208), .B2(G119), .ZN(new_n213));
  INV_X1    g027(.A(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n212), .A2(new_n215), .B1(new_n203), .B2(new_n204), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n189), .A2(G104), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n192), .B1(new_n217), .B2(new_n196), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n198), .B2(new_n201), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(KEYINPUT5), .ZN(new_n220));
  INV_X1    g034(.A(G113), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n221), .B1(new_n211), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n220), .A2(new_n223), .B1(new_n213), .B2(new_n214), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n206), .A2(new_n216), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G110), .B(G122), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT6), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n206), .A2(new_n216), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(new_n224), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT86), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n232), .A3(new_n226), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n227), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NOR3_X1   g048(.A1(new_n225), .A2(KEYINPUT6), .A3(new_n226), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G143), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n238), .B2(G146), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(KEYINPUT64), .A3(G143), .ZN(new_n246));
  INV_X1    g060(.A(new_n241), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n239), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G125), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n237), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G128), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n240), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n245), .A2(new_n246), .A3(new_n256), .A4(new_n239), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n250), .B1(new_n261), .B2(G125), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G224), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n262), .B(new_n264), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n234), .A2(new_n235), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n267));
  INV_X1    g081(.A(new_n264), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n267), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n250), .B(new_n270), .C1(new_n261), .C2(G125), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n226), .B(KEYINPUT8), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT88), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n219), .B2(new_n224), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n223), .B(KEYINPUT87), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n220), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n219), .A2(new_n277), .A3(new_n215), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n219), .A2(new_n224), .A3(new_n274), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n273), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AND4_X1   g095(.A1(new_n232), .A2(new_n228), .A3(new_n229), .A4(new_n226), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n232), .B1(new_n225), .B2(new_n226), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n272), .B(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n187), .B1(new_n266), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n269), .A2(new_n271), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(new_n231), .B2(new_n233), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n291), .B2(new_n281), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n228), .A2(new_n229), .ZN(new_n294));
  INV_X1    g108(.A(new_n226), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n282), .B2(new_n283), .ZN(new_n297));
  INV_X1    g111(.A(new_n235), .ZN(new_n298));
  INV_X1    g112(.A(new_n265), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n292), .A2(new_n300), .A3(KEYINPUT89), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n287), .A2(new_n289), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n292), .A2(new_n300), .A3(new_n288), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  NOR2_X1   g119(.A1(G237), .A2(G953), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT18), .B(G131), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G140), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G146), .ZN(new_n316));
  XNOR2_X1  g130(.A(G125), .B(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n236), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n263), .A3(G214), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n238), .ZN(new_n322));
  NAND2_X1  g136(.A1(KEYINPUT18), .A2(G131), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n307), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n310), .A2(new_n319), .A3(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(G113), .B(G122), .Z(new_n326));
  XOR2_X1   g140(.A(KEYINPUT92), .B(G104), .Z(new_n327));
  XOR2_X1   g141(.A(new_n326), .B(new_n327), .Z(new_n328));
  OAI21_X1  g142(.A(G131), .B1(new_n308), .B2(new_n309), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n322), .A2(new_n331), .A3(new_n307), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT16), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n311), .A3(G125), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n315), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n236), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT17), .B(G131), .C1(new_n308), .C2(new_n309), .ZN(new_n339));
  OAI211_X1 g153(.A(G146), .B(new_n336), .C1(new_n315), .C2(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n325), .B(new_n328), .C1(new_n334), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n333), .A2(new_n338), .A3(new_n340), .A4(new_n339), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n345), .A2(KEYINPUT93), .A3(new_n328), .A4(new_n325), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT91), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT19), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n315), .B2(KEYINPUT90), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n317), .A2(new_n350), .A3(KEYINPUT19), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n352), .B2(new_n236), .ZN(new_n353));
  AOI211_X1 g167(.A(KEYINPUT91), .B(G146), .C1(new_n349), .C2(new_n351), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n329), .A2(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n340), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n325), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n328), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n344), .A2(new_n346), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(G475), .A2(G902), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT20), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n344), .A2(new_n346), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n358), .A2(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n361), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n328), .B1(new_n345), .B2(new_n325), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n369), .B1(new_n344), .B2(new_n346), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(G902), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT94), .B(G475), .Z(new_n372));
  AOI22_X1  g186(.A1(new_n363), .A2(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  INV_X1    g188(.A(G217), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(G953), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n238), .A2(G128), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n255), .A2(G143), .ZN(new_n378));
  INV_X1    g192(.A(G134), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n378), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n383));
  INV_X1    g197(.A(new_n377), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(KEYINPUT13), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n377), .A2(KEYINPUT95), .A3(new_n381), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n208), .A2(G122), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n210), .A2(G122), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n189), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n189), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  OAI221_X1 g206(.A(new_n380), .B1(new_n387), .B2(new_n379), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n377), .A2(new_n378), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G134), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n380), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n388), .A2(new_n397), .A3(new_n389), .ZN(new_n398));
  OAI21_X1  g212(.A(G107), .B1(new_n388), .B2(new_n397), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n390), .B(new_n396), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n376), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n391), .A2(new_n392), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n380), .B1(new_n387), .B2(new_n379), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n400), .B(new_n376), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n285), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G478), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n400), .B1(new_n402), .B2(new_n403), .ZN(new_n410));
  INV_X1    g224(.A(new_n376), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(G902), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  INV_X1    g227(.A(new_n408), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n409), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n373), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(G234), .A2(G237), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n419), .A2(G952), .A3(new_n263), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(G902), .A3(G953), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT96), .Z(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(G898), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n304), .A2(new_n305), .A3(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT26), .B(G101), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n306), .A2(G210), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n212), .A2(new_n215), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n379), .B2(G137), .ZN(new_n435));
  INV_X1    g249(.A(G137), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT11), .A3(G134), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n379), .A2(G137), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G131), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n435), .A2(new_n437), .A3(new_n331), .A4(new_n438), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(KEYINPUT65), .A3(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n243), .A2(new_n248), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n444), .A3(G131), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n438), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n379), .A2(G137), .ZN(new_n449));
  OAI21_X1  g263(.A(G131), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n441), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n261), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n433), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n249), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n248), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(new_n457), .A3(new_n442), .A4(new_n445), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n433), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT28), .B1(new_n454), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n453), .A2(new_n458), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n432), .B1(new_n463), .B2(KEYINPUT72), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n453), .A2(new_n465), .A3(new_n458), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT28), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n431), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n246), .A2(new_n239), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(KEYINPUT66), .A3(new_n245), .A4(new_n256), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n257), .A2(new_n258), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n451), .B1(new_n473), .B2(new_n254), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n469), .B1(new_n446), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n453), .A2(KEYINPUT30), .A3(new_n458), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n432), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n476), .A3(new_n479), .A4(new_n432), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n431), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n459), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(KEYINPUT31), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT31), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n486), .B(new_n483), .C1(new_n478), .C2(new_n480), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n468), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G472), .A2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT73), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n464), .A2(new_n466), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n482), .B1(new_n497), .B2(new_n461), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n481), .A2(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n486), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n481), .A2(KEYINPUT31), .A3(new_n484), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n490), .A2(new_n493), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT75), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n463), .A2(KEYINPUT72), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n506), .A2(new_n433), .A3(new_n466), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n461), .B(new_n482), .C1(new_n507), .C2(KEYINPUT28), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT29), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n460), .B1(new_n478), .B2(new_n480), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n508), .B(new_n509), .C1(new_n482), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT74), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n463), .A2(new_n432), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n496), .B1(new_n513), .B2(new_n459), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n431), .A2(new_n509), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n467), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n512), .B1(new_n517), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n514), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n497), .A2(new_n519), .A3(new_n515), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT74), .A3(new_n285), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(G472), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n488), .A2(new_n524), .A3(new_n503), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n494), .A2(new_n505), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  INV_X1    g341(.A(G119), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n527), .B1(new_n528), .B2(G128), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(G128), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n255), .A2(KEYINPUT23), .A3(G119), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G110), .ZN(new_n533));
  INV_X1    g347(.A(G110), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G110), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n528), .B2(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n255), .A2(KEYINPUT76), .A3(G119), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n538), .A2(new_n540), .A3(new_n541), .A4(new_n530), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n338), .B2(new_n340), .ZN(new_n544));
  INV_X1    g358(.A(new_n532), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n541), .A3(new_n530), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n545), .A2(new_n534), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n340), .A2(new_n318), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT77), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n338), .A2(new_n340), .ZN(new_n552));
  INV_X1    g366(.A(new_n543), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n340), .A2(new_n318), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n546), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(G110), .B2(new_n532), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n551), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n554), .A2(new_n558), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(new_n564), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n552), .A2(new_n553), .B1(new_n555), .B2(new_n557), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT78), .A3(new_n563), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n565), .A2(new_n568), .A3(new_n285), .A4(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT78), .B1(new_n569), .B2(new_n563), .ZN(new_n574));
  AND4_X1   g388(.A1(KEYINPUT78), .A2(new_n554), .A3(new_n558), .A4(new_n563), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n576), .A2(KEYINPUT25), .A3(new_n285), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n375), .B1(G234), .B2(new_n285), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT79), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n582), .A3(new_n579), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n576), .A2(new_n565), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n579), .A2(G902), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT80), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n581), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n374), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G469), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  INV_X1    g408(.A(G227), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(G953), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n594), .B(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n470), .A2(new_n245), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n255), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n599));
  OAI22_X1  g413(.A1(new_n259), .A2(new_n260), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n219), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n199), .A2(new_n194), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(new_n204), .A3(G101), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n456), .A2(new_n605), .A3(new_n457), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n206), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n442), .A2(new_n445), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n261), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n603), .A2(new_n607), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT83), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n602), .B1(new_n473), .B2(new_n254), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n606), .A2(new_n206), .B1(new_n613), .B2(new_n219), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n614), .A2(KEYINPUT83), .A3(new_n608), .A4(new_n603), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n597), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n601), .B1(new_n261), .B2(new_n219), .ZN(new_n617));
  INV_X1    g431(.A(new_n608), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n597), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n615), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT84), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n202), .A2(new_n205), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n456), .A2(new_n605), .A3(new_n457), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n609), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT10), .B1(new_n219), .B2(new_n600), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n614), .A2(KEYINPUT84), .A3(new_n603), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n618), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n623), .B1(new_n624), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT85), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n622), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n614), .A2(new_n603), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n608), .B1(new_n636), .B2(new_n625), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(new_n631), .B1(new_n612), .B2(new_n615), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n638), .A2(KEYINPUT85), .A3(new_n623), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n593), .B(new_n285), .C1(new_n635), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n621), .A2(new_n624), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n641), .A2(new_n597), .B1(new_n632), .B2(new_n616), .ZN(new_n642));
  OAI21_X1  g456(.A(G469), .B1(new_n642), .B2(G902), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n592), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n426), .A2(new_n526), .A3(new_n590), .A4(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT97), .B(G101), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G3));
  INV_X1    g461(.A(new_n492), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n488), .A2(KEYINPUT98), .A3(new_n285), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n649), .A2(G472), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n488), .A2(new_n285), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n648), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n592), .B(new_n589), .C1(new_n640), .C2(new_n643), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n292), .A2(new_n300), .A3(new_n288), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n288), .B1(new_n292), .B2(new_n300), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n305), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n363), .A2(new_n368), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n372), .B1(new_n370), .B2(G902), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT33), .B1(new_n401), .B2(new_n405), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n412), .A2(new_n664), .A3(new_n404), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(G478), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n407), .A2(new_n285), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n413), .B2(new_n407), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n659), .A2(new_n671), .A3(new_n424), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n360), .A2(KEYINPUT20), .A3(new_n362), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n367), .B1(new_n366), .B2(new_n361), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n416), .B(new_n661), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n677), .B1(new_n680), .B2(new_n424), .ZN(new_n681));
  INV_X1    g495(.A(new_n424), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n373), .A2(KEYINPUT99), .A3(new_n682), .A4(new_n416), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n676), .B1(new_n684), .B2(new_n659), .ZN(new_n685));
  INV_X1    g499(.A(new_n305), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n292), .A2(new_n300), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n289), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n688), .B2(new_n303), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(KEYINPUT100), .A3(new_n681), .A4(new_n683), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n656), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT35), .B(G107), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n551), .A2(new_n560), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(KEYINPUT36), .A3(new_n564), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n564), .A2(KEYINPUT36), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n551), .B2(new_n560), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n695), .B1(new_n700), .B2(new_n586), .ZN(new_n701));
  INV_X1    g515(.A(new_n700), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT101), .A3(new_n587), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n581), .A2(new_n583), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n654), .A2(new_n426), .A3(new_n644), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT37), .B(G110), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G12));
  AOI211_X1 g521(.A(new_n592), .B(new_n659), .C1(new_n640), .C2(new_n643), .ZN(new_n708));
  INV_X1    g522(.A(new_n704), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n488), .A2(new_n524), .A3(new_n503), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n524), .B1(new_n488), .B2(new_n503), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n493), .A2(new_n492), .B1(new_n522), .B2(G472), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(G900), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n420), .B1(new_n422), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n680), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n708), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT102), .B(G128), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G30));
  AOI21_X1  g534(.A(new_n482), .B1(new_n513), .B2(new_n459), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n481), .B2(new_n484), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n722), .B2(G902), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n494), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n712), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n304), .A2(KEYINPUT38), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT38), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n302), .A2(new_n728), .A3(new_n303), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n373), .A2(new_n417), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n305), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n726), .A2(new_n730), .A3(new_n704), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n716), .B(KEYINPUT39), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n644), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT103), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n733), .A2(new_n740), .A3(new_n736), .A4(new_n737), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n238), .ZN(G45));
  INV_X1    g557(.A(new_n671), .ZN(new_n744));
  INV_X1    g558(.A(new_n716), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n708), .A2(new_n714), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  AOI21_X1  g563(.A(new_n589), .B1(new_n712), .B2(new_n713), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n285), .B1(new_n635), .B2(new_n639), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n752), .A2(new_n591), .A3(new_n640), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(new_n753), .A3(new_n672), .ZN(new_n754));
  XNOR2_X1  g568(.A(KEYINPUT41), .B(G113), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G15));
  NAND2_X1  g570(.A1(new_n526), .A2(new_n590), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n752), .A2(new_n591), .A3(new_n640), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n691), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NAND3_X1  g575(.A1(new_n526), .A2(new_n425), .A3(new_n704), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n752), .A2(new_n591), .A3(new_n640), .A4(new_n689), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n528), .ZN(G21));
  OAI21_X1  g579(.A(G472), .B1(new_n502), .B2(G902), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n431), .B1(new_n467), .B2(new_n514), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n485), .B2(new_n487), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n491), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n590), .A2(new_n766), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n689), .A2(new_n682), .A3(new_n731), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n753), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  NOR2_X1   g588(.A1(new_n763), .A2(new_n746), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n704), .A3(new_n769), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g592(.A1(new_n651), .A2(G472), .B1(new_n491), .B2(new_n768), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(KEYINPUT104), .A3(new_n704), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G125), .ZN(G27));
  AND2_X1   g597(.A1(new_n303), .A2(new_n305), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n302), .A2(new_n784), .A3(new_n591), .ZN(new_n785));
  NAND2_X1  g599(.A1(G469), .A2(G902), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT105), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n642), .B2(G469), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n785), .B1(new_n640), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n488), .A2(new_n503), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n589), .B1(new_n713), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n790), .A2(new_n792), .A3(KEYINPUT42), .A4(new_n747), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  INV_X1    g608(.A(new_n785), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n640), .A2(new_n789), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n526), .A2(new_n795), .A3(new_n590), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n794), .B1(new_n797), .B2(new_n747), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n750), .A2(new_n790), .A3(new_n794), .A4(new_n747), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n793), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G131), .ZN(G33));
  NAND3_X1  g617(.A1(new_n750), .A2(new_n790), .A3(new_n717), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND2_X1  g619(.A1(new_n302), .A2(new_n784), .ZN(new_n806));
  INV_X1    g620(.A(new_n654), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT107), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n373), .B(new_n670), .C1(new_n808), .C2(KEYINPUT43), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n662), .A2(new_n669), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n807), .A2(new_n704), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n806), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  INV_X1    g630(.A(new_n734), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n641), .A2(new_n597), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n616), .A2(new_n632), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT45), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n593), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n642), .A2(KEYINPUT45), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n787), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(KEYINPUT46), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n640), .B1(new_n826), .B2(KEYINPUT46), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n591), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n816), .A2(new_n817), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT108), .B(G137), .Z(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(G39));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(KEYINPUT47), .B(new_n591), .C1(new_n827), .C2(new_n828), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR4_X1   g650(.A1(new_n526), .A2(new_n746), .A3(new_n590), .A4(new_n806), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G140), .ZN(G42));
  NAND2_X1  g653(.A1(new_n263), .A2(G952), .ZN(new_n840));
  INV_X1    g654(.A(new_n763), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n812), .A2(new_n420), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n770), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n420), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n758), .A2(new_n845), .A3(new_n806), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n726), .A3(new_n590), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n844), .B1(new_n847), .B2(new_n671), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n846), .A2(new_n812), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n792), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT48), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n781), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n373), .A2(new_n669), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n847), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n640), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT85), .B1(new_n638), .B2(new_n623), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n633), .A2(new_n634), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n622), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n593), .B1(new_n863), .B2(new_n285), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n592), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n834), .A2(new_n835), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n842), .A2(new_n770), .A3(new_n806), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n856), .B(new_n859), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n758), .B2(new_n305), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n753), .A2(KEYINPUT114), .A3(new_n686), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n730), .A3(new_n872), .A4(new_n843), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT50), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n850), .B(new_n855), .C1(new_n869), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n866), .B(KEYINPUT113), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n834), .A2(new_n835), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n859), .B1(new_n880), .B2(new_n868), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n876), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n856), .ZN(new_n883));
  AOI211_X1 g697(.A(KEYINPUT116), .B(KEYINPUT51), .C1(new_n881), .C2(new_n876), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT104), .B1(new_n779), .B2(new_n704), .ZN(new_n886));
  AND4_X1   g700(.A1(KEYINPUT104), .A2(new_n766), .A3(new_n704), .A4(new_n769), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n747), .B(new_n790), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n640), .A2(new_n643), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n745), .A2(new_n591), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n806), .A2(new_n418), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n714), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n804), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n424), .B1(new_n671), .B2(new_n680), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n304), .A2(new_n305), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n654), .A2(new_n655), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n705), .A2(new_n645), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n802), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n526), .A2(new_n425), .A3(new_n704), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n759), .A2(new_n691), .B1(new_n900), .B2(new_n841), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n758), .A2(new_n770), .A3(new_n771), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n759), .B2(new_n672), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT111), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT111), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n865), .A2(new_n526), .A3(new_n590), .A4(new_n591), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n685), .A2(new_n690), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n906), .A2(new_n907), .B1(new_n762), .B2(new_n763), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n754), .A2(new_n773), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n904), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n708), .B(new_n714), .C1(new_n717), .C2(new_n747), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n659), .A2(new_n417), .A3(new_n373), .A4(new_n890), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n725), .A2(new_n709), .A3(new_n796), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n782), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT52), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n899), .A2(new_n911), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT53), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(KEYINPUT54), .C1(new_n918), .C2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n802), .A2(new_n904), .A3(new_n898), .A4(new_n910), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n915), .B(KEYINPUT52), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n901), .A2(new_n903), .A3(KEYINPUT53), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n899), .A2(new_n917), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  OAI22_X1  g744(.A1(new_n885), .A2(new_n930), .B1(G952), .B2(G953), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n590), .A2(new_n591), .A3(new_n305), .A4(new_n810), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT109), .ZN(new_n933));
  INV_X1    g747(.A(new_n865), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(KEYINPUT49), .B2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT110), .Z(new_n936));
  OAI211_X1 g750(.A(new_n726), .B(new_n730), .C1(KEYINPUT49), .C2(new_n934), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(G75));
  AOI21_X1  g752(.A(new_n299), .B1(new_n297), .B2(new_n298), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n266), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n285), .B1(new_n925), .B2(new_n928), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(G210), .ZN(new_n944));
  OR2_X1    g758(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n263), .A2(G952), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n944), .A2(new_n942), .A3(new_n945), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G51));
  AOI211_X1 g765(.A(new_n285), .B(new_n824), .C1(new_n925), .C2(new_n928), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n787), .B(KEYINPUT57), .Z(new_n953));
  AND3_X1   g767(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n926), .B1(new_n925), .B2(new_n928), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n952), .B1(new_n956), .B2(new_n863), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT120), .B1(new_n957), .B2(new_n947), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT120), .ZN(new_n959));
  INV_X1    g773(.A(new_n863), .ZN(new_n960));
  AND4_X1   g774(.A1(new_n802), .A2(new_n904), .A3(new_n898), .A4(new_n910), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n921), .B1(new_n961), .B2(new_n917), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n899), .A2(new_n917), .A3(new_n927), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT54), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n929), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n960), .B1(new_n965), .B2(new_n953), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n959), .B(new_n948), .C1(new_n966), .C2(new_n952), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n958), .A2(new_n967), .ZN(G54));
  NAND3_X1  g782(.A1(new_n943), .A2(KEYINPUT58), .A3(G475), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n969), .A2(KEYINPUT121), .A3(new_n360), .ZN(new_n970));
  OAI21_X1  g784(.A(KEYINPUT121), .B1(new_n969), .B2(new_n360), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n947), .B1(new_n969), .B2(new_n360), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G60));
  AND2_X1   g787(.A1(new_n663), .A2(new_n665), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n667), .B(KEYINPUT59), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n965), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n948), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n930), .A2(new_n977), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT122), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n974), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n976), .B1(new_n922), .B2(new_n929), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT122), .B1(new_n983), .B2(new_n975), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n982), .B2(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n925), .B2(new_n928), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n584), .B(KEYINPUT124), .Z(new_n990));
  AOI21_X1  g804(.A(new_n947), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n988), .A2(KEYINPUT123), .A3(new_n702), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT123), .B1(new_n988), .B2(new_n702), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n991), .B(KEYINPUT61), .C1(new_n992), .C2(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  INV_X1    g812(.A(new_n423), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n263), .B1(new_n999), .B2(G224), .ZN(new_n1000));
  INV_X1    g814(.A(new_n897), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n911), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n263), .ZN(new_n1003));
  OAI22_X1  g817(.A1(new_n234), .A2(new_n235), .B1(G898), .B2(new_n263), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(G69));
  AOI21_X1  g819(.A(new_n806), .B1(new_n671), .B2(new_n680), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n750), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n830), .B(new_n838), .C1(new_n735), .C2(new_n1007), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n782), .A2(new_n912), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(new_n741), .A3(new_n739), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT126), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR3_X1   g831(.A1(new_n1013), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n475), .A2(new_n476), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(new_n352), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g836(.A1(new_n836), .A2(new_n837), .B1(new_n717), .B2(new_n797), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n792), .A2(new_n689), .A3(new_n731), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n816), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n829), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1025), .A2(new_n734), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1023), .A2(new_n1027), .A3(new_n802), .A4(new_n1012), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1021), .ZN(new_n1030));
  AOI21_X1  g844(.A(G953), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1030), .A2(G227), .ZN(new_n1032));
  AOI211_X1 g846(.A(new_n715), .B(new_n263), .C1(new_n1021), .C2(new_n595), .ZN(new_n1033));
  AOI22_X1  g847(.A1(new_n1022), .A2(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(G72));
  NAND2_X1  g848(.A1(G472), .A2(G902), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1035), .B(KEYINPUT63), .Z(new_n1036));
  OAI21_X1  g850(.A(new_n1036), .B1(new_n1028), .B2(new_n1002), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n510), .B(KEYINPUT127), .Z(new_n1038));
  INV_X1    g852(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1037), .A2(new_n431), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1036), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n510), .A2(new_n482), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1042), .B2(new_n499), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n919), .B(new_n1043), .C1(new_n918), .C2(new_n921), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1040), .A2(new_n948), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1036), .B1(new_n1019), .B2(new_n1002), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1039), .A2(new_n431), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(G57));
endmodule


