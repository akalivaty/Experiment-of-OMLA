//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n813, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  OR3_X1    g001(.A1(new_n202), .A2(G29gat), .A3(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND4_X1  g004(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT86), .A4(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207));
  AND2_X1   g006(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(KEYINPUT15), .ZN(new_n209));
  OR3_X1    g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(KEYINPUT15), .A3(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT16), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G8gat), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n218), .A2(G8gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n219), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n212), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n221), .A2(new_n227), .A3(KEYINPUT18), .A4(new_n228), .ZN(new_n232));
  INV_X1    g031(.A(new_n226), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n233), .A2(new_n224), .A3(new_n211), .A4(new_n210), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n227), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n228), .B(KEYINPUT88), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(KEYINPUT13), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G169gat), .B(G197gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT12), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n239), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n238), .A3(new_n232), .A4(new_n245), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(G71gat), .B(G99gat), .Z(new_n251));
  XNOR2_X1  g050(.A(G15gat), .B(G43gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G227gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(G134gat), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G113gat), .B2(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(G113gat), .A2(G120gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n256), .A2(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n257), .A2(G127gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n255), .A2(G134gat), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n266), .A2(new_n261), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n273));
  NOR3_X1   g072(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n273), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  INV_X1    g076(.A(G169gat), .ZN(new_n278));
  INV_X1    g077(.A(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n281));
  OAI211_X1 g080(.A(KEYINPUT70), .B(new_n271), .C1(new_n276), .C2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n273), .A2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n280), .A2(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n274), .A2(new_n275), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT70), .B1(new_n287), .B2(new_n271), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT27), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n292));
  INV_X1    g091(.A(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT27), .B(G183gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NOR3_X1   g097(.A1(new_n283), .A2(new_n288), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n271), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT65), .ZN(new_n302));
  AND2_X1   g101(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G190gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT23), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(G169gat), .B2(G176gat), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n313), .A2(KEYINPUT25), .A3(new_n315), .A4(new_n272), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n272), .B1(new_n312), .B2(KEYINPUT23), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n314), .A2(G169gat), .A3(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT64), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT64), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n313), .A2(new_n321), .A3(new_n315), .A4(new_n272), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n305), .B1(new_n303), .B2(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n301), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT25), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n311), .A2(new_n317), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n270), .B1(new_n299), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n326), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n301), .B(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n317), .B1(new_n331), .B2(new_n309), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n271), .B1(new_n276), .B2(new_n281), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n298), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n282), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n263), .A2(new_n269), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n254), .B1(new_n328), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT33), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n253), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n254), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n339), .B1(new_n333), .B2(new_n338), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n342), .B1(new_n253), .B2(KEYINPUT33), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n328), .A2(new_n254), .A3(new_n340), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT34), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n328), .A2(KEYINPUT34), .A3(new_n254), .A4(new_n340), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT72), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n343), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n359), .A2(new_n253), .B1(new_n349), .B2(new_n350), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT71), .B1(new_n360), .B2(new_n362), .ZN(new_n364));
  AND4_X1   g163(.A1(KEYINPUT71), .A2(new_n362), .A3(new_n345), .A4(new_n351), .ZN(new_n365));
  OAI22_X1  g164(.A1(new_n358), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT36), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n357), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n345), .A3(new_n351), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT36), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G211gat), .B(G218gat), .Z(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n386), .A2(new_n381), .A3(new_n382), .A4(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(G148gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G141gat), .ZN(new_n392));
  INV_X1    g191(.A(G141gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(G148gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT74), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(G148gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(G141gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G155gat), .A2(G162gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT2), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G155gat), .ZN(new_n403));
  INV_X1    g202(.A(G162gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n400), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT75), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n391), .B2(G141gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT75), .A3(G148gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n397), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n400), .B1(new_n405), .B2(KEYINPUT2), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n402), .A2(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n377), .B1(new_n390), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G141gat), .B(G148gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n401), .B1(new_n415), .B2(new_n398), .ZN(new_n416));
  INV_X1    g215(.A(new_n399), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n407), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(new_n412), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n385), .B2(new_n387), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT79), .B(new_n420), .C1(new_n421), .C2(KEYINPUT3), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n376), .B1(new_n414), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n418), .A2(new_n425), .A3(new_n419), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT76), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n428), .A3(new_n425), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n424), .B1(new_n430), .B2(new_n388), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n413), .B2(new_n425), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n433), .B1(G155gat), .B2(G162gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n396), .A2(new_n397), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n434), .B1(new_n435), .B2(KEYINPUT74), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n406), .B1(new_n436), .B2(new_n399), .ZN(new_n437));
  INV_X1    g236(.A(new_n419), .ZN(new_n438));
  NOR4_X1   g237(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT76), .A4(KEYINPUT3), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n389), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n388), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n431), .A3(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n430), .A2(new_n388), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n390), .A2(new_n413), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n376), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n443), .B2(new_n446), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n375), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n443), .A2(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(G22gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n448), .A3(new_n374), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n271), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n275), .B1(new_n312), .B2(new_n277), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n273), .A2(new_n272), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n459), .B1(new_n462), .B2(new_n286), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n337), .B1(new_n463), .B2(KEYINPUT70), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n313), .A2(new_n272), .A3(new_n315), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(KEYINPUT64), .B1(new_n323), .B2(new_n301), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT25), .B1(new_n466), .B2(new_n322), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n316), .B1(new_n302), .B2(new_n310), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n464), .A2(new_n283), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n458), .B1(new_n469), .B2(new_n389), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n457), .B1(new_n333), .B2(new_n338), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n441), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G64gat), .ZN(new_n474));
  INV_X1    g273(.A(G92gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n298), .B1(new_n334), .B2(new_n335), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n282), .A2(new_n477), .B1(new_n329), .B2(new_n332), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n457), .B1(new_n478), .B2(KEYINPUT29), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n469), .A2(new_n458), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n388), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n472), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n472), .A2(new_n481), .A3(KEYINPUT30), .A4(new_n476), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n470), .A2(new_n441), .A3(new_n471), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n388), .B1(new_n479), .B2(new_n480), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n484), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n339), .B1(new_n420), .B2(KEYINPUT3), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(new_n432), .B2(new_n439), .ZN(new_n493));
  NAND2_X1  g292(.A1(G225gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n413), .B2(new_n339), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n497), .B2(KEYINPUT77), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n418), .A2(new_n339), .A3(new_n419), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n413), .A2(new_n496), .A3(new_n339), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n437), .A2(new_n438), .A3(new_n270), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n339), .B1(new_n418), .B2(new_n419), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n495), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n505), .B1(new_n508), .B2(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n270), .B1(new_n437), .B2(new_n438), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n494), .B1(new_n510), .B2(new_n499), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT5), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n511), .A2(KEYINPUT78), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n504), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G1gat), .B(G29gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT0), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G57gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G85gat), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n516), .B(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G85gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n427), .A2(new_n429), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n524), .A2(new_n492), .B1(new_n500), .B2(new_n501), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n514), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n505), .A3(KEYINPUT5), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT78), .B1(new_n511), .B2(new_n512), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(new_n504), .B1(new_n525), .B2(new_n526), .ZN(new_n533));
  INV_X1    g332(.A(new_n523), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n528), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n525), .A2(new_n526), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n514), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n491), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n368), .A2(new_n371), .B1(new_n456), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT37), .B1(new_n487), .B2(new_n488), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT38), .ZN(new_n543));
  XNOR2_X1  g342(.A(KEYINPUT83), .B(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n472), .A2(new_n481), .A3(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n542), .A2(new_n543), .A3(new_n486), .A4(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n535), .A2(new_n546), .A3(new_n482), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT84), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n537), .B2(KEYINPUT6), .ZN(new_n549));
  NOR4_X1   g348(.A1(new_n533), .A2(KEYINPUT84), .A3(new_n529), .A4(new_n534), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(new_n486), .A3(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT38), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n547), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT40), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n500), .A2(new_n501), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n493), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT81), .B1(new_n557), .B2(new_n495), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559));
  AOI211_X1 g358(.A(new_n559), .B(new_n494), .C1(new_n493), .C2(new_n556), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT39), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n506), .A2(new_n507), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n494), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n555), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n559), .B1(new_n525), .B2(new_n494), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n557), .A2(KEYINPUT81), .A3(new_n495), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT39), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT82), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n568), .A2(new_n569), .A3(new_n523), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n562), .B1(new_n558), .B2(new_n560), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT82), .B1(new_n571), .B2(new_n534), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n565), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n537), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n490), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n569), .B1(new_n568), .B2(new_n523), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(KEYINPUT82), .A3(new_n534), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT40), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n554), .B(new_n455), .C1(new_n576), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n541), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n369), .A2(new_n361), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n352), .A2(new_n357), .A3(KEYINPUT72), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT71), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n370), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n362), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n585), .A2(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n538), .A2(KEYINPUT84), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n537), .A2(new_n548), .A3(KEYINPUT6), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n535), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n590), .A2(new_n593), .A3(new_n455), .A4(new_n491), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n369), .A2(new_n370), .ZN(new_n595));
  AOI211_X1 g394(.A(new_n490), .B(new_n595), .C1(new_n454), .C2(new_n451), .ZN(new_n596));
  INV_X1    g395(.A(new_n539), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(new_n584), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n584), .A2(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n250), .B1(new_n583), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n521), .B2(new_n475), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT91), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT7), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT92), .B1(G99gat), .B2(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT8), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT92), .A2(G99gat), .A3(G106gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n613), .A2(new_n614), .B1(new_n521), .B2(new_n475), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G99gat), .B(G106gat), .Z(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT93), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT93), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n622), .B1(new_n618), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n213), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n213), .B(KEYINPUT94), .C1(new_n621), .C2(new_n623), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n618), .A2(new_n619), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n629), .A2(new_n212), .B1(KEYINPUT41), .B2(new_n601), .ZN(new_n630));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT90), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n633), .B1(new_n628), .B2(new_n630), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n605), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n604), .A3(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n519), .A2(G64gat), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n519), .A2(G64gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT89), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  NAND2_X1  g444(.A1(G71gat), .A2(G78gat), .ZN(new_n646));
  OR2_X1    g445(.A1(G71gat), .A2(G78gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT9), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n645), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT9), .B1(new_n642), .B2(new_n641), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n646), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(KEYINPUT21), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G211gat), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n225), .A2(new_n226), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n654), .A2(KEYINPUT21), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G183gat), .ZN(new_n663));
  INV_X1    g462(.A(G183gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n660), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n666));
  NAND2_X1  g465(.A1(G231gat), .A2(G233gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n663), .B2(new_n665), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n659), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n658), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n640), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n620), .A2(new_n653), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n618), .A2(new_n654), .A3(new_n619), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n629), .A2(KEYINPUT95), .A3(KEYINPUT10), .A4(new_n654), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(new_n680), .B2(new_n679), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n678), .B2(new_n680), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT96), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XOR2_X1   g490(.A(new_n690), .B(new_n691), .Z(new_n692));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n687), .A2(KEYINPUT97), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT97), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n685), .A2(new_n696), .A3(new_n686), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n688), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n699));
  INV_X1    g498(.A(new_n692), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n688), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n685), .A2(new_n696), .A3(new_n686), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n696), .B1(new_n685), .B2(new_n686), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT98), .B1(new_n705), .B2(new_n692), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n694), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n677), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n600), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n539), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n215), .ZN(G1324gat));
  INV_X1    g510(.A(new_n709), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n490), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n713), .A2(KEYINPUT99), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(G8gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n715), .B(KEYINPUT100), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n717), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(new_n714), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n722), .B2(new_n714), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n720), .B1(new_n724), .B2(new_n725), .ZN(G1325gat));
  NAND2_X1  g525(.A1(new_n368), .A2(new_n371), .ZN(new_n727));
  OAI21_X1  g526(.A(G15gat), .B1(new_n709), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n366), .A2(G15gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n709), .B2(new_n729), .ZN(G1326gat));
  NOR2_X1   g529(.A1(new_n709), .A2(new_n455), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT43), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G22gat), .ZN(G1327gat));
  INV_X1    g538(.A(new_n640), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n705), .A2(KEYINPUT98), .A3(new_n692), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n741), .A2(new_n742), .B1(new_n687), .B2(new_n693), .ZN(new_n743));
  INV_X1    g542(.A(new_n676), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n740), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(G29gat), .A3(new_n539), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n600), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n751), .A2(new_n250), .A3(new_n707), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n583), .A2(new_n599), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n740), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT44), .B(new_n640), .C1(new_n583), .C2(new_n599), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT104), .B(new_n752), .C1(new_n755), .C2(new_n756), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n597), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G29gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n762), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n748), .B1(new_n764), .B2(new_n765), .ZN(G1328gat));
  NAND3_X1  g565(.A1(new_n759), .A2(new_n490), .A3(new_n760), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G36gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n745), .A2(G36gat), .A3(new_n491), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n600), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT46), .Z(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1329gat));
  OAI21_X1  g571(.A(G43gat), .B1(new_n757), .B2(new_n727), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n745), .A2(G43gat), .A3(new_n366), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n600), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(KEYINPUT47), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n775), .ZN(new_n777));
  INV_X1    g576(.A(new_n727), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n759), .A2(new_n778), .A3(new_n760), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(G43gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT107), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n784), .B(new_n776), .C1(new_n780), .C2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1330gat));
  OR3_X1    g585(.A1(new_n757), .A2(KEYINPUT108), .A3(new_n455), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT108), .B1(new_n757), .B2(new_n455), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(G50gat), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT48), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n745), .A2(G50gat), .A3(new_n455), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n600), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n790), .B1(new_n789), .B2(new_n793), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n456), .A3(new_n760), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n796), .A2(G50gat), .B1(new_n600), .B2(new_n792), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(KEYINPUT48), .B2(new_n797), .ZN(G1331gat));
  NOR3_X1   g597(.A1(new_n677), .A2(new_n743), .A3(new_n249), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT110), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n583), .B2(new_n599), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n597), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g602(.A(new_n491), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n805), .B(new_n806), .Z(G1333gat));
  INV_X1    g606(.A(G71gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n801), .A2(new_n808), .A3(new_n590), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n801), .A2(new_n778), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n808), .ZN(new_n811));
  XOR2_X1   g610(.A(new_n811), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g611(.A1(new_n801), .A2(new_n456), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g613(.A1(new_n744), .A2(new_n250), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT111), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n754), .A2(new_n740), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(KEYINPUT112), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n640), .B1(new_n583), .B2(new_n599), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(KEYINPUT51), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n824));
  INV_X1    g623(.A(new_n822), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n743), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n521), .A3(new_n597), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n820), .B(new_n753), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n817), .A2(new_n743), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n597), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n834), .B2(new_n521), .ZN(G1336gat));
  AOI21_X1  g634(.A(new_n475), .B1(new_n832), .B2(new_n490), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  INV_X1    g636(.A(new_n828), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n491), .A2(G92gat), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g640(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n825), .B2(new_n826), .ZN(new_n844));
  AOI211_X1 g643(.A(new_n743), .B(new_n840), .C1(new_n823), .C2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n845), .B2(new_n836), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n841), .A2(new_n846), .ZN(G1337gat));
  AOI21_X1  g646(.A(G99gat), .B1(new_n828), .B2(new_n590), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n832), .A2(G99gat), .A3(new_n778), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n848), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1338gat));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n743), .A2(G106gat), .A3(new_n455), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT115), .Z(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n823), .B2(new_n844), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n831), .B(new_n456), .C1(new_n755), .C2(new_n756), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G106gat), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT53), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n823), .B2(new_n827), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n855), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n862), .B(KEYINPUT116), .C1(new_n866), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1339gat));
  NOR3_X1   g669(.A1(new_n677), .A2(new_n707), .A3(new_n249), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n235), .A2(new_n237), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n228), .B1(new_n221), .B2(new_n227), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n244), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n248), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n637), .A2(new_n639), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n695), .A2(new_n879), .A3(new_n697), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n685), .A2(new_n686), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n685), .B2(new_n686), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n700), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n880), .A2(new_n883), .A3(KEYINPUT55), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n694), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT55), .B1(new_n880), .B2(new_n883), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n878), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT55), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n687), .A2(KEYINPUT54), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n685), .A2(new_n686), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n692), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n888), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(new_n249), .A3(new_n694), .A4(new_n884), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n743), .B2(new_n876), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n887), .B1(new_n895), .B2(new_n640), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n872), .B1(new_n896), .B2(new_n751), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n597), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n456), .A2(new_n595), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n898), .A2(new_n490), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(G113gat), .B1(new_n901), .B2(new_n249), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n539), .A2(new_n490), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n895), .A2(new_n640), .ZN(new_n906));
  INV_X1    g705(.A(new_n887), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n751), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n871), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n910), .B2(new_n456), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n897), .A2(KEYINPUT117), .A3(new_n455), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n366), .B(new_n904), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n250), .A2(new_n264), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n902), .B1(new_n913), .B2(new_n914), .ZN(G1340gat));
  AOI21_X1  g714(.A(G120gat), .B1(new_n901), .B2(new_n707), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n743), .A2(new_n265), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n913), .B2(new_n917), .ZN(G1341gat));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n255), .A3(new_n676), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n913), .A2(new_n751), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n255), .ZN(G1342gat));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n257), .A3(new_n740), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT56), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n257), .B1(new_n913), .B2(new_n740), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n923), .A2(new_n924), .ZN(G1343gat));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT58), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(KEYINPUT58), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n778), .A2(new_n904), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT118), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n896), .B2(new_n676), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n707), .A2(new_n877), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n740), .B1(new_n933), .B2(new_n894), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT118), .B(new_n744), .C1(new_n934), .C2(new_n887), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n935), .A3(new_n872), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n455), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n937), .B1(new_n910), .B2(new_n455), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n393), .B1(new_n941), .B2(new_n249), .ZN(new_n942));
  NOR4_X1   g741(.A1(new_n898), .A2(new_n490), .A3(new_n455), .A4(new_n778), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(new_n393), .A3(new_n249), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n927), .B(new_n928), .C1(new_n942), .C2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n938), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n744), .B1(new_n934), .B2(new_n887), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n871), .B1(new_n947), .B2(new_n931), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n935), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT57), .B1(new_n897), .B2(new_n456), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n249), .B(new_n929), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G141gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n943), .A2(new_n393), .A3(new_n249), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n952), .A2(new_n926), .A3(KEYINPUT58), .A4(new_n953), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n945), .A2(new_n954), .ZN(G1344gat));
  NAND2_X1  g754(.A1(new_n941), .A2(new_n707), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT59), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(G148gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n959));
  OAI21_X1  g758(.A(KEYINPUT57), .B1(new_n910), .B2(new_n455), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n947), .A2(new_n872), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n937), .A3(new_n456), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n960), .A2(new_n962), .A3(new_n707), .A4(new_n929), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G148gat), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n959), .B1(new_n964), .B2(KEYINPUT59), .ZN(new_n965));
  AOI211_X1 g764(.A(KEYINPUT120), .B(new_n957), .C1(new_n963), .C2(G148gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n943), .A2(new_n391), .A3(new_n707), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1345gat));
  NAND3_X1  g768(.A1(new_n943), .A2(new_n403), .A3(new_n676), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n941), .A2(new_n751), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n403), .ZN(G1346gat));
  NAND3_X1  g771(.A1(new_n943), .A2(new_n404), .A3(new_n740), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n941), .A2(new_n740), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n974), .B2(new_n404), .ZN(G1347gat));
  NAND2_X1  g774(.A1(new_n911), .A2(new_n912), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n597), .A2(new_n491), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(new_n590), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n980), .A2(new_n278), .A3(new_n250), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n897), .A2(new_n539), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT121), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n900), .A2(new_n491), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n983), .A2(KEYINPUT122), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT122), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n249), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n981), .B1(new_n987), .B2(new_n278), .ZN(G1348gat));
  OAI211_X1 g787(.A(new_n279), .B(new_n707), .C1(new_n985), .C2(new_n986), .ZN(new_n989));
  OAI21_X1  g788(.A(G176gat), .B1(new_n980), .B2(new_n743), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1349gat));
  OAI21_X1  g790(.A(G183gat), .B1(new_n980), .B2(new_n909), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n983), .A2(new_n296), .A3(new_n676), .A4(new_n984), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(KEYINPUT60), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT60), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n992), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1350gat));
  OAI211_X1 g797(.A(new_n293), .B(new_n740), .C1(new_n985), .C2(new_n986), .ZN(new_n999));
  XOR2_X1   g798(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n978), .B1(new_n911), .B2(new_n912), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1002), .A2(new_n740), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n1003), .B2(G190gat), .ZN(new_n1004));
  AOI211_X1 g803(.A(new_n293), .B(new_n1000), .C1(new_n1002), .C2(new_n740), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n999), .B1(new_n1004), .B2(new_n1005), .ZN(G1351gat));
  NAND2_X1  g805(.A1(new_n960), .A2(new_n962), .ZN(new_n1007));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n960), .A2(new_n962), .A3(KEYINPUT125), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n727), .A2(new_n977), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1012), .A2(G197gat), .A3(new_n249), .ZN(new_n1013));
  NOR2_X1   g812(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n727), .A2(new_n490), .A3(new_n456), .ZN(new_n1015));
  XOR2_X1   g814(.A(new_n1015), .B(KEYINPUT124), .Z(new_n1016));
  AND2_X1   g815(.A1(new_n983), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(G197gat), .B1(new_n1017), .B2(new_n249), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1014), .A2(new_n1018), .ZN(G1352gat));
  NOR2_X1   g818(.A1(new_n743), .A2(G204gat), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g821(.A1(new_n1012), .A2(new_n707), .ZN(new_n1023));
  OAI21_X1  g822(.A(G204gat), .B1(new_n1011), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g823(.A(KEYINPUT62), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1017), .A2(new_n1025), .A3(new_n1020), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .ZN(G1353gat));
  INV_X1    g826(.A(G211gat), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1017), .A2(new_n1028), .A3(new_n676), .ZN(new_n1029));
  NAND4_X1  g828(.A1(new_n960), .A2(new_n962), .A3(new_n676), .A4(new_n1012), .ZN(new_n1030));
  AND3_X1   g829(.A1(new_n1030), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1031));
  AOI21_X1  g830(.A(KEYINPUT63), .B1(new_n1030), .B2(G211gat), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G1354gat));
  NAND3_X1  g832(.A1(new_n983), .A2(new_n740), .A3(new_n1016), .ZN(new_n1034));
  INV_X1    g833(.A(G218gat), .ZN(new_n1035));
  AND3_X1   g834(.A1(new_n1034), .A2(KEYINPUT126), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g835(.A(KEYINPUT126), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n640), .A2(new_n1035), .ZN(new_n1038));
  XNOR2_X1  g837(.A(new_n1038), .B(KEYINPUT127), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1039), .A2(new_n1012), .ZN(new_n1040));
  AOI21_X1  g839(.A(new_n1040), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1041));
  NOR3_X1   g840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(G1355gat));
endmodule


