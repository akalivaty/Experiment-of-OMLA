

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n472), .B(n471), .ZN(n571) );
  XNOR2_X1 U325 ( .A(n447), .B(n446), .ZN(n576) );
  XOR2_X1 U326 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n292) );
  AND2_X1 U327 ( .A1(G228GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U328 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n294) );
  XNOR2_X1 U329 ( .A(n373), .B(n293), .ZN(n374) );
  XNOR2_X1 U330 ( .A(n375), .B(n374), .ZN(n376) );
  INV_X1 U331 ( .A(KEYINPUT22), .ZN(n381) );
  XNOR2_X1 U332 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U333 ( .A(n384), .B(n383), .ZN(n388) );
  INV_X1 U334 ( .A(KEYINPUT66), .ZN(n471) );
  NOR2_X1 U335 ( .A1(n412), .A2(n411), .ZN(n480) );
  XNOR2_X1 U336 ( .A(n405), .B(KEYINPUT26), .ZN(n570) );
  NOR2_X1 U337 ( .A1(n533), .A2(n564), .ZN(n477) );
  XNOR2_X1 U338 ( .A(KEYINPUT38), .B(n448), .ZN(n495) );
  XNOR2_X1 U339 ( .A(n449), .B(G29GAT), .ZN(n450) );
  XNOR2_X1 U340 ( .A(n451), .B(n450), .ZN(G1328GAT) );
  XOR2_X1 U341 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n419) );
  XOR2_X1 U344 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n298) );
  XNOR2_X1 U345 ( .A(G218GAT), .B(KEYINPUT67), .ZN(n297) );
  XOR2_X1 U346 ( .A(n298), .B(n297), .Z(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n300) );
  XNOR2_X1 U348 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U351 ( .A(G106GAT), .B(G92GAT), .Z(n304) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U354 ( .A(KEYINPUT11), .B(n305), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n309) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G85GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n308), .B(KEYINPUT76), .ZN(n445) );
  XNOR2_X1 U358 ( .A(n309), .B(n445), .ZN(n311) );
  XOR2_X1 U359 ( .A(G134GAT), .B(KEYINPUT81), .Z(n341) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XOR2_X1 U361 ( .A(n341), .B(n373), .Z(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n419), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(G36GAT), .B(G190GAT), .Z(n313) );
  XOR2_X1 U365 ( .A(KEYINPUT82), .B(n313), .Z(n395) );
  XNOR2_X1 U366 ( .A(n314), .B(n395), .ZN(n552) );
  INV_X1 U367 ( .A(n552), .ZN(n455) );
  XNOR2_X1 U368 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n455), .B(n315), .ZN(n585) );
  XOR2_X1 U370 ( .A(G78GAT), .B(G64GAT), .Z(n317) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G183GAT), .ZN(n316) );
  XNOR2_X1 U372 ( .A(n317), .B(n316), .ZN(n331) );
  XOR2_X1 U373 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n319) );
  XNOR2_X1 U374 ( .A(KEYINPUT14), .B(KEYINPUT83), .ZN(n318) );
  XNOR2_X1 U375 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G155GAT), .Z(n380) );
  XOR2_X1 U377 ( .A(n380), .B(G211GAT), .Z(n321) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G127GAT), .Z(n364) );
  XNOR2_X1 U379 ( .A(n364), .B(G8GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n325) );
  AND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U384 ( .A(n326), .B(KEYINPUT15), .Z(n329) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n294), .B(n327), .ZN(n437) );
  XNOR2_X1 U387 ( .A(n437), .B(KEYINPUT12), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n580) );
  INV_X1 U390 ( .A(n580), .ZN(n533) );
  XOR2_X1 U391 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n333) );
  XNOR2_X1 U392 ( .A(KEYINPUT4), .B(KEYINPUT5), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n352) );
  XOR2_X1 U394 ( .A(G155GAT), .B(G148GAT), .Z(n335) );
  XNOR2_X1 U395 ( .A(G1GAT), .B(G127GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U397 ( .A(G57GAT), .B(G85GAT), .Z(n337) );
  XNOR2_X1 U398 ( .A(G29GAT), .B(G162GAT), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U400 ( .A(n339), .B(n338), .ZN(n350) );
  XNOR2_X1 U401 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n292), .B(n340), .ZN(n375) );
  XOR2_X1 U403 ( .A(n375), .B(n341), .Z(n343) );
  NAND2_X1 U404 ( .A1(G225GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U405 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U406 ( .A(n344), .B(KEYINPUT93), .Z(n348) );
  XOR2_X1 U407 ( .A(KEYINPUT86), .B(KEYINPUT0), .Z(n346) );
  XNOR2_X1 U408 ( .A(G113GAT), .B(G120GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n346), .B(n345), .ZN(n365) );
  XNOR2_X1 U410 ( .A(n365), .B(KEYINPUT94), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n523) );
  INV_X1 U414 ( .A(n523), .ZN(n401) );
  XOR2_X1 U415 ( .A(KEYINPUT18), .B(KEYINPUT89), .Z(n354) );
  XNOR2_X1 U416 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U418 ( .A(KEYINPUT19), .B(n355), .Z(n396) );
  XOR2_X1 U419 ( .A(G99GAT), .B(G190GAT), .Z(n357) );
  XNOR2_X1 U420 ( .A(G43GAT), .B(G134GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U422 ( .A(KEYINPUT87), .B(G71GAT), .Z(n359) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G176GAT), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U425 ( .A(n361), .B(n360), .Z(n371) );
  XOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT90), .Z(n363) );
  XNOR2_X1 U427 ( .A(KEYINPUT20), .B(KEYINPUT88), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n369) );
  XOR2_X1 U429 ( .A(n365), .B(n364), .Z(n367) );
  NAND2_X1 U430 ( .A1(G227GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n396), .B(n372), .ZN(n515) );
  XOR2_X1 U435 ( .A(n376), .B(KEYINPUT24), .Z(n379) );
  XNOR2_X1 U436 ( .A(G148GAT), .B(G106GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n377), .B(G78GAT), .ZN(n436) );
  XNOR2_X1 U438 ( .A(n436), .B(KEYINPUT23), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n380), .B(G204GAT), .ZN(n382) );
  XOR2_X1 U441 ( .A(KEYINPUT21), .B(KEYINPUT91), .Z(n386) );
  XNOR2_X1 U442 ( .A(G218GAT), .B(G211GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(G197GAT), .B(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n388), .B(n389), .ZN(n473) );
  XOR2_X1 U446 ( .A(n473), .B(KEYINPUT28), .Z(n528) );
  XOR2_X1 U447 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XNOR2_X1 U448 ( .A(n389), .B(n418), .ZN(n391) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n394) );
  XOR2_X1 U451 ( .A(G204GAT), .B(G64GAT), .Z(n393) );
  XNOR2_X1 U452 ( .A(G176GAT), .B(G92GAT), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n444) );
  XOR2_X1 U454 ( .A(n394), .B(n444), .Z(n398) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n513) );
  XOR2_X1 U457 ( .A(n513), .B(KEYINPUT27), .Z(n406) );
  INV_X1 U458 ( .A(n406), .ZN(n522) );
  NAND2_X1 U459 ( .A1(n528), .A2(n522), .ZN(n399) );
  NOR2_X1 U460 ( .A1(n515), .A2(n399), .ZN(n400) );
  NOR2_X1 U461 ( .A1(n401), .A2(n400), .ZN(n412) );
  AND2_X1 U462 ( .A1(n515), .A2(n513), .ZN(n402) );
  NOR2_X1 U463 ( .A1(n473), .A2(n402), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT25), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n404), .B(KEYINPUT95), .ZN(n408) );
  INV_X1 U466 ( .A(n515), .ZN(n526) );
  NAND2_X1 U467 ( .A1(n473), .A2(n526), .ZN(n405) );
  NOR2_X1 U468 ( .A1(n570), .A2(n406), .ZN(n407) );
  NOR2_X1 U469 ( .A1(n408), .A2(n407), .ZN(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT96), .B(n409), .Z(n410) );
  NOR2_X1 U471 ( .A1(n523), .A2(n410), .ZN(n411) );
  NAND2_X1 U472 ( .A1(n533), .A2(n480), .ZN(n413) );
  NOR2_X1 U473 ( .A1(n585), .A2(n413), .ZN(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT99), .B(KEYINPUT37), .Z(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n510) );
  XOR2_X1 U476 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n417) );
  XNOR2_X1 U477 ( .A(G197GAT), .B(G22GAT), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n432) );
  XOR2_X1 U479 ( .A(n418), .B(G36GAT), .Z(n421) );
  XNOR2_X1 U480 ( .A(n419), .B(G50GAT), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U482 ( .A(G141GAT), .B(G1GAT), .Z(n423) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U485 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U486 ( .A(G113GAT), .B(KEYINPUT30), .Z(n427) );
  XNOR2_X1 U487 ( .A(KEYINPUT70), .B(KEYINPUT29), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n428), .B(G15GAT), .ZN(n429) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n554) );
  INV_X1 U492 ( .A(n554), .ZN(n572) );
  XOR2_X1 U493 ( .A(KEYINPUT74), .B(KEYINPUT77), .Z(n434) );
  NAND2_X1 U494 ( .A1(G230GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(KEYINPUT75), .Z(n439) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n443) );
  XOR2_X1 U499 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n441) );
  XNOR2_X1 U500 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U504 ( .A1(n572), .A2(n576), .ZN(n482) );
  NOR2_X1 U505 ( .A1(n510), .A2(n482), .ZN(n448) );
  NAND2_X1 U506 ( .A1(n495), .A2(n523), .ZN(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n449) );
  INV_X1 U508 ( .A(KEYINPUT54), .ZN(n469) );
  XOR2_X1 U509 ( .A(KEYINPUT107), .B(KEYINPUT47), .Z(n458) );
  XNOR2_X1 U510 ( .A(n576), .B(KEYINPUT65), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(KEYINPUT41), .ZN(n558) );
  NOR2_X1 U512 ( .A1(n558), .A2(n554), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(KEYINPUT46), .ZN(n454) );
  NOR2_X1 U514 ( .A1(n454), .A2(n580), .ZN(n456) );
  NAND2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n533), .A2(n585), .ZN(n459) );
  XNOR2_X1 U518 ( .A(KEYINPUT45), .B(n459), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n460), .A2(n576), .ZN(n461) );
  NOR2_X1 U520 ( .A1(n572), .A2(n461), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n466) );
  XNOR2_X1 U522 ( .A(KEYINPUT48), .B(KEYINPUT108), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT64), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n521) );
  XOR2_X1 U525 ( .A(KEYINPUT116), .B(n513), .Z(n467) );
  NOR2_X1 U526 ( .A1(n521), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n470), .A2(n523), .ZN(n472) );
  NOR2_X1 U529 ( .A1(n571), .A2(n473), .ZN(n475) );
  XNOR2_X1 U530 ( .A(KEYINPUT117), .B(KEYINPUT55), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n476), .A2(n515), .ZN(n564) );
  XNOR2_X1 U533 ( .A(KEYINPUT122), .B(n477), .ZN(n478) );
  XOR2_X1 U534 ( .A(G183GAT), .B(n478), .Z(G1350GAT) );
  NOR2_X1 U535 ( .A1(n552), .A2(n533), .ZN(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT16), .B(n479), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n481), .A2(n480), .ZN(n500) );
  NOR2_X1 U538 ( .A1(n482), .A2(n500), .ZN(n483) );
  XOR2_X1 U539 ( .A(KEYINPUT97), .B(n483), .Z(n489) );
  NAND2_X1 U540 ( .A1(n523), .A2(n489), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n489), .A2(n513), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U546 ( .A1(n489), .A2(n515), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(G1326GAT) );
  INV_X1 U548 ( .A(n528), .ZN(n518) );
  NAND2_X1 U549 ( .A1(n518), .A2(n489), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n495), .A2(n513), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n491), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U554 ( .A1(n495), .A2(n515), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(KEYINPUT102), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n518), .A2(n495), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(KEYINPUT103), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n499), .Z(n502) );
  INV_X1 U563 ( .A(n558), .ZN(n544) );
  NAND2_X1 U564 ( .A1(n554), .A2(n544), .ZN(n509) );
  NOR2_X1 U565 ( .A1(n500), .A2(n509), .ZN(n505) );
  NAND2_X1 U566 ( .A1(n505), .A2(n523), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n505), .A2(n513), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U570 ( .A1(n515), .A2(n505), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U573 ( .A1(n505), .A2(n518), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n508), .Z(G1335GAT) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n512) );
  NOR2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n517), .A2(n523), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n513), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n515), .A2(n517), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U588 ( .A1(n521), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT109), .B(n525), .ZN(n541) );
  NOR2_X1 U590 ( .A1(n541), .A2(n526), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(KEYINPUT110), .B(n529), .ZN(n537) );
  NOR2_X1 U593 ( .A1(n537), .A2(n554), .ZN(n530) );
  XOR2_X1 U594 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  XNOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n558), .A2(n537), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT111), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n533), .A2(n537), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n537), .A2(n455), .ZN(n539) );
  XNOR2_X1 U603 ( .A(KEYINPUT51), .B(KEYINPUT112), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n570), .A2(n541), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(n542), .Z(n551) );
  NAND2_X1 U608 ( .A1(n572), .A2(n551), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XNOR2_X1 U610 ( .A(KEYINPUT114), .B(KEYINPUT52), .ZN(n548) );
  XOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .Z(n546) );
  NAND2_X1 U612 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  XOR2_X1 U615 ( .A(G155GAT), .B(KEYINPUT115), .Z(n550) );
  NAND2_X1 U616 ( .A1(n551), .A2(n580), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n553), .ZN(G1347GAT) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n557) );
  NOR2_X1 U621 ( .A1(n564), .A2(n554), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(KEYINPUT119), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n564), .ZN(n563) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(KEYINPUT56), .B(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n455), .ZN(n566) );
  XNOR2_X1 U631 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n575) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(n573), .Z(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n578) );
  INV_X1 U642 ( .A(n581), .ZN(n584) );
  OR2_X1 U643 ( .A1(n584), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT127), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

