//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT2), .A2(G113), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n190), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT2), .A2(G113), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(KEYINPUT67), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n194), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n192), .B(KEYINPUT67), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n196), .A2(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n189), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n216), .A3(G101), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n204), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n208), .A2(G104), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n205), .A2(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(G101), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n214), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G113), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n197), .A2(G119), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT5), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n196), .A2(new_n198), .A3(KEYINPUT5), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n226), .A2(KEYINPUT80), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT80), .B1(new_n226), .B2(new_n227), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n222), .B(new_n203), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n188), .B1(new_n218), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n231), .A2(KEYINPUT6), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n230), .A3(new_n188), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT81), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n218), .A2(new_n230), .A3(new_n235), .A4(new_n188), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n231), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT6), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(G128), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n241), .B(new_n243), .C1(KEYINPUT1), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G125), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(KEYINPUT82), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT82), .B1(new_n249), .B2(new_n250), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n241), .A2(new_n243), .A3(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT0), .B(G128), .Z(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI22_X1  g071(.A1(new_n251), .A2(new_n252), .B1(new_n250), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n259));
  INV_X1    g073(.A(G224), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G953), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(KEYINPUT84), .A3(G224), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n264), .B(KEYINPUT83), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n258), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n214), .A2(new_n221), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n226), .A2(new_n227), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n203), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n188), .B(KEYINPUT8), .Z(new_n271));
  NOR2_X1   g085(.A1(new_n228), .A2(new_n229), .ZN(new_n272));
  INV_X1    g086(.A(new_n203), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n270), .B(new_n271), .C1(new_n274), .C2(new_n268), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n263), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n258), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n258), .A2(new_n277), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n275), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n234), .A2(new_n236), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(G210), .B1(G237), .B2(G902), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n267), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n285), .B1(new_n267), .B2(new_n282), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n187), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  XNOR2_X1  g105(.A(G110), .B(G140), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n262), .A2(G227), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g108(.A(KEYINPUT65), .ZN(new_n295));
  INV_X1    g109(.A(G137), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(G134), .ZN(new_n297));
  INV_X1    g111(.A(G134), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT65), .A3(G137), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n296), .A2(KEYINPUT11), .A3(G134), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT11), .B1(new_n296), .B2(G134), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G131), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT11), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n298), .B2(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(KEYINPUT11), .A3(G134), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n297), .A2(new_n307), .A3(new_n299), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT79), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n312), .A2(new_n215), .A3(new_n257), .A4(new_n217), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n217), .A2(new_n257), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n314), .B2(new_n215), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n249), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT10), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n268), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n246), .A2(new_n320), .A3(new_n248), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n249), .A2(new_n268), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(KEYINPUT10), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n311), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n215), .A2(new_n257), .A3(new_n217), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT79), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n312), .A3(new_n215), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n246), .A2(new_n320), .A3(new_n248), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n320), .B1(new_n246), .B2(new_n248), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n222), .A2(new_n248), .A3(new_n246), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n332), .A2(new_n319), .B1(new_n333), .B2(new_n318), .ZN(new_n334));
  INV_X1    g148(.A(new_n311), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n294), .B1(new_n325), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n246), .A2(new_n248), .B1(new_n214), .B2(new_n221), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n311), .B1(new_n323), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT12), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(KEYINPUT12), .B(new_n311), .C1(new_n323), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n336), .A2(new_n343), .A3(new_n294), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n290), .B(new_n291), .C1(new_n337), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(G469), .A2(G902), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n336), .A2(new_n343), .ZN(new_n347));
  INV_X1    g161(.A(new_n294), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n325), .A2(new_n336), .A3(new_n294), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(G469), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G475), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n250), .A2(G140), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(new_n354), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n240), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n250), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  XNOR2_X1  g176(.A(G125), .B(G140), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n363), .B2(KEYINPUT16), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G146), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n369));
  AOI21_X1  g183(.A(G143), .B1(new_n368), .B2(G214), .ZN(new_n370));
  OAI21_X1  g184(.A(G131), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT17), .ZN(new_n373));
  OR3_X1    g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n242), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n304), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n378), .A3(new_n373), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n372), .B1(new_n371), .B2(new_n373), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n367), .A2(new_n374), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n369), .A2(new_n370), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT18), .A2(G131), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n359), .A2(G146), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n363), .A2(new_n240), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n382), .A2(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT18), .B(G131), .C1(new_n369), .C2(new_n370), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(new_n377), .A3(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT86), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(G113), .B(G122), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(new_n205), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n381), .A2(new_n394), .A3(new_n397), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n353), .B1(new_n401), .B2(new_n291), .ZN(new_n402));
  NOR2_X1   g216(.A1(G475), .A2(G902), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n371), .A2(new_n378), .B1(new_n364), .B2(G146), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT19), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT19), .B1(new_n357), .B2(new_n358), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n240), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT87), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT19), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n359), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n363), .A2(KEYINPUT19), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT87), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(new_n240), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n404), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n387), .B1(new_n386), .B2(new_n388), .ZN(new_n416));
  AND4_X1   g230(.A1(new_n387), .A2(new_n388), .A3(new_n390), .A4(new_n391), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(new_n398), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n400), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n418), .B2(new_n398), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n403), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n398), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT88), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n420), .A3(new_n400), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n403), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n402), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT9), .B(G234), .ZN(new_n431));
  OAI21_X1  g245(.A(G221), .B1(new_n431), .B2(G902), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT77), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT78), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G116), .B(G122), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(new_n208), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n247), .A2(G143), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n247), .A2(G143), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n298), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n438), .B1(KEYINPUT13), .B2(new_n440), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n438), .A2(KEYINPUT13), .ZN(new_n444));
  OAI21_X1  g258(.A(G134), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n437), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G217), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n431), .A2(new_n447), .A3(G953), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n197), .A2(G122), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n197), .A2(G122), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n452), .B2(KEYINPUT90), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(KEYINPUT90), .B2(new_n452), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n454), .A2(G107), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n436), .A2(new_n208), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n298), .B1(new_n439), .B2(new_n440), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n441), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n446), .B(new_n448), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n448), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n454), .B2(G107), .ZN(new_n461));
  INV_X1    g275(.A(new_n446), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n291), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT15), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(G478), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n464), .B(new_n291), .C1(KEYINPUT15), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n262), .A2(G952), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(G234), .B2(G237), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n291), .B(new_n262), .C1(G234), .C2(G237), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT21), .B(G898), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n352), .A2(new_n430), .A3(new_n435), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n289), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n368), .A2(G210), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(KEYINPUT27), .Z(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT26), .B(G101), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n480), .B(new_n481), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT71), .B(KEYINPUT28), .ZN(new_n484));
  INV_X1    g298(.A(new_n204), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n298), .A2(G137), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n296), .A2(G134), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n304), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n309), .B2(G131), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n249), .ZN(new_n491));
  OR2_X1    g305(.A1(KEYINPUT0), .A2(G128), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n241), .A2(new_n243), .B1(new_n492), .B2(new_n253), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n241), .A2(new_n243), .A3(new_n253), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT64), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n495), .A2(new_n497), .B1(new_n305), .B2(new_n310), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT66), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n491), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n495), .A2(new_n497), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n311), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT66), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n485), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AND4_X1   g318(.A1(new_n297), .A2(new_n307), .A3(new_n299), .A4(new_n308), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n488), .B1(new_n505), .B2(new_n304), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n317), .A2(new_n506), .A3(new_n321), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n311), .A2(new_n257), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n204), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n200), .A2(new_n203), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT72), .B(new_n484), .C1(new_n504), .C2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n501), .A2(new_n311), .A3(new_n499), .ZN(new_n518));
  INV_X1    g332(.A(new_n491), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n498), .A2(new_n499), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n204), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n512), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT72), .B1(new_n523), .B2(new_n484), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n483), .B1(new_n517), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n520), .B2(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n507), .A2(new_n508), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n526), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT69), .A4(KEYINPUT30), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(new_n530), .A3(new_n204), .A4(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n482), .A3(new_n512), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n532), .A2(new_n535), .A3(new_n482), .A4(new_n512), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(KEYINPUT32), .A3(new_n538), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n511), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n513), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n516), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT29), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n483), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(G902), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n517), .A2(new_n524), .A3(new_n483), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n532), .A2(new_n512), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n483), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(G472), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n541), .A2(new_n542), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G234), .ZN(new_n558));
  OAI21_X1  g372(.A(G217), .B1(new_n558), .B2(G902), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT73), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OR3_X1    g375(.A1(new_n247), .A2(KEYINPUT74), .A3(G119), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n195), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT74), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n562), .A2(new_n564), .B1(G119), .B2(new_n247), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n247), .A2(G119), .ZN(new_n568));
  OR2_X1    g382(.A1(new_n568), .A2(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n563), .A3(KEYINPUT23), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(G110), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n366), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n565), .A2(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(G110), .B1(new_n569), .B2(new_n570), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n365), .B(new_n385), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n581), .B(new_n580), .C1(new_n572), .C2(new_n575), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n561), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n582), .A2(new_n580), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n581), .B1(new_n572), .B2(new_n575), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n291), .B1(new_n591), .B2(new_n584), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n583), .A2(new_n585), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n559), .A2(new_n291), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n588), .A2(new_n593), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n557), .A2(KEYINPUT76), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT76), .B1(new_n557), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n478), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n352), .A2(new_n435), .ZN(new_n602));
  INV_X1    g416(.A(new_n597), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n537), .A2(new_n291), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT91), .B1(new_n605), .B2(G472), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT91), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n607), .B(new_n608), .C1(new_n537), .C2(new_n291), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n539), .B(new_n604), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n402), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n423), .A2(KEYINPUT20), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n428), .B1(new_n427), .B2(new_n403), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT92), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n468), .A2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n459), .A2(new_n463), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n459), .B2(new_n463), .ZN(new_n620));
  OAI211_X1 g434(.A(new_n615), .B(new_n616), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n616), .ZN(new_n622));
  INV_X1    g436(.A(new_n620), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n622), .B1(new_n623), .B2(new_n618), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT92), .B1(new_n465), .B2(new_n468), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n267), .A2(new_n282), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n283), .ZN(new_n629));
  INV_X1    g443(.A(new_n475), .ZN(new_n630));
  INV_X1    g444(.A(new_n283), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n267), .A2(new_n282), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n629), .A2(new_n187), .A3(new_n630), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n610), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  NAND3_X1  g450(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT93), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n423), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n611), .A4(new_n470), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n610), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT94), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT35), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G9));
  NOR2_X1   g457(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n576), .B(new_n644), .Z(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(new_n595), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n588), .B2(new_n593), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n289), .A2(new_n477), .A3(new_n647), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n648), .B(new_n539), .C1(new_n606), .C2(new_n609), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  NAND2_X1  g465(.A1(new_n629), .A2(new_n632), .ZN(new_n652));
  INV_X1    g466(.A(new_n187), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n653), .A3(new_n647), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n557), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n473), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n472), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n639), .A2(new_n602), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NAND2_X1  g477(.A1(new_n628), .A2(new_n284), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n286), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n647), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n470), .A2(new_n187), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n430), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n483), .B1(new_n513), .B2(new_n543), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n533), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n674), .B2(G902), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n541), .A2(new_n542), .A3(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n672), .A2(KEYINPUT96), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT96), .B1(new_n672), .B2(new_n676), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n659), .B(KEYINPUT39), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n352), .A2(new_n435), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT40), .ZN(new_n681));
  OR3_X1    g495(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NAND3_X1  g497(.A1(new_n614), .A2(new_n626), .A3(new_n659), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n602), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n655), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NOR2_X1   g501(.A1(new_n633), .A2(new_n627), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n291), .B1(new_n337), .B2(new_n344), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n691), .A3(new_n345), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n689), .A2(KEYINPUT97), .A3(G469), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n433), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n557), .A2(new_n597), .A3(new_n688), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NOR2_X1   g511(.A1(new_n633), .A2(new_n639), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n557), .A2(new_n597), .A3(new_n698), .A4(new_n694), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NAND2_X1  g514(.A1(new_n430), .A2(new_n476), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n557), .A2(new_n702), .A3(new_n654), .A4(new_n694), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  INV_X1    g518(.A(new_n538), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n533), .A2(KEYINPUT31), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n482), .B1(new_n544), .B2(new_n516), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT98), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n536), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n707), .B1(new_n533), .B2(KEYINPUT31), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT98), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n705), .B1(new_n708), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n608), .B1(new_n537), .B2(new_n291), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n603), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n671), .A2(new_n652), .A3(new_n475), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n694), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AND3_X1   g532(.A1(new_n629), .A2(new_n187), .A3(new_n632), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n614), .A2(new_n626), .A3(new_n659), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n694), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n713), .A2(new_n714), .A3(new_n647), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT102), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n352), .A2(KEYINPUT99), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n345), .A2(new_n728), .A3(new_n346), .A4(new_n351), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n433), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n664), .A2(new_n187), .A3(new_n286), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n557), .A2(new_n597), .A3(new_n733), .A4(new_n720), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n542), .A2(KEYINPUT100), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT100), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n537), .A2(new_n737), .A3(KEYINPUT32), .A4(new_n538), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n541), .A3(new_n556), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n597), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n730), .A2(new_n732), .A3(new_n684), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT42), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n735), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NOR4_X1   g557(.A1(new_n730), .A2(new_n732), .A3(new_n684), .A4(new_n726), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT101), .A3(new_n739), .A4(new_n597), .ZN(new_n745));
  AOI221_X4 g559(.A(new_n725), .B1(new_n726), .B2(new_n734), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n734), .A2(new_n726), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT102), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT103), .B(G131), .Z(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G33));
  NOR2_X1   g566(.A1(new_n639), .A2(new_n660), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n557), .A2(new_n597), .A3(new_n733), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  OAI21_X1  g569(.A(new_n539), .B1(new_n606), .B2(new_n609), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n668), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT105), .A3(new_n668), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n430), .A2(new_n626), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT43), .Z(new_n762));
  NAND3_X1  g576(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n664), .A2(new_n187), .A3(new_n286), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n763), .A2(new_n764), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n351), .B1(new_n769), .B2(new_n290), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n349), .A2(KEYINPUT45), .A3(new_n350), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n346), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n345), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT46), .B1(new_n775), .B2(new_n346), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n731), .B(new_n679), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n765), .A2(new_n767), .A3(new_n768), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  OAI21_X1  g596(.A(new_n731), .B1(new_n777), .B2(new_n778), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n557), .A2(new_n597), .A3(new_n684), .A4(new_n766), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  OR2_X1    g602(.A1(new_n676), .A2(new_n603), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n692), .A2(new_n693), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT49), .Z(new_n791));
  INV_X1    g605(.A(new_n667), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n430), .A2(new_n187), .A3(new_n435), .A4(new_n626), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n789), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT106), .Z(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n557), .B(new_n654), .C1(new_n661), .C2(new_n685), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n731), .A2(new_n659), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n646), .B(new_n798), .C1(new_n588), .C2(new_n593), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n670), .A2(new_n799), .A3(new_n629), .A4(new_n632), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n730), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n676), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n797), .A2(new_n723), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n797), .A2(new_n723), .A3(new_n802), .A4(KEYINPUT52), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n695), .A2(new_n699), .ZN(new_n808));
  INV_X1    g622(.A(new_n470), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n627), .B1(new_n614), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n665), .A3(new_n187), .A4(new_n630), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n610), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n649), .A2(new_n717), .A3(new_n703), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n722), .A2(new_n741), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n470), .A2(new_n402), .A3(new_n660), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n638), .A3(new_n637), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT107), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT107), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n816), .A2(new_n819), .A3(new_n638), .A4(new_n637), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n766), .A2(new_n602), .A3(new_n647), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n557), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n754), .A2(new_n815), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n813), .A2(new_n600), .A3(new_n814), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n807), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n750), .A2(new_n826), .A3(KEYINPUT53), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT53), .B1(new_n750), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(KEYINPUT108), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n747), .A2(new_n748), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n725), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n747), .A2(KEYINPUT102), .A3(new_n748), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n814), .A2(new_n600), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n805), .A2(new_n806), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n813), .A4(new_n824), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT108), .B(new_n830), .C1(new_n834), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n796), .B(KEYINPUT54), .C1(new_n829), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n830), .B1(new_n834), .B2(new_n837), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT110), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n828), .A2(KEYINPUT110), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n831), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT108), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n838), .A3(new_n827), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n796), .B1(new_n851), .B2(KEYINPUT54), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n790), .A2(new_n434), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n784), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n762), .A2(new_n472), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(new_n715), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n766), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n667), .A2(new_n653), .A3(new_n694), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n857), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n857), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n767), .A2(new_n731), .A3(new_n790), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n789), .A2(new_n658), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n614), .A2(new_n626), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n855), .A2(new_n865), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n866), .A2(new_n867), .B1(new_n722), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(KEYINPUT112), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n864), .B2(new_n869), .ZN(new_n873));
  OAI211_X1 g687(.A(KEYINPUT51), .B(new_n859), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n471), .B(KEYINPUT113), .ZN(new_n875));
  INV_X1    g689(.A(new_n857), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n694), .A2(new_n719), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n866), .A2(new_n614), .A3(new_n626), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n868), .A2(new_n597), .A3(new_n739), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n878), .B(new_n879), .C1(new_n881), .C2(KEYINPUT48), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n883), .A2(KEYINPUT48), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n882), .B1(new_n884), .B2(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n859), .A2(KEYINPUT111), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT111), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n854), .A2(new_n887), .A3(new_n858), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n870), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n874), .B(new_n885), .C1(new_n889), .C2(KEYINPUT51), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n848), .A2(new_n852), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n795), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT115), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT115), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n795), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(G75));
  NAND3_X1  g711(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(G210), .A3(G902), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n239), .B(new_n266), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n899), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n899), .B2(new_n900), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n262), .A2(G952), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT116), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(G51));
  NAND2_X1  g722(.A1(new_n898), .A2(G902), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n775), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT117), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n346), .B(KEYINPUT57), .Z(new_n912));
  AND2_X1   g726(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n913));
  INV_X1    g727(.A(new_n847), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n337), .B2(new_n344), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n905), .B1(new_n911), .B2(new_n916), .ZN(G54));
  NAND4_X1  g731(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n918));
  INV_X1    g732(.A(new_n427), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n905), .ZN(G60));
  OR2_X1    g736(.A1(new_n913), .A2(new_n914), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n619), .A2(new_n620), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n907), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n848), .A2(new_n852), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n926), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  XNOR2_X1  g745(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n447), .A2(new_n291), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n898), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n585), .A3(new_n583), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n645), .B(KEYINPUT119), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n936), .B(new_n906), .C1(new_n935), .C2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  NOR3_X1   g754(.A1(new_n474), .A2(new_n260), .A3(new_n262), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n835), .A2(new_n813), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n262), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT120), .ZN(new_n944));
  INV_X1    g758(.A(new_n239), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(G898), .B2(new_n262), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  AOI21_X1  g761(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n527), .A2(new_n531), .A3(new_n530), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n412), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n797), .A2(new_n723), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n682), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n682), .A2(KEYINPUT62), .A3(new_n953), .ZN(new_n957));
  AOI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(new_n785), .B2(new_n786), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n766), .A2(new_n680), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n810), .B(new_n959), .C1(new_n598), .C2(new_n599), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n781), .A2(KEYINPUT121), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT121), .B1(new_n781), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n952), .B1(new_n963), .B2(new_n262), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI211_X1 g780(.A(KEYINPUT122), .B(new_n952), .C1(new_n963), .C2(new_n262), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n949), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OR4_X1    g782(.A1(new_n652), .A2(new_n779), .A3(new_n671), .A4(new_n740), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n750), .A2(new_n787), .A3(new_n754), .A4(new_n969), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n781), .A2(KEYINPUT124), .A3(new_n953), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT124), .B1(new_n781), .B2(new_n953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n970), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(KEYINPUT125), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT125), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n970), .B(new_n975), .C1(new_n971), .C2(new_n972), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n262), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n951), .B1(G900), .B2(G953), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n948), .B1(new_n968), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n964), .B(new_n965), .ZN(new_n982));
  INV_X1    g796(.A(new_n948), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n982), .A2(new_n949), .A3(new_n983), .A4(new_n979), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(G72));
  XNOR2_X1  g799(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n608), .A2(new_n291), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n986), .B(new_n987), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n553), .B2(new_n533), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n905), .B1(new_n851), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n552), .A2(new_n482), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n958), .B(new_n942), .C1(new_n962), .C2(new_n961), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n992), .B1(new_n993), .B2(new_n988), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n974), .A2(new_n942), .A3(new_n976), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n482), .B(new_n552), .C1(new_n999), .C2(new_n988), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(G57));
endmodule


