

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  OR2_X1 U324 ( .A1(n451), .A2(n538), .ZN(n573) );
  XNOR2_X2 U325 ( .A(n346), .B(n293), .ZN(n584) );
  NOR2_X1 U326 ( .A1(n537), .A2(n530), .ZN(n393) );
  XOR2_X1 U327 ( .A(G71GAT), .B(KEYINPUT13), .Z(n350) );
  OR2_X1 U328 ( .A1(n562), .A2(n538), .ZN(n292) );
  XNOR2_X1 U329 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n368) );
  XNOR2_X1 U330 ( .A(n329), .B(n400), .ZN(n331) );
  XNOR2_X1 U331 ( .A(n376), .B(n375), .ZN(n537) );
  XNOR2_X1 U332 ( .A(KEYINPUT111), .B(KEYINPUT48), .ZN(n375) );
  XOR2_X1 U333 ( .A(n363), .B(n362), .Z(n565) );
  XNOR2_X1 U334 ( .A(n584), .B(KEYINPUT41), .ZN(n562) );
  XOR2_X1 U335 ( .A(n345), .B(n344), .Z(n293) );
  AND2_X1 U336 ( .A1(G231GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n330) );
  XNOR2_X1 U338 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U339 ( .A(n355), .B(n294), .ZN(n356) );
  XOR2_X1 U340 ( .A(G1GAT), .B(G127GAT), .Z(n408) );
  XNOR2_X1 U341 ( .A(n357), .B(n356), .ZN(n358) );
  INV_X1 U342 ( .A(G218GAT), .ZN(n467) );
  INV_X1 U343 ( .A(n573), .ZN(n570) );
  XNOR2_X1 U344 ( .A(n467), .B(KEYINPUT62), .ZN(n468) );
  XNOR2_X1 U345 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U346 ( .A(n469), .B(n468), .ZN(G1355GAT) );
  XNOR2_X1 U347 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT11), .B(KEYINPUT77), .Z(n296) );
  XNOR2_X1 U349 ( .A(KEYINPUT76), .B(KEYINPUT9), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n310) );
  XOR2_X1 U351 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n298) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n299), .B(KEYINPUT10), .Z(n304) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n300), .B(KEYINPUT7), .ZN(n321) );
  XOR2_X1 U357 ( .A(G92GAT), .B(G218GAT), .Z(n302) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n386) );
  XNOR2_X1 U360 ( .A(n321), .B(n386), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U362 ( .A(G99GAT), .B(G106GAT), .Z(n327) );
  XOR2_X1 U363 ( .A(n305), .B(n327), .Z(n308) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(G134GAT), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n306), .B(G85GAT), .ZN(n401) );
  XNOR2_X1 U367 ( .A(n420), .B(n401), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n568) );
  INV_X1 U370 ( .A(n568), .ZN(n367) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G29GAT), .Z(n312) );
  XNOR2_X1 U372 ( .A(G50GAT), .B(G36GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U374 ( .A(KEYINPUT29), .B(G1GAT), .Z(n314) );
  XNOR2_X1 U375 ( .A(G197GAT), .B(G113GAT), .ZN(n313) );
  XNOR2_X1 U376 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n325) );
  XOR2_X1 U378 ( .A(G169GAT), .B(G8GAT), .Z(n377) );
  XNOR2_X1 U379 ( .A(G22GAT), .B(G15GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n317), .B(KEYINPUT69), .ZN(n359) );
  XOR2_X1 U381 ( .A(n377), .B(n359), .Z(n319) );
  NAND2_X1 U382 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U384 ( .A(n320), .B(KEYINPUT68), .Z(n323) );
  XNOR2_X1 U385 ( .A(n321), .B(KEYINPUT30), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n578) );
  AND2_X1 U388 ( .A1(G230GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n329) );
  XNOR2_X1 U390 ( .A(G120GAT), .B(G148GAT), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n328), .B(G57GAT), .ZN(n400) );
  XOR2_X1 U392 ( .A(n350), .B(G92GAT), .Z(n333) );
  XOR2_X1 U393 ( .A(KEYINPUT71), .B(G78GAT), .Z(n417) );
  XNOR2_X1 U394 ( .A(n417), .B(G85GAT), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U396 ( .A(n334), .B(KEYINPUT72), .Z(n335) );
  XNOR2_X1 U397 ( .A(n336), .B(n335), .ZN(n341) );
  INV_X1 U398 ( .A(n341), .ZN(n339) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(G64GAT), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n337), .B(KEYINPUT73), .ZN(n380) );
  XOR2_X1 U401 ( .A(n380), .B(KEYINPUT31), .Z(n340) );
  INV_X1 U402 ( .A(n340), .ZN(n338) );
  NAND2_X1 U403 ( .A1(n339), .A2(n338), .ZN(n343) );
  NAND2_X1 U404 ( .A1(n341), .A2(n340), .ZN(n342) );
  NAND2_X1 U405 ( .A1(n343), .A2(n342), .ZN(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n345) );
  XNOR2_X1 U407 ( .A(KEYINPUT70), .B(KEYINPUT75), .ZN(n344) );
  NOR2_X1 U408 ( .A1(n578), .A2(n562), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n347), .B(KEYINPUT46), .ZN(n364) );
  XOR2_X1 U410 ( .A(G64GAT), .B(G211GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(G183GAT), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n363) );
  XOR2_X1 U413 ( .A(n350), .B(n408), .Z(n352) );
  XNOR2_X1 U414 ( .A(G155GAT), .B(G78GAT), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n357) );
  XOR2_X1 U416 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n354) );
  XNOR2_X1 U417 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U419 ( .A(n358), .B(KEYINPUT15), .Z(n361) );
  XNOR2_X1 U420 ( .A(n359), .B(G57GAT), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  INV_X1 U422 ( .A(n565), .ZN(n587) );
  NOR2_X1 U423 ( .A1(n364), .A2(n587), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT109), .ZN(n366) );
  NOR2_X1 U425 ( .A1(n367), .A2(n366), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U427 ( .A(KEYINPUT78), .B(n568), .ZN(n572) );
  XNOR2_X1 U428 ( .A(KEYINPUT36), .B(n572), .ZN(n500) );
  NOR2_X1 U429 ( .A1(n565), .A2(n500), .ZN(n370) );
  XOR2_X1 U430 ( .A(KEYINPUT45), .B(n370), .Z(n371) );
  NOR2_X1 U431 ( .A1(n584), .A2(n371), .ZN(n372) );
  NAND2_X1 U432 ( .A1(n372), .A2(n578), .ZN(n373) );
  NAND2_X1 U433 ( .A1(n374), .A2(n373), .ZN(n376) );
  XOR2_X1 U434 ( .A(KEYINPUT93), .B(n377), .Z(n379) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U437 ( .A(n381), .B(n380), .Z(n388) );
  XNOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT86), .ZN(n383) );
  XOR2_X1 U440 ( .A(n383), .B(KEYINPUT87), .Z(n385) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G204GAT), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n425) );
  XNOR2_X1 U443 ( .A(n425), .B(n386), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U445 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U448 ( .A(KEYINPUT19), .B(n391), .ZN(n450) );
  XNOR2_X1 U449 ( .A(n392), .B(n450), .ZN(n530) );
  XNOR2_X1 U450 ( .A(KEYINPUT54), .B(n393), .ZN(n412) );
  XOR2_X1 U451 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n395) );
  XNOR2_X1 U452 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U454 ( .A(G141GAT), .B(n396), .Z(n429) );
  XOR2_X1 U455 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n398) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U458 ( .A(n399), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U460 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT90), .B(KEYINPUT1), .Z(n405) );
  XNOR2_X1 U462 ( .A(G162GAT), .B(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U464 ( .A(n407), .B(n406), .Z(n410) );
  XOR2_X1 U465 ( .A(G113GAT), .B(KEYINPUT0), .Z(n442) );
  XNOR2_X1 U466 ( .A(n442), .B(n408), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n429), .B(n411), .ZN(n483) );
  XNOR2_X1 U469 ( .A(KEYINPUT92), .B(n483), .ZN(n528) );
  NAND2_X1 U470 ( .A1(n412), .A2(n528), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n413), .B(KEYINPUT64), .ZN(n464) );
  XOR2_X1 U472 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n415) );
  XNOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U475 ( .A(n416), .B(G106GAT), .Z(n419) );
  XNOR2_X1 U476 ( .A(n417), .B(G218GAT), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U478 ( .A(n420), .B(G148GAT), .Z(n422) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n427) );
  XNOR2_X1 U482 ( .A(G22GAT), .B(n425), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n478) );
  NOR2_X1 U485 ( .A1(n464), .A2(n478), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n430), .B(KEYINPUT55), .ZN(n451) );
  XOR2_X1 U487 ( .A(KEYINPUT81), .B(KEYINPUT65), .Z(n432) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U490 ( .A(G71GAT), .B(KEYINPUT83), .Z(n434) );
  XNOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n448) );
  XOR2_X1 U494 ( .A(G120GAT), .B(G127GAT), .Z(n438) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G176GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n446) );
  XOR2_X1 U497 ( .A(G99GAT), .B(G134GAT), .Z(n440) );
  XNOR2_X1 U498 ( .A(G43GAT), .B(G190GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U500 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U501 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n538) );
  OR2_X1 U506 ( .A1(n292), .A2(n451), .ZN(n457) );
  XOR2_X1 U507 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n452) );
  XOR2_X1 U509 ( .A(n453), .B(n452), .Z(n455) );
  XOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT121), .Z(n454) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  INV_X1 U512 ( .A(n578), .ZN(n515) );
  NAND2_X1 U513 ( .A1(n515), .A2(n570), .ZN(n461) );
  XNOR2_X1 U514 ( .A(G169GAT), .B(KEYINPUT119), .ZN(n459) );
  INV_X1 U515 ( .A(KEYINPUT120), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U517 ( .A(KEYINPUT126), .ZN(n466) );
  XOR2_X1 U518 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n463) );
  NAND2_X1 U519 ( .A1(n538), .A2(n478), .ZN(n462) );
  XNOR2_X1 U520 ( .A(n463), .B(n462), .ZN(n555) );
  NOR2_X1 U521 ( .A1(n464), .A2(n555), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n583) );
  NOR2_X1 U523 ( .A1(n583), .A2(n500), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n471) );
  XNOR2_X1 U525 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(n489) );
  NOR2_X1 U527 ( .A1(n578), .A2(n584), .ZN(n503) );
  NAND2_X1 U528 ( .A1(n572), .A2(n587), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT16), .B(n472), .Z(n487) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(n478), .ZN(n494) );
  XNOR2_X1 U531 ( .A(n530), .B(KEYINPUT94), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT27), .ZN(n480) );
  NOR2_X1 U533 ( .A1(n480), .A2(n528), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT95), .ZN(n554) );
  NOR2_X1 U535 ( .A1(n494), .A2(n554), .ZN(n540) );
  XNOR2_X1 U536 ( .A(KEYINPUT96), .B(n540), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n475), .A2(n538), .ZN(n486) );
  NOR2_X1 U538 ( .A1(n538), .A2(n530), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  NOR2_X1 U540 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n479), .B(KEYINPUT25), .ZN(n482) );
  OR2_X1 U542 ( .A1(n555), .A2(n480), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n482), .A2(n481), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n498) );
  AND2_X1 U546 ( .A1(n487), .A2(n498), .ZN(n516) );
  NAND2_X1 U547 ( .A1(n503), .A2(n516), .ZN(n495) );
  NOR2_X1 U548 ( .A1(n528), .A2(n495), .ZN(n488) );
  XOR2_X1 U549 ( .A(n489), .B(n488), .Z(G1324GAT) );
  NOR2_X1 U550 ( .A1(n530), .A2(n495), .ZN(n490) );
  XOR2_X1 U551 ( .A(G8GAT), .B(n490), .Z(G1325GAT) );
  NOR2_X1 U552 ( .A1(n538), .A2(n495), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U555 ( .A(G15GAT), .B(n493), .Z(G1326GAT) );
  INV_X1 U556 ( .A(n494), .ZN(n534) );
  NOR2_X1 U557 ( .A1(n534), .A2(n495), .ZN(n496) );
  XOR2_X1 U558 ( .A(KEYINPUT102), .B(n496), .Z(n497) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XNOR2_X1 U560 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n506) );
  NAND2_X1 U561 ( .A1(n565), .A2(n498), .ZN(n499) );
  NOR2_X1 U562 ( .A1(n500), .A2(n499), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n527) );
  NAND2_X1 U565 ( .A1(n503), .A2(n527), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(KEYINPUT38), .ZN(n513) );
  NOR2_X1 U567 ( .A1(n528), .A2(n513), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G29GAT), .B(n507), .ZN(G1328GAT) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n530), .A2(n513), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  XNOR2_X1 U573 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n511) );
  NOR2_X1 U574 ( .A1(n538), .A2(n513), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U576 ( .A(G43GAT), .B(n512), .Z(G1330GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n534), .ZN(n514) );
  XOR2_X1 U578 ( .A(G50GAT), .B(n514), .Z(G1331GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n562), .ZN(n526) );
  AND2_X1 U580 ( .A1(n516), .A2(n526), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(KEYINPUT107), .ZN(n523) );
  NOR2_X1 U582 ( .A1(n528), .A2(n523), .ZN(n519) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U585 ( .A(G57GAT), .B(n520), .Z(G1332GAT) );
  NOR2_X1 U586 ( .A1(n530), .A2(n523), .ZN(n521) );
  XOR2_X1 U587 ( .A(G64GAT), .B(n521), .Z(G1333GAT) );
  NOR2_X1 U588 ( .A1(n538), .A2(n523), .ZN(n522) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n522), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n534), .A2(n523), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n528), .A2(n533), .ZN(n529) );
  XOR2_X1 U595 ( .A(G85GAT), .B(n529), .Z(G1336GAT) );
  NOR2_X1 U596 ( .A1(n530), .A2(n533), .ZN(n531) );
  XOR2_X1 U597 ( .A(G92GAT), .B(n531), .Z(G1337GAT) );
  NOR2_X1 U598 ( .A1(n538), .A2(n533), .ZN(n532) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n532), .Z(G1338GAT) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n535), .Z(n536) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n538), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(KEYINPUT112), .B(n541), .ZN(n549) );
  NOR2_X1 U606 ( .A1(n578), .A2(n549), .ZN(n542) );
  XOR2_X1 U607 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U608 ( .A1(n549), .A2(n562), .ZN(n544) );
  XNOR2_X1 U609 ( .A(KEYINPUT113), .B(KEYINPUT49), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U611 ( .A(G120GAT), .B(n545), .Z(G1341GAT) );
  XNOR2_X1 U612 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n547) );
  NOR2_X1 U613 ( .A1(n565), .A2(n549), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n572), .ZN(n553) );
  XOR2_X1 U617 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n551) );
  XNOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT115), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  INV_X1 U621 ( .A(n537), .ZN(n557) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n567) );
  NOR2_X1 U624 ( .A1(n578), .A2(n567), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n561) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n562), .A2(n567), .ZN(n563) );
  XOR2_X1 U631 ( .A(n564), .B(n563), .Z(G1345GAT) );
  NOR2_X1 U632 ( .A1(n565), .A2(n567), .ZN(n566) );
  XOR2_X1 U633 ( .A(G155GAT), .B(n566), .Z(G1346GAT) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(G162GAT), .B(n569), .Z(G1347GAT) );
  NAND2_X1 U636 ( .A1(n587), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n577) );
  XNOR2_X1 U639 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT58), .B(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1351GAT) );
  NOR2_X1 U643 ( .A1(n583), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U649 ( .A(n583), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n584), .A2(n588), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
endmodule

