//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(KEYINPUT25), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n206), .B1(KEYINPUT23), .B2(new_n202), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(new_n214), .C1(new_n208), .C2(KEYINPUT64), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n204), .B(new_n207), .C1(new_n210), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(new_n206), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT26), .ZN(new_n222));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT27), .B(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT68), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n219), .B(new_n224), .C1(new_n228), .C2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT27), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(G183gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n233), .A2(new_n225), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n229), .B(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n216), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n205), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n213), .A2(new_n214), .ZN(new_n247));
  OR2_X1    g046(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n249), .A3(new_n223), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n203), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n240), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n239), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n255));
  XNOR2_X1  g054(.A(G127gat), .B(G134gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(G127gat), .A2(G134gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n260));
  INV_X1    g059(.A(G134gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT70), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G113gat), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT1), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n258), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n264), .ZN(new_n275));
  OAI21_X1  g074(.A(G134gat), .B1(new_n275), .B2(new_n262), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n257), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n222), .B(new_n223), .C1(new_n218), .C2(new_n206), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n235), .B2(new_n237), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n228), .A2(new_n230), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n243), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n284), .A2(new_n247), .A3(new_n209), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n281), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n247), .A2(new_n250), .ZN(new_n287));
  INV_X1    g086(.A(new_n203), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n242), .A2(KEYINPUT65), .A3(new_n205), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT65), .B1(new_n242), .B2(new_n205), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT25), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT70), .B1(new_n260), .B2(new_n265), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n267), .A3(new_n276), .ZN(new_n295));
  AOI22_X1  g094(.A1(new_n294), .A2(new_n295), .B1(new_n255), .B2(new_n256), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G227gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n279), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT32), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT33), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G15gat), .B(G43gat), .Z(new_n305));
  XNOR2_X1  g104(.A(G71gat), .B(G99gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n301), .B(KEYINPUT32), .C1(new_n303), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n300), .B1(new_n279), .B2(new_n297), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT34), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI211_X1 g113(.A(KEYINPUT34), .B(new_n300), .C1(new_n279), .C2(new_n297), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n311), .B1(KEYINPUT71), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n314), .A2(new_n315), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n308), .A4(new_n310), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n308), .A3(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n311), .A2(new_n316), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT36), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n286), .B2(new_n292), .ZN(new_n328));
  INV_X1    g127(.A(G226gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(new_n299), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT73), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n239), .B2(new_n252), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n337), .A2(KEYINPUT22), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G197gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G197gat), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n341), .A2(new_n343), .A3(G204gat), .ZN(new_n344));
  AOI21_X1  g143(.A(G204gat), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(G211gat), .A2(G218gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G204gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n342), .A2(G197gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n340), .A2(KEYINPUT72), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n341), .A2(new_n343), .A3(G204gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n348), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n339), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n293), .B2(new_n330), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n336), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  NOR2_X1   g165(.A1(new_n328), .A2(new_n330), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n253), .A2(new_n335), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n359), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT74), .A4(new_n360), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n363), .A2(new_n366), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n370), .A2(new_n369), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n366), .A4(new_n363), .ZN(new_n375));
  INV_X1    g174(.A(new_n366), .ZN(new_n376));
  INV_X1    g175(.A(new_n363), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n369), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n373), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  INV_X1    g180(.A(G141gat), .ZN(new_n382));
  INV_X1    g181(.A(G148gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G162gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G155gat), .ZN(new_n386));
  INV_X1    g185(.A(G155gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G162gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(G141gat), .A2(G148gat), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n384), .A2(new_n386), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G155gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n393));
  OAI21_X1  g192(.A(G162gat), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n390), .B1(new_n394), .B2(KEYINPUT2), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n384), .A2(new_n389), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT2), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n396), .A2(new_n397), .B1(new_n386), .B2(new_n388), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n381), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n386), .A2(new_n388), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n389), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n400), .B1(new_n401), .B2(KEYINPUT2), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT75), .B(G155gat), .Z(new_n403));
  AOI21_X1  g202(.A(new_n397), .B1(new_n403), .B2(G162gat), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT77), .B(new_n402), .C1(new_n404), .C2(new_n390), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT4), .B1(new_n406), .B2(new_n278), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n395), .A2(new_n398), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n296), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n395), .B2(new_n398), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n413), .B(new_n402), .C1(new_n404), .C2(new_n390), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT76), .B1(new_n415), .B2(new_n296), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n278), .A2(new_n417), .A3(new_n414), .A4(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n411), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT78), .ZN(new_n422));
  INV_X1    g221(.A(new_n409), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n278), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n296), .A2(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n420), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n422), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n294), .A2(new_n295), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n430), .A2(new_n409), .A3(new_n257), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n409), .B1(new_n430), .B2(new_n257), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n421), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n429), .B1(new_n416), .B2(new_n418), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT4), .B1(new_n278), .B2(new_n423), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n296), .A2(new_n408), .A3(new_n399), .A4(new_n405), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n439), .B1(new_n437), .B2(new_n438), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n427), .B(new_n436), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G1gat), .B(G29gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n444), .B(KEYINPUT0), .ZN(new_n445));
  XNOR2_X1  g244(.A(G57gat), .B(G85gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n445), .B(new_n446), .Z(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n435), .A2(new_n442), .A3(new_n447), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n447), .B1(new_n435), .B2(new_n442), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n380), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT31), .B(G50gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n409), .B2(new_n413), .ZN(new_n459));
  OAI211_X1 g258(.A(G228gat), .B(G233gat), .C1(new_n459), .C2(new_n358), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n356), .B1(new_n355), .B2(new_n339), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n348), .B(new_n338), .C1(new_n353), .C2(new_n354), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n332), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT80), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n358), .A2(KEYINPUT80), .A3(new_n332), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n413), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n460), .B1(new_n467), .B2(new_n423), .ZN(new_n468));
  INV_X1    g267(.A(new_n414), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n359), .B1(new_n469), .B2(KEYINPUT29), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n349), .B2(new_n357), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n406), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n470), .A2(new_n472), .B1(G228gat), .B2(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G22gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n463), .A2(new_n413), .B1(new_n399), .B2(new_n405), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n459), .A2(new_n358), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT3), .B1(new_n463), .B2(new_n464), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n409), .B1(new_n481), .B2(new_n466), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n480), .B1(new_n482), .B2(new_n460), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(G22gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n458), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n468), .B2(new_n473), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n480), .B(KEYINPUT81), .C1(new_n482), .C2(new_n460), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(KEYINPUT82), .A3(G22gat), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n458), .B1(new_n474), .B2(new_n475), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n475), .B1(new_n483), .B2(new_n486), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT82), .B1(new_n492), .B2(new_n488), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n485), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n327), .B1(new_n455), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n447), .B(KEYINPUT83), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n419), .B1(new_n440), .B2(new_n441), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n429), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(KEYINPUT39), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT40), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n424), .A2(new_n425), .A3(new_n420), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT39), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n498), .B2(new_n429), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n500), .A2(new_n501), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n443), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n435), .A2(KEYINPUT84), .A3(new_n442), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(new_n496), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n373), .A2(new_n375), .A3(new_n379), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n501), .B1(new_n500), .B2(new_n504), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n505), .A2(new_n509), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n512), .A2(new_n494), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n377), .A2(new_n378), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT37), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n366), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n515), .B2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT38), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n451), .A3(new_n450), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n367), .A2(new_n368), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n515), .B1(new_n520), .B2(new_n358), .ZN(new_n521));
  INV_X1    g320(.A(new_n368), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(new_n331), .A3(new_n336), .A4(new_n359), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n516), .A2(new_n524), .B1(new_n366), .B2(new_n514), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n518), .A2(new_n519), .A3(new_n449), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n495), .B1(new_n513), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n494), .A2(new_n380), .A3(new_n454), .A4(new_n321), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n528), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n323), .A2(new_n324), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n534), .A2(new_n510), .A3(KEYINPUT35), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n449), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n494), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n527), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT87), .B(G36gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n541), .A2(G29gat), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G43gat), .ZN(new_n549));
  INV_X1    g348(.A(G43gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G50gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n551), .A3(KEYINPUT15), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n554), .A3(KEYINPUT15), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n547), .A3(new_n553), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT86), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n546), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n559), .A3(new_n545), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n541), .A2(G29gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n556), .A2(new_n564), .A3(KEYINPUT89), .ZN(new_n568));
  XNOR2_X1  g367(.A(G15gat), .B(G22gat), .ZN(new_n569));
  INV_X1    g368(.A(G1gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT16), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(G1gat), .B2(new_n569), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G8gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n568), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT90), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT90), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n567), .A2(new_n577), .A3(new_n568), .A4(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n565), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n574), .B1(new_n582), .B2(KEYINPUT17), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n584), .A3(new_n568), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(KEYINPUT18), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n568), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT89), .B1(new_n556), .B2(new_n564), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n590), .A2(new_n574), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n580), .B(KEYINPUT13), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n587), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n586), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n598), .A3(new_n586), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n594), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n596), .A2(new_n597), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT92), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n340), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT11), .B(G169gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  INV_X1    g409(.A(KEYINPUT93), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n612), .B(new_n587), .C1(new_n592), .C2(new_n593), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n603), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n587), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n593), .B1(new_n579), .B2(new_n591), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n615), .A2(new_n610), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT93), .A3(new_n600), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n605), .A2(new_n610), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n538), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT100), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n628), .A2(new_n631), .A3(new_n632), .A4(new_n624), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT7), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G99gat), .B(G106gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(G85gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n637), .A2(new_n630), .B1(KEYINPUT8), .B2(new_n638), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n636), .B1(new_n635), .B2(new_n639), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n623), .B1(new_n590), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n582), .A2(KEYINPUT17), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT102), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n635), .A2(new_n639), .ZN(new_n646));
  INV_X1    g445(.A(new_n636), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n585), .A2(new_n644), .A3(new_n645), .A4(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n622), .B1(new_n643), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n643), .A2(new_n652), .A3(new_n622), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G134gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n385), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n653), .B2(KEYINPUT103), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n654), .A2(KEYINPUT103), .A3(new_n655), .A4(new_n659), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n665));
  NAND2_X1  g464(.A1(G71gat), .A2(G78gat), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT95), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT9), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G57gat), .A2(G64gat), .ZN(new_n670));
  OR2_X1    g469(.A1(G57gat), .A2(G64gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n667), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n665), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g473(.A1(G71gat), .A2(G78gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n666), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n666), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n665), .B(new_n677), .C1(new_n672), .C2(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n574), .B1(KEYINPUT21), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT98), .ZN(new_n681));
  XNOR2_X1  g480(.A(G127gat), .B(G155gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NAND2_X1  g482(.A1(G231gat), .A2(G233gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT96), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n683), .B(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n681), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n679), .A2(KEYINPUT21), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(G183gat), .B(G211gat), .Z(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n687), .A2(new_n695), .A3(new_n696), .A4(new_n688), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n664), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT104), .B1(new_n663), .B2(new_n700), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n676), .B(new_n678), .C1(new_n640), .C2(new_n641), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n679), .A2(new_n648), .A3(new_n650), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT10), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n642), .A2(KEYINPUT10), .A3(new_n679), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(G230gat), .A2(G233gat), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n706), .ZN(new_n713));
  INV_X1    g512(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(G120gat), .B(G148gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(G176gat), .B(G204gat), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n710), .B2(new_n711), .ZN(new_n721));
  AOI211_X1 g520(.A(KEYINPUT105), .B(new_n714), .C1(new_n708), .C2(new_n709), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n713), .B2(new_n714), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n719), .B1(new_n724), .B2(new_n718), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n704), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n620), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n454), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(new_n570), .ZN(G1324gat));
  NOR2_X1   g530(.A1(new_n729), .A2(new_n380), .ZN(new_n732));
  XOR2_X1   g531(.A(KEYINPUT16), .B(G8gat), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(G8gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n732), .ZN(new_n736));
  MUX2_X1   g535(.A(new_n734), .B(new_n736), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g536(.A(G15gat), .B1(new_n729), .B2(new_n327), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n534), .A2(G15gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n729), .B2(new_n739), .ZN(G1326gat));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n729), .B2(new_n494), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n742));
  INV_X1    g541(.A(new_n494), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n620), .A2(new_n742), .A3(new_n743), .A4(new_n728), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT43), .B(G22gat), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n745), .B(new_n746), .Z(G1327gat));
  NAND4_X1  g546(.A1(new_n620), .A2(new_n663), .A3(new_n700), .A4(new_n726), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n748), .A2(G29gat), .A3(new_n454), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT44), .B1(new_n538), .B2(new_n664), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n528), .A2(KEYINPUT85), .A3(KEYINPUT35), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT85), .B1(new_n528), .B2(KEYINPUT35), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n537), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT108), .B(new_n537), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n527), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n664), .A2(KEYINPUT44), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n752), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n619), .A2(new_n701), .A3(new_n725), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n454), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n751), .B1(new_n543), .B2(new_n766), .ZN(G1328gat));
  AOI21_X1  g566(.A(new_n541), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n510), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n770), .B(new_n771), .Z(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n510), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n541), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(G1329gat));
  INV_X1    g574(.A(new_n327), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n762), .A2(new_n776), .A3(new_n763), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G43gat), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n748), .A2(G43gat), .A3(new_n534), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n779), .A3(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1330gat));
  NAND4_X1  g583(.A1(new_n762), .A2(G50gat), .A3(new_n743), .A4(new_n763), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n548), .B1(new_n748), .B2(new_n494), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g587(.A1(new_n703), .A2(new_n619), .A3(new_n704), .A4(new_n725), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n759), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n765), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G57gat), .ZN(G1332gat));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n793));
  INV_X1    g592(.A(G64gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n510), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT110), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n794), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1333gat));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n534), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n790), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n759), .A2(new_n327), .A3(new_n789), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n800), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n743), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  INV_X1    g606(.A(new_n619), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n701), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n726), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n762), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n454), .ZN(new_n813));
  INV_X1    g612(.A(new_n527), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT108), .B1(new_n533), .B2(new_n537), .ZN(new_n815));
  INV_X1    g614(.A(new_n758), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n663), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n757), .A2(new_n758), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n664), .B1(new_n822), .B2(new_n814), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n819), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n817), .A2(new_n663), .A3(new_n809), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n821), .A2(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n765), .A2(new_n637), .A3(new_n725), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n813), .A2(new_n637), .B1(new_n828), .B2(new_n829), .ZN(G1336gat));
  NAND3_X1  g629(.A1(new_n762), .A2(new_n510), .A3(new_n811), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(new_n831), .B2(G92gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n726), .A2(G92gat), .A3(new_n380), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n828), .B2(new_n834), .ZN(new_n835));
  XOR2_X1   g634(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n827), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n824), .B1(new_n823), .B2(new_n819), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n759), .A2(KEYINPUT111), .A3(new_n664), .A4(new_n818), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n840), .A2(new_n833), .B1(G92gat), .B2(new_n831), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n835), .B1(new_n841), .B2(new_n842), .ZN(G1337gat));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n826), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(new_n838), .B2(new_n839), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT113), .B(G99gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n801), .A3(new_n725), .A4(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n812), .A2(new_n327), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n848), .B2(new_n846), .ZN(G1338gat));
  NOR3_X1   g648(.A1(new_n726), .A2(G106gat), .A3(new_n494), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n821), .A2(new_n825), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n837), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n761), .B1(new_n822), .B2(new_n814), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT44), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n814), .A2(new_n755), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n663), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n743), .B(new_n811), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(G106gat), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT53), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n762), .A2(KEYINPUT114), .A3(new_n743), .A4(new_n811), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(G106gat), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n850), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n860), .A2(new_n867), .ZN(G1339gat));
  NAND2_X1  g667(.A1(new_n728), .A2(new_n619), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n614), .A2(new_n618), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n592), .A2(new_n593), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n583), .A2(new_n585), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n579), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n580), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n609), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n719), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n718), .B1(new_n723), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT55), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n710), .B2(new_n711), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n708), .A2(new_n714), .A3(new_n709), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n712), .A2(KEYINPUT105), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n710), .A2(new_n720), .A3(new_n711), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n878), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n718), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n881), .A2(new_n882), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n880), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n663), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n870), .A2(new_n725), .A3(new_n875), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n884), .A2(new_n891), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n619), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n896), .B2(new_n664), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n869), .B1(new_n897), .B2(new_n701), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n454), .A2(new_n510), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n898), .A2(new_n494), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n801), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n270), .A3(new_n619), .ZN(new_n902));
  INV_X1    g701(.A(new_n898), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(new_n454), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n494), .A2(new_n321), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n905), .A2(new_n510), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n808), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n270), .B2(new_n908), .ZN(G1340gat));
  AOI21_X1  g708(.A(G120gat), .B1(new_n907), .B2(new_n725), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n726), .A2(new_n268), .A3(new_n534), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n900), .B2(new_n911), .ZN(G1341gat));
  NAND4_X1  g711(.A1(new_n907), .A2(new_n263), .A3(new_n264), .A4(new_n701), .ZN(new_n913));
  OAI22_X1  g712(.A1(new_n901), .A2(new_n700), .B1(new_n262), .B2(new_n275), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1342gat));
  NOR2_X1   g714(.A1(new_n664), .A2(G134gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n904), .A2(new_n906), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n917), .A2(KEYINPUT56), .ZN(new_n918));
  OAI21_X1  g717(.A(G134gat), .B1(new_n901), .B2(new_n664), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(KEYINPUT56), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n918), .A2(KEYINPUT115), .A3(new_n919), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1343gat));
  NAND2_X1  g724(.A1(new_n327), .A2(new_n899), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT116), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n743), .A2(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n896), .A2(new_n664), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n930), .A2(KEYINPUT118), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n893), .B1(new_n930), .B2(KEYINPUT118), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n701), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n727), .A2(new_n808), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n929), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n936), .B1(new_n903), .B2(new_n494), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n927), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n382), .B1(new_n938), .B2(new_n808), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n776), .A2(new_n494), .A3(new_n510), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n904), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(G141gat), .A3(new_n619), .ZN(new_n942));
  OAI21_X1  g741(.A(KEYINPUT58), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n942), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT58), .ZN(new_n945));
  AOI211_X1 g744(.A(new_n619), .B(new_n927), .C1(new_n935), .C2(new_n937), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n382), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(new_n947), .ZN(G1344gat));
  OAI21_X1  g747(.A(KEYINPUT59), .B1(new_n941), .B2(new_n726), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n726), .A2(KEYINPUT59), .ZN(new_n950));
  AOI22_X1  g749(.A1(new_n949), .A2(new_n383), .B1(new_n938), .B2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n884), .A2(new_n891), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n614), .A2(new_n618), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n612), .B1(new_n602), .B2(new_n604), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n663), .B1(new_n955), .B2(new_n894), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n892), .A2(KEYINPUT120), .ZN(new_n957));
  AOI22_X1  g756(.A1(new_n614), .A2(new_n618), .B1(new_n609), .B2(new_n874), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n884), .A2(new_n663), .A3(new_n891), .A4(new_n959), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n700), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n494), .B1(new_n962), .B2(new_n869), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT121), .B1(new_n963), .B2(KEYINPUT57), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n930), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n934), .B1(new_n968), .B2(new_n700), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(new_n494), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n964), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n494), .A2(new_n936), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n898), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n898), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AOI211_X1 g778(.A(new_n726), .B(new_n927), .C1(new_n972), .C2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n951), .B1(new_n980), .B2(new_n981), .ZN(G1345gat));
  NAND2_X1  g781(.A1(new_n938), .A2(new_n701), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n403), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n700), .A2(new_n403), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n984), .B1(new_n941), .B2(new_n985), .ZN(G1346gat));
  AND2_X1   g785(.A1(new_n938), .A2(new_n663), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n663), .A2(new_n385), .ZN(new_n988));
  OAI22_X1  g787(.A1(new_n987), .A2(new_n385), .B1(new_n941), .B2(new_n988), .ZN(G1347gat));
  NOR2_X1   g788(.A1(new_n903), .A2(new_n765), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n905), .A2(new_n380), .ZN(new_n991));
  AND2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n992), .A2(new_n220), .A3(new_n808), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n903), .A2(new_n743), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n454), .A2(new_n510), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT123), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n999), .A2(new_n534), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(G169gat), .B1(new_n1001), .B2(new_n619), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n995), .A2(new_n1002), .ZN(G1348gat));
  NAND3_X1  g802(.A1(new_n992), .A2(new_n221), .A3(new_n725), .ZN(new_n1004));
  OAI21_X1  g803(.A(G176gat), .B1(new_n1001), .B2(new_n726), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT124), .ZN(G1349gat));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n227), .A3(new_n701), .ZN(new_n1008));
  OAI21_X1  g807(.A(G183gat), .B1(new_n1001), .B2(new_n700), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g810(.A1(new_n992), .A2(new_n212), .A3(new_n663), .ZN(new_n1012));
  OAI21_X1  g811(.A(G190gat), .B1(new_n1001), .B2(new_n664), .ZN(new_n1013));
  AND2_X1   g812(.A1(new_n1013), .A2(KEYINPUT61), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1013), .A2(KEYINPUT61), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1351gat));
  NAND3_X1  g815(.A1(new_n327), .A2(new_n743), .A3(new_n510), .ZN(new_n1017));
  XNOR2_X1  g816(.A(new_n1017), .B(KEYINPUT125), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n990), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g818(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g819(.A(G197gat), .B1(new_n1020), .B2(new_n808), .ZN(new_n1021));
  NOR2_X1   g820(.A1(new_n999), .A2(new_n776), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1022), .B1(new_n971), .B2(new_n978), .ZN(new_n1023));
  INV_X1    g822(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g823(.A1(new_n619), .A2(new_n340), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(G1352gat));
  NOR3_X1   g825(.A1(new_n1019), .A2(G204gat), .A3(new_n726), .ZN(new_n1027));
  XNOR2_X1  g826(.A(new_n1027), .B(KEYINPUT62), .ZN(new_n1028));
  OAI21_X1  g827(.A(G204gat), .B1(new_n1023), .B2(new_n726), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1353gat));
  OR3_X1    g829(.A1(new_n1019), .A2(G211gat), .A3(new_n700), .ZN(new_n1031));
  OAI211_X1 g830(.A(new_n701), .B(new_n1022), .C1(new_n971), .C2(new_n978), .ZN(new_n1032));
  AND3_X1   g831(.A1(new_n1032), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1033));
  AOI21_X1  g832(.A(KEYINPUT63), .B1(new_n1032), .B2(G211gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(G1354gat));
  AOI21_X1  g834(.A(G218gat), .B1(new_n1020), .B2(new_n663), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n663), .A2(G218gat), .ZN(new_n1037));
  XNOR2_X1  g836(.A(new_n1037), .B(KEYINPUT126), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n1036), .B1(new_n1024), .B2(new_n1038), .ZN(G1355gat));
endmodule


