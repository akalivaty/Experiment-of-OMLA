

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821;

  XOR2_X1 U376 ( .A(KEYINPUT7), .B(G107), .Z(n536) );
  XNOR2_X1 U377 ( .A(G146), .B(G101), .ZN(n565) );
  XNOR2_X1 U378 ( .A(KEYINPUT16), .B(G122), .ZN(n519) );
  NAND2_X2 U379 ( .A1(n405), .A2(n777), .ZN(n736) );
  NAND2_X2 U380 ( .A1(n744), .A2(G953), .ZN(n799) );
  XNOR2_X2 U381 ( .A(n486), .B(n740), .ZN(n742) );
  XNOR2_X2 U382 ( .A(n424), .B(n417), .ZN(n790) );
  INV_X2 U383 ( .A(G125), .ZN(n513) );
  XNOR2_X2 U384 ( .A(n513), .B(G146), .ZN(n407) );
  XNOR2_X2 U385 ( .A(n355), .B(KEYINPUT72), .ZN(n562) );
  INV_X4 U386 ( .A(G131), .ZN(n355) );
  XNOR2_X1 U387 ( .A(G125), .B(G146), .ZN(n359) );
  NAND2_X1 U388 ( .A1(G234), .A2(G237), .ZN(n515) );
  INV_X1 U389 ( .A(G237), .ZN(n528) );
  XOR2_X1 U390 ( .A(G122), .B(KEYINPUT12), .Z(n543) );
  XNOR2_X1 U391 ( .A(G116), .B(G122), .ZN(n535) );
  INV_X1 U392 ( .A(G104), .ZN(n751) );
  NAND2_X2 U393 ( .A1(n796), .A2(n760), .ZN(n428) );
  XNOR2_X2 U394 ( .A(n734), .B(KEYINPUT85), .ZN(n487) );
  NOR2_X1 U395 ( .A1(n711), .A2(n483), .ZN(n482) );
  INV_X4 U396 ( .A(G953), .ZN(n778) );
  NAND2_X1 U397 ( .A1(n365), .A2(n381), .ZN(n364) );
  NAND2_X1 U398 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U399 ( .A1(n476), .A2(n482), .ZN(n777) );
  NAND2_X1 U400 ( .A1(n361), .A2(n360), .ZN(n711) );
  AND2_X1 U401 ( .A1(n375), .A2(n373), .ZN(n360) );
  XNOR2_X1 U402 ( .A(n510), .B(n509), .ZN(n820) );
  XNOR2_X1 U403 ( .A(n607), .B(n606), .ZN(n726) );
  NOR2_X1 U404 ( .A1(n600), .A2(n633), .ZN(n545) );
  INV_X1 U405 ( .A(n594), .ZN(n679) );
  OR2_X1 U406 ( .A1(KEYINPUT32), .A2(n647), .ZN(n409) );
  BUF_X1 U407 ( .A(n583), .Z(n714) );
  XNOR2_X1 U408 ( .A(n716), .B(KEYINPUT38), .ZN(n594) );
  NOR2_X1 U409 ( .A1(n644), .A2(n643), .ZN(n489) );
  NOR2_X1 U410 ( .A1(n441), .A2(G902), .ZN(n455) );
  NAND2_X1 U411 ( .A1(n416), .A2(KEYINPUT84), .ZN(n381) );
  INV_X1 U412 ( .A(G113), .ZN(n492) );
  NAND2_X1 U413 ( .A1(n390), .A2(n387), .ZN(n395) );
  NAND2_X1 U414 ( .A1(n389), .A2(n388), .ZN(n387) );
  AND2_X1 U415 ( .A1(n393), .A2(n391), .ZN(n390) );
  NAND2_X1 U416 ( .A1(n368), .A2(n364), .ZN(n737) );
  XNOR2_X1 U417 ( .A(n657), .B(n656), .ZN(n733) );
  NAND2_X1 U418 ( .A1(n448), .A2(n445), .ZN(n657) );
  XNOR2_X1 U419 ( .A(n446), .B(n511), .ZN(n445) );
  NAND2_X1 U420 ( .A1(n447), .A2(n468), .ZN(n446) );
  NAND2_X1 U421 ( .A1(n711), .A2(KEYINPUT48), .ZN(n479) );
  INV_X1 U422 ( .A(n480), .ZN(n477) );
  AND2_X1 U423 ( .A1(n374), .A2(n699), .ZN(n361) );
  AND2_X1 U424 ( .A1(n641), .A2(n759), .ZN(n468) );
  NOR2_X1 U425 ( .A1(n821), .A2(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U426 ( .A1(n702), .A2(n679), .ZN(n681) );
  XNOR2_X1 U427 ( .A(n671), .B(KEYINPUT42), .ZN(n821) );
  XNOR2_X1 U428 ( .A(n404), .B(KEYINPUT101), .ZN(n626) );
  AND2_X1 U429 ( .A1(n379), .A2(n629), .ZN(n378) );
  NAND2_X1 U430 ( .A1(n594), .A2(n684), .ZN(n600) );
  XNOR2_X1 U431 ( .A(n489), .B(KEYINPUT105), .ZN(n633) );
  XNOR2_X1 U432 ( .A(n507), .B(n506), .ZN(n629) );
  NOR2_X1 U433 ( .A1(n586), .A2(n632), .ZN(n507) );
  XNOR2_X1 U434 ( .A(n455), .B(n490), .ZN(n643) );
  AND2_X1 U435 ( .A1(n392), .A2(n799), .ZN(n391) );
  INV_X1 U436 ( .A(n788), .ZN(n388) );
  OR2_X1 U437 ( .A1(n788), .A2(G472), .ZN(n392) );
  XNOR2_X1 U438 ( .A(n540), .B(n539), .ZN(n441) );
  INV_X1 U439 ( .A(n416), .ZN(n382) );
  NAND2_X1 U440 ( .A1(n735), .A2(KEYINPUT2), .ZN(n416) );
  NAND2_X1 U441 ( .A1(n530), .A2(G210), .ZN(n529) );
  XNOR2_X1 U442 ( .A(n492), .B(G143), .ZN(n491) );
  INV_X1 U443 ( .A(n359), .ZN(n442) );
  XNOR2_X1 U444 ( .A(G110), .B(KEYINPUT96), .ZN(n546) );
  XNOR2_X1 U445 ( .A(G119), .B(G128), .ZN(n549) );
  XNOR2_X1 U446 ( .A(KEYINPUT11), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U447 ( .A(G902), .B(KEYINPUT15), .ZN(n732) );
  XNOR2_X2 U448 ( .A(n356), .B(n518), .ZN(n579) );
  XNOR2_X2 U449 ( .A(n358), .B(n357), .ZN(n356) );
  XNOR2_X2 U450 ( .A(G101), .B(KEYINPUT73), .ZN(n357) );
  XNOR2_X2 U451 ( .A(G116), .B(G113), .ZN(n358) );
  XNOR2_X1 U452 ( .A(n570), .B(n386), .ZN(n385) );
  NAND2_X1 U453 ( .A1(n798), .A2(n555), .ZN(n508) );
  XNOR2_X1 U454 ( .A(n362), .B(n775), .ZN(n798) );
  XNOR2_X1 U455 ( .A(n363), .B(n553), .ZN(n362) );
  XNOR2_X1 U456 ( .A(n551), .B(n550), .ZN(n363) );
  NOR2_X1 U457 ( .A1(n482), .A2(n382), .ZN(n366) );
  INV_X1 U458 ( .A(n476), .ZN(n367) );
  NAND2_X1 U459 ( .A1(n371), .A2(n369), .ZN(n368) );
  NAND2_X1 U460 ( .A1(n487), .A2(n370), .ZN(n369) );
  NAND2_X1 U461 ( .A1(n478), .A2(n472), .ZN(n370) );
  NAND2_X1 U462 ( .A1(n372), .A2(KEYINPUT84), .ZN(n371) );
  INV_X1 U463 ( .A(n487), .ZN(n372) );
  NAND2_X1 U464 ( .A1(n820), .A2(KEYINPUT46), .ZN(n373) );
  NAND2_X1 U465 ( .A1(n821), .A2(KEYINPUT46), .ZN(n374) );
  NAND2_X1 U466 ( .A1(n377), .A2(n376), .ZN(n375) );
  INV_X1 U467 ( .A(n820), .ZN(n377) );
  NAND2_X1 U468 ( .A1(n629), .A2(n423), .ZN(n676) );
  NAND2_X1 U469 ( .A1(n677), .A2(n378), .ZN(n678) );
  AND2_X1 U470 ( .A1(n423), .A2(n380), .ZN(n379) );
  INV_X1 U471 ( .A(n675), .ZN(n380) );
  NAND2_X1 U472 ( .A1(n527), .A2(n732), .ZN(n444) );
  XNOR2_X1 U473 ( .A(n383), .B(n514), .ZN(n527) );
  XNOR2_X1 U474 ( .A(n485), .B(n384), .ZN(n383) );
  XNOR2_X1 U475 ( .A(n523), .B(n522), .ZN(n384) );
  XNOR2_X2 U476 ( .A(n532), .B(n526), .ZN(n485) );
  XNOR2_X1 U477 ( .A(n579), .B(n385), .ZN(n514) );
  INV_X1 U478 ( .A(n519), .ZN(n386) );
  INV_X1 U479 ( .A(n421), .ZN(n389) );
  NAND2_X1 U480 ( .A1(n421), .A2(n394), .ZN(n393) );
  AND2_X1 U481 ( .A1(n788), .A2(G472), .ZN(n394) );
  XNOR2_X1 U482 ( .A(n395), .B(n789), .ZN(G57) );
  INV_X1 U483 ( .A(n597), .ZN(n396) );
  BUF_X1 U484 ( .A(n460), .Z(n397) );
  NAND2_X1 U485 ( .A1(n454), .A2(n453), .ZN(n398) );
  BUF_X1 U486 ( .A(n451), .Z(n399) );
  AND2_X2 U487 ( .A1(n494), .A2(n495), .ZN(n454) );
  INV_X1 U488 ( .A(n716), .ZN(n400) );
  XNOR2_X1 U489 ( .A(n508), .B(n559), .ZN(n586) );
  XNOR2_X1 U490 ( .A(n444), .B(n529), .ZN(n401) );
  XNOR2_X1 U491 ( .A(n444), .B(n529), .ZN(n617) );
  BUF_X1 U492 ( .A(n760), .Z(n402) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n403) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n552) );
  NAND2_X1 U495 ( .A1(n605), .A2(n672), .ZN(n404) );
  AND2_X1 U496 ( .A1(n766), .A2(KEYINPUT2), .ZN(n405) );
  AND2_X1 U497 ( .A1(n766), .A2(n777), .ZN(n722) );
  NOR2_X1 U498 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U499 ( .A1(n397), .A2(n458), .ZN(n406) );
  NAND2_X1 U500 ( .A1(n460), .A2(n458), .ZN(n694) );
  BUF_X1 U501 ( .A(n411), .Z(n408) );
  NOR2_X1 U502 ( .A1(n692), .A2(n647), .ZN(n410) );
  NOR2_X1 U503 ( .A1(n409), .A2(n692), .ZN(n470) );
  XNOR2_X2 U504 ( .A(n637), .B(n412), .ZN(n411) );
  XOR2_X1 U505 ( .A(KEYINPUT74), .B(KEYINPUT22), .Z(n412) );
  NAND2_X1 U506 ( .A1(n430), .A2(n429), .ZN(n796) );
  BUF_X1 U507 ( .A(n733), .Z(n766) );
  XNOR2_X2 U508 ( .A(n419), .B(KEYINPUT65), .ZN(n421) );
  XNOR2_X2 U509 ( .A(n418), .B(KEYINPUT65), .ZN(n422) );
  XNOR2_X2 U510 ( .A(n738), .B(KEYINPUT65), .ZN(n801) );
  OR2_X1 U511 ( .A1(n480), .A2(n475), .ZN(n474) );
  XNOR2_X1 U512 ( .A(n434), .B(n432), .ZN(n747) );
  XNOR2_X1 U513 ( .A(n544), .B(n433), .ZN(n432) );
  XNOR2_X1 U514 ( .A(n554), .B(n435), .ZN(n434) );
  XNOR2_X1 U515 ( .A(n491), .B(n493), .ZN(n433) );
  INV_X1 U516 ( .A(KEYINPUT19), .ZN(n462) );
  OR2_X1 U517 ( .A1(n684), .A2(n462), .ZN(n461) );
  INV_X1 U518 ( .A(n482), .ZN(n478) );
  NOR2_X1 U519 ( .A1(n474), .A2(n473), .ZN(n472) );
  INV_X1 U520 ( .A(KEYINPUT69), .ZN(n506) );
  XNOR2_X1 U521 ( .A(n443), .B(n624), .ZN(n636) );
  XNOR2_X1 U522 ( .A(n623), .B(KEYINPUT0), .ZN(n624) );
  NAND2_X1 U523 ( .A1(n694), .A2(n622), .ZN(n443) );
  NAND2_X1 U524 ( .A1(n778), .A2(G234), .ZN(n439) );
  OR2_X2 U525 ( .A1(n747), .A2(G902), .ZN(n456) );
  INV_X1 U526 ( .A(G478), .ZN(n490) );
  XNOR2_X1 U527 ( .A(n747), .B(n746), .ZN(n748) );
  INV_X1 U528 ( .A(KEYINPUT88), .ZN(n511) );
  INV_X1 U529 ( .A(n479), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT95), .B(KEYINPUT77), .Z(n566) );
  NAND2_X1 U531 ( .A1(n502), .A2(n501), .ZN(n500) );
  INV_X1 U532 ( .A(G469), .ZN(n502) );
  INV_X1 U533 ( .A(G902), .ZN(n501) );
  NAND2_X1 U534 ( .A1(G902), .A2(G469), .ZN(n504) );
  INV_X1 U535 ( .A(G902), .ZN(n555) );
  XNOR2_X1 U536 ( .A(G146), .B(G137), .ZN(n574) );
  XOR2_X1 U537 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n575) );
  NAND2_X1 U538 ( .A1(n481), .A2(n414), .ZN(n480) );
  OR2_X1 U539 ( .A1(n710), .A2(KEYINPUT48), .ZN(n483) );
  XOR2_X1 U540 ( .A(G137), .B(G140), .Z(n568) );
  XNOR2_X1 U541 ( .A(n562), .B(n436), .ZN(n435) );
  XNOR2_X1 U542 ( .A(n541), .B(n437), .ZN(n436) );
  INV_X1 U543 ( .A(G140), .ZN(n541) );
  INV_X1 U544 ( .A(G104), .ZN(n437) );
  XNOR2_X1 U545 ( .A(KEYINPUT70), .B(KEYINPUT4), .ZN(n526) );
  AND2_X1 U546 ( .A1(n684), .A2(n462), .ZN(n459) );
  XNOR2_X1 U547 ( .A(KEYINPUT3), .B(G119), .ZN(n518) );
  INV_X1 U548 ( .A(n726), .ZN(n498) );
  OR2_X1 U549 ( .A1(n721), .A2(n720), .ZN(n723) );
  XNOR2_X1 U550 ( .A(n628), .B(n627), .ZN(n761) );
  XNOR2_X1 U551 ( .A(n678), .B(KEYINPUT76), .ZN(n702) );
  XNOR2_X1 U552 ( .A(n787), .B(n786), .ZN(n788) );
  INV_X1 U553 ( .A(n771), .ZN(n431) );
  XOR2_X1 U554 ( .A(G134), .B(KEYINPUT9), .Z(n537) );
  INV_X1 U555 ( .A(KEYINPUT40), .ZN(n509) );
  NAND2_X1 U556 ( .A1(n470), .A2(n411), .ZN(n429) );
  BUF_X1 U557 ( .A(n761), .Z(n764) );
  NAND2_X1 U558 ( .A1(n408), .A2(n471), .ZN(n760) );
  NOR2_X1 U559 ( .A1(n714), .A2(n648), .ZN(n471) );
  INV_X1 U560 ( .A(KEYINPUT60), .ZN(n466) );
  INV_X1 U561 ( .A(KEYINPUT124), .ZN(n464) );
  XNOR2_X1 U562 ( .A(n814), .B(G146), .ZN(G48) );
  XOR2_X1 U563 ( .A(KEYINPUT13), .B(G475), .Z(n413) );
  AND2_X1 U564 ( .A1(n817), .A2(n818), .ZN(n414) );
  OR2_X1 U565 ( .A1(KEYINPUT44), .A2(KEYINPUT89), .ZN(n415) );
  XOR2_X1 U566 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n417) );
  INV_X1 U567 ( .A(KEYINPUT84), .ZN(n475) );
  NAND2_X1 U568 ( .A1(n737), .A2(n736), .ZN(n418) );
  NAND2_X1 U569 ( .A1(n737), .A2(n736), .ZN(n419) );
  NAND2_X1 U570 ( .A1(n737), .A2(n736), .ZN(n738) );
  BUF_X1 U571 ( .A(n654), .Z(n420) );
  OR2_X1 U572 ( .A1(n499), .A2(n503), .ZN(n423) );
  AND2_X1 U573 ( .A1(n583), .A2(n629), .ZN(n605) );
  BUF_X1 U574 ( .A(n527), .Z(n424) );
  XNOR2_X1 U575 ( .A(n451), .B(n573), .ZN(n425) );
  XNOR2_X1 U576 ( .A(n452), .B(n646), .ZN(n426) );
  INV_X1 U577 ( .A(n498), .ZN(n427) );
  XNOR2_X1 U578 ( .A(n451), .B(n573), .ZN(n741) );
  XNOR2_X1 U579 ( .A(n398), .B(n646), .ZN(n795) );
  NAND2_X1 U580 ( .A1(n454), .A2(n453), .ZN(n452) );
  AND2_X1 U581 ( .A1(n514), .A2(n431), .ZN(n772) );
  XNOR2_X1 U582 ( .A(n442), .B(n521), .ZN(n522) );
  XNOR2_X2 U583 ( .A(n428), .B(KEYINPUT90), .ZN(n654) );
  NAND2_X1 U584 ( .A1(n469), .A2(KEYINPUT32), .ZN(n430) );
  XNOR2_X1 U585 ( .A(n583), .B(KEYINPUT91), .ZN(n692) );
  XNOR2_X2 U586 ( .A(n669), .B(KEYINPUT1), .ZN(n583) );
  XNOR2_X1 U587 ( .A(n407), .B(KEYINPUT10), .ZN(n554) );
  XNOR2_X2 U588 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n440) );
  XNOR2_X1 U589 ( .A(n802), .B(n441), .ZN(n804) );
  AND2_X2 U590 ( .A1(n463), .A2(n461), .ZN(n460) );
  NAND2_X1 U591 ( .A1(n512), .A2(KEYINPUT44), .ZN(n447) );
  NAND2_X1 U592 ( .A1(n449), .A2(n655), .ZN(n448) );
  NAND2_X1 U593 ( .A1(n450), .A2(KEYINPUT66), .ZN(n449) );
  NAND2_X1 U594 ( .A1(n651), .A2(n650), .ZN(n450) );
  NAND2_X1 U595 ( .A1(n626), .A2(n625), .ZN(n628) );
  XNOR2_X1 U596 ( .A(n399), .B(n776), .ZN(n780) );
  XNOR2_X2 U597 ( .A(n582), .B(n564), .ZN(n451) );
  NAND2_X1 U598 ( .A1(n497), .A2(n498), .ZN(n453) );
  XNOR2_X2 U599 ( .A(n456), .B(n413), .ZN(n644) );
  NAND2_X1 U600 ( .A1(n457), .A2(n459), .ZN(n458) );
  INV_X1 U601 ( .A(n401), .ZN(n457) );
  NAND2_X1 U602 ( .A1(n617), .A2(KEYINPUT19), .ZN(n463) );
  XNOR2_X1 U603 ( .A(n465), .B(n464), .ZN(G54) );
  NAND2_X1 U604 ( .A1(n745), .A2(n799), .ZN(n465) );
  XNOR2_X1 U605 ( .A(n467), .B(n466), .ZN(G60) );
  NAND2_X1 U606 ( .A1(n750), .A2(n799), .ZN(n467) );
  OR2_X2 U607 ( .A1(n499), .A2(n503), .ZN(n669) );
  XNOR2_X2 U608 ( .A(n485), .B(n563), .ZN(n582) );
  NAND2_X1 U609 ( .A1(n411), .A2(n410), .ZN(n469) );
  NAND2_X1 U610 ( .A1(n710), .A2(KEYINPUT48), .ZN(n481) );
  NAND2_X1 U611 ( .A1(n477), .A2(n479), .ZN(n476) );
  NAND2_X1 U612 ( .A1(n672), .A2(n684), .ZN(n673) );
  XNOR2_X2 U613 ( .A(n484), .B(G472), .ZN(n672) );
  OR2_X2 U614 ( .A1(n787), .A2(G902), .ZN(n484) );
  XNOR2_X1 U615 ( .A(n582), .B(n581), .ZN(n787) );
  BUF_X1 U616 ( .A(n425), .Z(n486) );
  NAND2_X1 U617 ( .A1(n505), .A2(n504), .ZN(n503) );
  XNOR2_X2 U618 ( .A(n488), .B(n751), .ZN(n570) );
  XNOR2_X2 U619 ( .A(G110), .B(G107), .ZN(n488) );
  NAND2_X1 U620 ( .A1(n726), .A2(KEYINPUT34), .ZN(n494) );
  AND2_X1 U621 ( .A1(n496), .A2(n645), .ZN(n495) );
  NAND2_X1 U622 ( .A1(n642), .A2(KEYINPUT34), .ZN(n496) );
  NOR2_X1 U623 ( .A1(n642), .A2(KEYINPUT34), .ZN(n497) );
  NOR2_X1 U624 ( .A1(n425), .A2(n500), .ZN(n499) );
  NAND2_X1 U625 ( .A1(n741), .A2(G469), .ZN(n505) );
  NAND2_X1 U626 ( .A1(n712), .A2(n682), .ZN(n510) );
  INV_X1 U627 ( .A(n795), .ZN(n512) );
  XNOR2_X2 U628 ( .A(n525), .B(n524), .ZN(n532) );
  XNOR2_X1 U629 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n556) );
  INV_X1 U630 ( .A(KEYINPUT23), .ZN(n548) );
  XNOR2_X1 U631 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U632 ( .A(n731), .B(n730), .ZN(G75) );
  XOR2_X1 U633 ( .A(KEYINPUT93), .B(KEYINPUT14), .Z(n517) );
  XNOR2_X1 U634 ( .A(KEYINPUT75), .B(n515), .ZN(n516) );
  XNOR2_X1 U635 ( .A(n517), .B(n516), .ZN(n659) );
  NAND2_X1 U636 ( .A1(n778), .A2(G224), .ZN(n520) );
  XNOR2_X1 U637 ( .A(n520), .B(KEYINPUT18), .ZN(n523) );
  XNOR2_X1 U638 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n521) );
  XNOR2_X2 U639 ( .A(G143), .B(KEYINPUT80), .ZN(n525) );
  INV_X1 U640 ( .A(G128), .ZN(n524) );
  NAND2_X1 U641 ( .A1(n555), .A2(n528), .ZN(n530) );
  BUF_X1 U642 ( .A(n401), .Z(n716) );
  NAND2_X1 U643 ( .A1(n530), .A2(G214), .ZN(n531) );
  XNOR2_X1 U644 ( .A(n531), .B(KEYINPUT92), .ZN(n684) );
  NAND2_X1 U645 ( .A1(n552), .A2(G217), .ZN(n534) );
  INV_X1 U646 ( .A(n532), .ZN(n533) );
  XNOR2_X1 U647 ( .A(n534), .B(n533), .ZN(n540) );
  XNOR2_X1 U648 ( .A(n536), .B(n535), .ZN(n538) );
  XNOR2_X1 U649 ( .A(n538), .B(n537), .ZN(n539) );
  NOR2_X2 U650 ( .A1(G953), .A2(G237), .ZN(n576) );
  NAND2_X1 U651 ( .A1(G214), .A2(n576), .ZN(n542) );
  XNOR2_X1 U652 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U653 ( .A(n545), .B(KEYINPUT41), .ZN(n727) );
  XOR2_X1 U654 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n547) );
  XNOR2_X1 U655 ( .A(n547), .B(n546), .ZN(n551) );
  NAND2_X1 U656 ( .A1(n403), .A2(G221), .ZN(n553) );
  XNOR2_X1 U657 ( .A(n554), .B(n568), .ZN(n775) );
  NAND2_X1 U658 ( .A1(n732), .A2(G234), .ZN(n557) );
  XNOR2_X1 U659 ( .A(n557), .B(n556), .ZN(n560) );
  NAND2_X1 U660 ( .A1(G217), .A2(n560), .ZN(n558) );
  XNOR2_X1 U661 ( .A(n558), .B(KEYINPUT25), .ZN(n559) );
  NAND2_X1 U662 ( .A1(n560), .A2(G221), .ZN(n561) );
  XNOR2_X1 U663 ( .A(n561), .B(KEYINPUT21), .ZN(n665) );
  XOR2_X1 U664 ( .A(n665), .B(KEYINPUT99), .Z(n632) );
  XNOR2_X1 U665 ( .A(n562), .B(G134), .ZN(n563) );
  INV_X1 U666 ( .A(KEYINPUT94), .ZN(n564) );
  XNOR2_X1 U667 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U668 ( .A(n568), .B(n567), .Z(n572) );
  NAND2_X1 U669 ( .A1(n778), .A2(G227), .ZN(n569) );
  XNOR2_X1 U670 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U672 ( .A(n575), .B(n574), .ZN(n578) );
  NAND2_X1 U673 ( .A1(n576), .A2(G210), .ZN(n577) );
  XNOR2_X1 U674 ( .A(n578), .B(n577), .ZN(n580) );
  XNOR2_X1 U675 ( .A(n579), .B(n580), .ZN(n581) );
  INV_X1 U676 ( .A(n672), .ZN(n667) );
  NOR2_X1 U677 ( .A1(n629), .A2(n714), .ZN(n585) );
  XNOR2_X1 U678 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n584) );
  XNOR2_X1 U679 ( .A(n585), .B(n584), .ZN(n590) );
  BUF_X1 U680 ( .A(n586), .Z(n683) );
  NAND2_X1 U681 ( .A1(n665), .A2(n683), .ZN(n587) );
  XOR2_X1 U682 ( .A(KEYINPUT49), .B(n587), .Z(n588) );
  NAND2_X1 U683 ( .A1(n667), .A2(n588), .ZN(n589) );
  NOR2_X1 U684 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U685 ( .A1(n626), .A2(n591), .ZN(n592) );
  XOR2_X1 U686 ( .A(KEYINPUT51), .B(n592), .Z(n593) );
  NOR2_X1 U687 ( .A1(n727), .A2(n593), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n594), .A2(n684), .ZN(n595) );
  XOR2_X1 U689 ( .A(KEYINPUT119), .B(n595), .Z(n596) );
  NOR2_X1 U690 ( .A1(n633), .A2(n596), .ZN(n602) );
  INV_X1 U691 ( .A(n643), .ZN(n597) );
  AND2_X1 U692 ( .A1(n644), .A2(n597), .ZN(n682) );
  INV_X1 U693 ( .A(n682), .ZN(n599) );
  INV_X1 U694 ( .A(n644), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n598), .A2(n396), .ZN(n763) );
  AND2_X1 U696 ( .A1(n599), .A2(n763), .ZN(n703) );
  NOR2_X1 U697 ( .A1(n703), .A2(n600), .ZN(n601) );
  NOR2_X1 U698 ( .A1(n602), .A2(n601), .ZN(n608) );
  XNOR2_X1 U699 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n603) );
  XNOR2_X1 U700 ( .A(n672), .B(n603), .ZN(n688) );
  INV_X1 U701 ( .A(n688), .ZN(n604) );
  NAND2_X1 U702 ( .A1(n605), .A2(n604), .ZN(n607) );
  INV_X1 U703 ( .A(KEYINPUT33), .ZN(n606) );
  NOR2_X1 U704 ( .A1(n608), .A2(n427), .ZN(n609) );
  NOR2_X1 U705 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U706 ( .A(n611), .B(KEYINPUT52), .Z(n612) );
  XOR2_X1 U707 ( .A(KEYINPUT120), .B(n612), .Z(n613) );
  NOR2_X1 U708 ( .A1(n659), .A2(n613), .ZN(n614) );
  NAND2_X1 U709 ( .A1(n614), .A2(G952), .ZN(n615) );
  XNOR2_X1 U710 ( .A(KEYINPUT121), .B(n615), .ZN(n616) );
  NOR2_X1 U711 ( .A1(G953), .A2(n616), .ZN(n725) );
  NAND2_X1 U712 ( .A1(n778), .A2(G952), .ZN(n618) );
  NOR2_X1 U713 ( .A1(n659), .A2(n618), .ZN(n664) );
  INV_X1 U714 ( .A(G898), .ZN(n619) );
  AND2_X1 U715 ( .A1(n619), .A2(G953), .ZN(n771) );
  NAND2_X1 U716 ( .A1(n771), .A2(G902), .ZN(n620) );
  NOR2_X1 U717 ( .A1(n659), .A2(n620), .ZN(n621) );
  OR2_X1 U718 ( .A1(n664), .A2(n621), .ZN(n622) );
  INV_X1 U719 ( .A(KEYINPUT68), .ZN(n623) );
  BUF_X1 U720 ( .A(n636), .Z(n625) );
  XOR2_X1 U721 ( .A(KEYINPUT102), .B(KEYINPUT31), .Z(n627) );
  NOR2_X1 U722 ( .A1(n676), .A2(n672), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n630), .A2(n625), .ZN(n756) );
  NAND2_X1 U724 ( .A1(n761), .A2(n756), .ZN(n631) );
  INV_X1 U725 ( .A(n703), .ZN(n696) );
  NAND2_X1 U726 ( .A1(n631), .A2(n696), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n634), .B(KEYINPUT106), .ZN(n635) );
  NAND2_X1 U728 ( .A1(n636), .A2(n635), .ZN(n637) );
  INV_X1 U729 ( .A(n683), .ZN(n638) );
  NAND2_X1 U730 ( .A1(n688), .A2(n638), .ZN(n639) );
  NOR2_X1 U731 ( .A1(n714), .A2(n639), .ZN(n640) );
  NAND2_X1 U732 ( .A1(n408), .A2(n640), .ZN(n759) );
  INV_X1 U733 ( .A(n625), .ZN(n642) );
  NAND2_X1 U734 ( .A1(n644), .A2(n396), .ZN(n700) );
  XNOR2_X1 U735 ( .A(KEYINPUT79), .B(n700), .ZN(n645) );
  XOR2_X1 U736 ( .A(KEYINPUT86), .B(KEYINPUT35), .Z(n646) );
  INV_X1 U737 ( .A(KEYINPUT44), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n688), .A2(n683), .ZN(n647) );
  NAND2_X1 U739 ( .A1(n683), .A2(n667), .ZN(n648) );
  XNOR2_X1 U740 ( .A(n654), .B(n415), .ZN(n651) );
  NOR2_X1 U741 ( .A1(n426), .A2(KEYINPUT44), .ZN(n649) );
  INV_X1 U742 ( .A(n649), .ZN(n650) );
  NOR2_X1 U743 ( .A1(n652), .A2(KEYINPUT66), .ZN(n653) );
  NAND2_X1 U744 ( .A1(n420), .A2(n653), .ZN(n655) );
  XNOR2_X1 U745 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n656) );
  NAND2_X1 U746 ( .A1(G953), .A2(G902), .ZN(n658) );
  NOR2_X1 U747 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U748 ( .A(KEYINPUT108), .B(n660), .Z(n661) );
  NOR2_X1 U749 ( .A1(G900), .A2(n661), .ZN(n662) );
  XOR2_X1 U750 ( .A(KEYINPUT109), .B(n662), .Z(n663) );
  NOR2_X1 U751 ( .A1(n664), .A2(n663), .ZN(n675) );
  NOR2_X1 U752 ( .A1(n665), .A2(n675), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n686), .A2(n683), .ZN(n666) );
  NOR2_X1 U754 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U755 ( .A(KEYINPUT28), .B(n668), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n670), .A2(n423), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n727), .A2(n693), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n674) );
  XNOR2_X1 U759 ( .A(n674), .B(n673), .ZN(n677) );
  INV_X1 U760 ( .A(KEYINPUT39), .ZN(n680) );
  XNOR2_X1 U761 ( .A(n681), .B(n680), .ZN(n712) );
  XNOR2_X1 U762 ( .A(n682), .B(KEYINPUT107), .ZN(n810) );
  AND2_X1 U763 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U765 ( .A1(n810), .A2(n687), .ZN(n689) );
  NAND2_X1 U766 ( .A1(n689), .A2(n604), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n713), .A2(n716), .ZN(n690) );
  XOR2_X1 U768 ( .A(KEYINPUT36), .B(n690), .Z(n691) );
  NOR2_X1 U769 ( .A1(n692), .A2(n691), .ZN(n815) );
  INV_X1 U770 ( .A(n693), .ZN(n695) );
  NAND2_X1 U771 ( .A1(n695), .A2(n406), .ZN(n705) );
  INV_X1 U772 ( .A(n705), .ZN(n812) );
  NAND2_X1 U773 ( .A1(n812), .A2(n696), .ZN(n697) );
  NOR2_X1 U774 ( .A1(KEYINPUT47), .A2(n697), .ZN(n698) );
  NOR2_X1 U775 ( .A1(n815), .A2(n698), .ZN(n699) );
  OR2_X1 U776 ( .A1(n700), .A2(n716), .ZN(n701) );
  NOR2_X1 U777 ( .A1(n702), .A2(n701), .ZN(n808) );
  NAND2_X1 U778 ( .A1(n703), .A2(KEYINPUT47), .ZN(n704) );
  XOR2_X1 U779 ( .A(n704), .B(KEYINPUT83), .Z(n707) );
  NAND2_X1 U780 ( .A1(n705), .A2(KEYINPUT47), .ZN(n706) );
  NAND2_X1 U781 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U782 ( .A1(n808), .A2(n708), .ZN(n709) );
  XOR2_X1 U783 ( .A(KEYINPUT82), .B(n709), .Z(n710) );
  INV_X1 U784 ( .A(n763), .ZN(n805) );
  NAND2_X1 U785 ( .A1(n712), .A2(n805), .ZN(n817) );
  NOR2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U787 ( .A(n715), .B(KEYINPUT43), .ZN(n717) );
  OR2_X1 U788 ( .A1(n717), .A2(n400), .ZN(n818) );
  NOR2_X1 U789 ( .A1(n722), .A2(KEYINPUT81), .ZN(n718) );
  NOR2_X1 U790 ( .A1(n718), .A2(KEYINPUT2), .ZN(n721) );
  INV_X1 U791 ( .A(KEYINPUT2), .ZN(n719) );
  NOR2_X1 U792 ( .A1(n719), .A2(KEYINPUT81), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n723), .A2(n736), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n727), .A2(n427), .ZN(n728) );
  NOR2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U797 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n730) );
  INV_X1 U798 ( .A(n732), .ZN(n735) );
  NAND2_X1 U799 ( .A1(n733), .A2(n735), .ZN(n734) );
  NAND2_X1 U800 ( .A1(n801), .A2(G469), .ZN(n743) );
  XNOR2_X1 U801 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n739) );
  XOR2_X1 U802 ( .A(n739), .B(KEYINPUT58), .Z(n740) );
  XNOR2_X1 U803 ( .A(n743), .B(n742), .ZN(n745) );
  INV_X1 U804 ( .A(G952), .ZN(n744) );
  NAND2_X1 U805 ( .A1(n422), .A2(G475), .ZN(n749) );
  XOR2_X1 U806 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n746) );
  XNOR2_X1 U807 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U808 ( .A1(n756), .A2(n810), .ZN(n752) );
  XNOR2_X1 U809 ( .A(n752), .B(n751), .ZN(G6) );
  XOR2_X1 U810 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n754) );
  XNOR2_X1 U811 ( .A(G107), .B(KEYINPUT113), .ZN(n753) );
  XNOR2_X1 U812 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U813 ( .A(KEYINPUT26), .B(n755), .Z(n758) );
  NOR2_X1 U814 ( .A1(n756), .A2(n763), .ZN(n757) );
  XOR2_X1 U815 ( .A(n758), .B(n757), .Z(G9) );
  XNOR2_X1 U816 ( .A(n759), .B(G101), .ZN(G3) );
  XNOR2_X1 U817 ( .A(n402), .B(G110), .ZN(G12) );
  NOR2_X1 U818 ( .A1(n764), .A2(n810), .ZN(n762) );
  XOR2_X1 U819 ( .A(G113), .B(n762), .Z(G15) );
  NOR2_X1 U820 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U821 ( .A(G116), .B(n765), .Z(G18) );
  NAND2_X1 U822 ( .A1(n766), .A2(n778), .ZN(n770) );
  NAND2_X1 U823 ( .A1(G953), .A2(G224), .ZN(n767) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n767), .ZN(n768) );
  NAND2_X1 U825 ( .A1(n768), .A2(G898), .ZN(n769) );
  NAND2_X1 U826 ( .A1(n770), .A2(n769), .ZN(n774) );
  XOR2_X1 U827 ( .A(KEYINPUT125), .B(n772), .Z(n773) );
  XNOR2_X1 U828 ( .A(n774), .B(n773), .ZN(G69) );
  XNOR2_X1 U829 ( .A(n775), .B(KEYINPUT126), .ZN(n776) );
  XOR2_X1 U830 ( .A(n780), .B(n777), .Z(n779) );
  NAND2_X1 U831 ( .A1(n779), .A2(n778), .ZN(n785) );
  XNOR2_X1 U832 ( .A(G227), .B(n780), .ZN(n781) );
  NAND2_X1 U833 ( .A1(n781), .A2(G900), .ZN(n782) );
  NAND2_X1 U834 ( .A1(G953), .A2(n782), .ZN(n783) );
  XOR2_X1 U835 ( .A(KEYINPUT127), .B(n783), .Z(n784) );
  NAND2_X1 U836 ( .A1(n785), .A2(n784), .ZN(G72) );
  XNOR2_X1 U837 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n786) );
  XNOR2_X1 U838 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n789) );
  NAND2_X1 U839 ( .A1(n801), .A2(G210), .ZN(n791) );
  XNOR2_X1 U840 ( .A(n791), .B(n790), .ZN(n792) );
  NAND2_X1 U841 ( .A1(n792), .A2(n799), .ZN(n794) );
  XNOR2_X1 U842 ( .A(KEYINPUT87), .B(KEYINPUT56), .ZN(n793) );
  XNOR2_X1 U843 ( .A(n794), .B(n793), .ZN(G51) );
  XNOR2_X1 U844 ( .A(n426), .B(G122), .ZN(G24) );
  XNOR2_X1 U845 ( .A(n796), .B(G119), .ZN(G21) );
  NAND2_X1 U846 ( .A1(n422), .A2(G217), .ZN(n797) );
  XOR2_X1 U847 ( .A(n798), .B(n797), .Z(n800) );
  INV_X1 U848 ( .A(n799), .ZN(n803) );
  NOR2_X1 U849 ( .A1(n800), .A2(n803), .ZN(G66) );
  NAND2_X1 U850 ( .A1(n421), .A2(G478), .ZN(n802) );
  NOR2_X1 U851 ( .A1(n804), .A2(n803), .ZN(G63) );
  XOR2_X1 U852 ( .A(G128), .B(KEYINPUT29), .Z(n807) );
  NAND2_X1 U853 ( .A1(n812), .A2(n805), .ZN(n806) );
  XNOR2_X1 U854 ( .A(n807), .B(n806), .ZN(G30) );
  XNOR2_X1 U855 ( .A(G143), .B(n808), .ZN(n809) );
  XNOR2_X1 U856 ( .A(n809), .B(KEYINPUT115), .ZN(G45) );
  INV_X1 U857 ( .A(n810), .ZN(n811) );
  NAND2_X1 U858 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U859 ( .A(n813), .B(KEYINPUT116), .ZN(n814) );
  XNOR2_X1 U860 ( .A(G125), .B(n815), .ZN(n816) );
  XNOR2_X1 U861 ( .A(n816), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U862 ( .A(G134), .B(n817), .ZN(G36) );
  XOR2_X1 U863 ( .A(n818), .B(G140), .Z(n819) );
  XNOR2_X1 U864 ( .A(n819), .B(KEYINPUT117), .ZN(G42) );
  XOR2_X1 U865 ( .A(G131), .B(n820), .Z(G33) );
  XOR2_X1 U866 ( .A(G137), .B(n821), .Z(G39) );
endmodule

