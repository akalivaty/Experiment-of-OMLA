//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(G107), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G104), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT3), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT77), .B(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT78), .B1(new_n187), .B2(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G107), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT79), .B1(new_n193), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n191), .B(G104), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n194), .A2(new_n197), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(new_n189), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n199), .A2(G101), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n202), .A2(new_n203), .A3(new_n207), .A4(new_n189), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT4), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n199), .A2(new_n205), .A3(KEYINPUT4), .A4(G101), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G116), .ZN(new_n222));
  INV_X1    g036(.A(G116), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G119), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT2), .B(G113), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT66), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n217), .B2(new_n218), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n220), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n225), .B2(new_n226), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n218), .A3(new_n228), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n220), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n212), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n190), .A2(new_n196), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n188), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n208), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n243));
  INV_X1    g057(.A(new_n222), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n213), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n225), .B2(new_n243), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n234), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G122), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n238), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n210), .A2(new_n211), .B1(new_n236), .B2(new_n231), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n248), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n254), .A3(KEYINPUT6), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n256), .B(new_n252), .C1(new_n253), .C2(new_n248), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT64), .A3(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT0), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n261), .A2(G146), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  OR2_X1    g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n259), .A2(G143), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n264), .B(new_n269), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G125), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  OAI21_X1  g088(.A(G128), .B1(new_n266), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n266), .B2(new_n270), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n263), .A2(new_n274), .A3(G128), .A4(new_n267), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT82), .B(G224), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n284), .A3(new_n280), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n255), .A2(new_n257), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n242), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT5), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n245), .B1(new_n294), .B2(new_n225), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n234), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n250), .B(KEYINPUT8), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n297), .B(new_n298), .C1(new_n293), .C2(new_n247), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n273), .A2(new_n280), .A3(new_n290), .A4(new_n284), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n292), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n301), .B2(new_n251), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n289), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G210), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n289), .A2(new_n302), .A3(new_n304), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(KEYINPUT83), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n303), .A2(new_n309), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT84), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n308), .A2(new_n315), .A3(new_n312), .A4(new_n310), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT70), .B(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n321), .B(KEYINPUT76), .ZN(new_n322));
  INV_X1    g136(.A(G227), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(G953), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n322), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n212), .A2(new_n272), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n276), .A2(new_n277), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT10), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n242), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n266), .B1(new_n260), .B2(new_n262), .ZN(new_n331));
  INV_X1    g145(.A(new_n275), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n277), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n241), .A3(new_n208), .ZN(new_n334));
  XOR2_X1   g148(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n330), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT65), .ZN(new_n340));
  INV_X1    g154(.A(G134), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G137), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT11), .ZN(new_n343));
  INV_X1    g157(.A(G137), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n344), .A2(G134), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT11), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n340), .B(new_n347), .C1(new_n341), .C2(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n343), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G131), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n343), .A2(new_n351), .A3(new_n346), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n268), .A2(new_n271), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n210), .B2(new_n211), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n337), .ZN(new_n357));
  INV_X1    g171(.A(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(new_n330), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n325), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n242), .A2(new_n327), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n361), .B2(new_n334), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n362), .B(new_n363), .ZN(new_n364));
  NOR4_X1   g178(.A1(new_n356), .A2(new_n337), .A3(new_n353), .A4(new_n329), .ZN(new_n365));
  INV_X1    g179(.A(new_n325), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n318), .B(new_n320), .C1(new_n360), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(G469), .A2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n354), .A2(new_n359), .A3(new_n325), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n366), .B1(new_n364), .B2(new_n365), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G469), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT9), .B(G234), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G221), .B1(new_n375), .B2(G902), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(KEYINPUT75), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(G234), .A2(G237), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(G952), .A3(new_n283), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n319), .A2(G953), .A3(new_n380), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT21), .B(G898), .Z(new_n383));
  OAI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G140), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G125), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n386), .A2(KEYINPUT73), .A3(G125), .ZN(new_n390));
  XNOR2_X1  g204(.A(G125), .B(G140), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  OAI211_X1 g208(.A(G146), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(G237), .A2(G953), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n396), .A2(G143), .A3(G214), .ZN(new_n397));
  AOI21_X1  g211(.A(G143), .B1(new_n396), .B2(G214), .ZN(new_n398));
  OAI21_X1  g212(.A(G131), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n283), .A3(G214), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n261), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n396), .A2(G143), .A3(G214), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n351), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n279), .A2(G140), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n387), .A2(new_n406), .A3(new_n392), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n386), .A2(KEYINPUT73), .A3(G125), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT19), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n391), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n259), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n391), .A2(new_n259), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n408), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT85), .B(new_n414), .C1(new_n415), .C2(new_n259), .ZN(new_n416));
  NAND2_X1  g230(.A1(KEYINPUT18), .A2(G131), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n397), .B2(new_n398), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n402), .A2(KEYINPUT18), .A3(G131), .A4(new_n403), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n393), .A2(new_n421), .A3(G146), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n196), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT86), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n424), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n394), .B1(new_n407), .B2(new_n408), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n259), .B1(new_n433), .B2(new_n388), .ZN(new_n434));
  OAI211_X1 g248(.A(KEYINPUT17), .B(G131), .C1(new_n397), .C2(new_n398), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n395), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT87), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n405), .A2(KEYINPUT17), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n395), .A3(new_n435), .A4(KEYINPUT87), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n426), .A3(new_n423), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G475), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n445), .B2(KEYINPUT20), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(KEYINPUT89), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n441), .A2(new_n426), .A3(new_n423), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n430), .B1(new_n424), .B2(new_n427), .ZN(new_n450));
  AOI211_X1 g264(.A(KEYINPUT86), .B(new_n426), .C1(new_n413), .C2(new_n423), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT88), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n432), .A2(new_n454), .A3(new_n442), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n445), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n448), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(KEYINPUT90), .B(G475), .Z(new_n459));
  AOI21_X1  g273(.A(new_n426), .B1(new_n441), .B2(new_n423), .ZN(new_n460));
  OR2_X1    g274(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G902), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n458), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n223), .A3(G122), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT92), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G116), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(G116), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n466), .ZN(new_n472));
  OAI21_X1  g286(.A(G107), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n470), .ZN(new_n475));
  XNOR2_X1  g289(.A(G128), .B(G143), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(G134), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n476), .A2(new_n341), .ZN(new_n479));
  OAI221_X1 g293(.A(new_n473), .B1(new_n190), .B2(new_n475), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n475), .B(new_n190), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n477), .A2(KEYINPUT91), .A3(G134), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT13), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n261), .A3(G128), .ZN(new_n484));
  OAI211_X1 g298(.A(G134), .B(new_n484), .C1(new_n477), .C2(new_n483), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT91), .B1(new_n477), .B2(G134), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n481), .A2(new_n482), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n374), .A2(G217), .A3(new_n283), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n480), .B2(new_n487), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n320), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT93), .B(new_n320), .C1(new_n491), .C2(new_n492), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n493), .A2(new_n497), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR4_X1   g315(.A1(new_n379), .A2(new_n385), .A3(new_n465), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n353), .A2(new_n272), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n341), .A2(G137), .ZN(new_n504));
  OAI21_X1  g318(.A(G131), .B1(new_n345), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n278), .A2(new_n352), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n503), .A2(new_n231), .A3(new_n236), .A4(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(G101), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n396), .A2(G210), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n352), .A2(new_n505), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n276), .B2(new_n277), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n355), .B1(new_n350), .B2(new_n352), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT30), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n503), .B2(new_n506), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n237), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT68), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n507), .A2(new_n521), .A3(new_n511), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT31), .ZN(new_n524));
  INV_X1    g338(.A(new_n511), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  AOI211_X1 g340(.A(KEYINPUT67), .B(new_n219), .C1(new_n233), .C2(new_n232), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n235), .B1(new_n234), .B2(new_n220), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n515), .A2(new_n516), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n526), .B1(new_n529), .B2(new_n507), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n515), .A2(new_n516), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT28), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n525), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT31), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n513), .A2(new_n520), .A3(new_n535), .A4(new_n522), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n524), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(G472), .A2(G902), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT32), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G472), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n507), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT28), .ZN(new_n543));
  INV_X1    g357(.A(new_n533), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n511), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n546), .A2(KEYINPUT29), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n520), .ZN(new_n550));
  INV_X1    g364(.A(new_n507), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n525), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n543), .A2(new_n547), .A3(new_n544), .A4(new_n511), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n541), .B1(new_n554), .B2(new_n320), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT32), .B1(new_n537), .B2(new_n538), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n540), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G128), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT23), .B1(new_n558), .B2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(G119), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(KEYINPUT71), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT71), .ZN(new_n562));
  OAI211_X1 g376(.A(G119), .B(new_n558), .C1(new_n562), .C2(KEYINPUT23), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT72), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT72), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G110), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT24), .B(G110), .Z(new_n569));
  XNOR2_X1  g383(.A(G119), .B(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n572));
  AOI21_X1  g386(.A(G146), .B1(new_n572), .B2(new_n389), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n433), .A2(new_n259), .A3(new_n388), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n568), .B(new_n571), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n564), .A2(G110), .B1(new_n570), .B2(new_n569), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n395), .A3(new_n414), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n575), .A2(KEYINPUT74), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT74), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT22), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n344), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AND4_X1   g397(.A1(KEYINPUT74), .A2(new_n575), .A3(new_n577), .A4(new_n582), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n320), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT25), .ZN(new_n586));
  INV_X1    g400(.A(G217), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n320), .B2(G234), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n575), .A2(new_n577), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT74), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n575), .A2(KEYINPUT74), .A3(new_n577), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n584), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n320), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n586), .A2(new_n588), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n588), .A2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n557), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n317), .A2(new_n502), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n537), .A2(new_n538), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n537), .A2(new_n320), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(G472), .ZN(new_n608));
  AOI211_X1 g422(.A(KEYINPUT94), .B(new_n541), .C1(new_n537), .C2(new_n320), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n610), .A2(new_n601), .A3(new_n379), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n480), .A2(new_n487), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n488), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n616), .B2(new_n490), .ZN(new_n617));
  OAI211_X1 g431(.A(G478), .B(new_n320), .C1(new_n613), .C2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n458), .B2(new_n464), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n304), .B1(new_n289), .B2(new_n302), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n313), .B1(new_n621), .B2(KEYINPUT95), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n306), .A2(new_n623), .A3(new_n307), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n620), .A2(new_n384), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n611), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT96), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n622), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n432), .A2(new_n454), .A3(new_n442), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n454), .B1(new_n432), .B2(new_n442), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n444), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT20), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n453), .A2(new_n455), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n457), .A3(new_n444), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n384), .A3(new_n464), .ZN(new_n639));
  INV_X1    g453(.A(new_n501), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n631), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n611), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  INV_X1    g458(.A(new_n610), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n589), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n599), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n598), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n317), .A2(new_n502), .A3(new_n645), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT37), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(G110), .Z(G12));
  NOR2_X1   g466(.A1(new_n557), .A2(new_n379), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n624), .A2(new_n622), .A3(new_n649), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n463), .B1(new_n635), .B2(new_n637), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n381), .B(KEYINPUT97), .ZN(new_n657));
  INV_X1    g471(.A(new_n382), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n656), .A2(new_n501), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XOR2_X1   g478(.A(new_n311), .B(KEYINPUT38), .Z(new_n665));
  INV_X1    g479(.A(new_n448), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n634), .B2(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n463), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n640), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n540), .A2(new_n556), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n542), .A2(new_n525), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n523), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n649), .A2(new_n313), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n665), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT98), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n660), .B(KEYINPUT39), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT40), .B1(new_n379), .B2(new_n680), .ZN(new_n681));
  OR3_X1    g495(.A1(new_n379), .A2(KEYINPUT40), .A3(new_n680), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT99), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(new_n261), .ZN(G45));
  NAND2_X1  g499(.A1(new_n612), .A2(new_n618), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n686), .B(new_n661), .C1(new_n667), .C2(new_n463), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n655), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G146), .ZN(G48));
  OAI21_X1  g504(.A(new_n320), .B1(new_n360), .B2(new_n367), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n378), .A3(new_n368), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n557), .A2(new_n601), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n626), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT41), .B(G113), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G15));
  NAND2_X1  g511(.A1(new_n641), .A2(new_n694), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G116), .ZN(G18));
  NOR3_X1   g513(.A1(new_n465), .A2(new_n385), .A3(new_n501), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n554), .A2(new_n320), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G472), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT32), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n605), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n704), .A3(new_n539), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n358), .B1(new_n357), .B2(new_n330), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n366), .B1(new_n706), .B2(new_n365), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n362), .B(KEYINPUT12), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n359), .A2(new_n708), .A3(new_n325), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n318), .B1(new_n710), .B2(new_n320), .ZN(new_n711));
  AOI211_X1 g525(.A(G469), .B(new_n319), .C1(new_n707), .C2(new_n709), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n377), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n654), .A2(new_n700), .A3(new_n705), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NAND2_X1  g529(.A1(new_n607), .A2(G472), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n605), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n601), .A3(new_n385), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n624), .A2(new_n622), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n669), .A4(new_n713), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G122), .ZN(G24));
  NAND3_X1  g535(.A1(new_n649), .A2(new_n716), .A3(new_n605), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n631), .A2(new_n722), .A3(new_n693), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n687), .A2(KEYINPUT100), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n465), .A2(new_n725), .A3(new_n686), .A4(new_n661), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  NAND2_X1  g543(.A1(new_n539), .A2(KEYINPUT102), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n537), .A2(new_n731), .A3(KEYINPUT32), .A4(new_n538), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n730), .A2(new_n702), .A3(new_n704), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  INV_X1    g548(.A(new_n601), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT42), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n311), .A2(new_n312), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n369), .B(KEYINPUT101), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n368), .A2(new_n372), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n378), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n727), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n739), .A2(new_n601), .A3(new_n557), .A4(new_n742), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT42), .B1(new_n746), .B2(new_n727), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n351), .ZN(G33));
  AND3_X1   g563(.A1(new_n743), .A2(new_n602), .A3(new_n662), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n341), .ZN(G36));
  NAND2_X1  g565(.A1(new_n610), .A2(new_n649), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT106), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n668), .A2(new_n686), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT105), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n680), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n370), .A2(new_n371), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n768), .B2(new_n740), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n740), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(KEYINPUT104), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n368), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n378), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n762), .A2(new_n763), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n313), .B1(new_n308), .B2(new_n310), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n760), .B2(new_n761), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT47), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n773), .B2(new_n378), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n773), .A2(new_n378), .A3(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n739), .A2(new_n705), .A3(new_n687), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n783), .A2(new_n601), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  NOR4_X1   g603(.A1(new_n754), .A2(new_n601), .A3(new_n313), .A4(new_n377), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT108), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n711), .A2(new_n712), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n674), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  INV_X1    g611(.A(new_n665), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n792), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n653), .B(new_n654), .C1(new_n662), .C2(new_n688), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n465), .A2(new_n624), .A3(new_n501), .A4(new_n622), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n649), .B1(new_n670), .B2(new_n673), .ZN(new_n803));
  INV_X1    g617(.A(new_n742), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n803), .A3(new_n804), .A4(new_n661), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n801), .A2(new_n728), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n801), .A2(new_n728), .A3(new_n805), .A4(KEYINPUT52), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n719), .A2(new_n384), .A3(new_n501), .A4(new_n656), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n713), .A2(new_n705), .A3(new_n735), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n714), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n719), .A2(new_n669), .A3(new_n713), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n717), .A2(new_n601), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n384), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n814), .A2(new_n816), .B1(new_n625), .B2(new_n812), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n656), .A2(new_n640), .A3(new_n661), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT111), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n649), .A3(new_n653), .A4(new_n776), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n818), .B(new_n821), .C1(new_n745), .C2(new_n747), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n810), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n465), .A2(new_n385), .A3(new_n640), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n317), .A2(new_n611), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n650), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT110), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n317), .A2(new_n384), .A3(new_n611), .A4(new_n620), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(new_n603), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n650), .A2(new_n825), .A3(KEYINPUT110), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n722), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n743), .A2(new_n727), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n743), .A2(KEYINPUT112), .A3(new_n727), .A4(new_n833), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n750), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n823), .A2(KEYINPUT53), .A3(new_n832), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n808), .A2(new_n809), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n698), .A2(new_n695), .A3(new_n714), .A4(new_n720), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n733), .A2(new_n735), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT103), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(KEYINPUT42), .A3(new_n727), .A4(new_n743), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT42), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n602), .A2(new_n776), .A3(new_n804), .ZN(new_n849));
  INV_X1    g663(.A(new_n727), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n842), .B1(new_n847), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n841), .A2(new_n852), .A3(new_n838), .A4(new_n821), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n828), .A2(new_n603), .A3(new_n829), .A4(new_n831), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n840), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT54), .B1(new_n839), .B2(new_n855), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n739), .A2(new_n693), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n735), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n381), .A3(new_n674), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n620), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n759), .A2(new_n657), .A3(new_n859), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n864), .A2(new_n722), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(new_n668), .A3(new_n619), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n757), .A2(new_n657), .A3(new_n815), .A4(new_n758), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n312), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n665), .A2(new_n693), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n868), .A2(KEYINPUT50), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT50), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n865), .B(new_n866), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n793), .A2(new_n377), .ZN(new_n873));
  INV_X1    g687(.A(new_n786), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n782), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n867), .A2(new_n739), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n863), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(G952), .A3(new_n283), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT113), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(KEYINPUT113), .B(new_n873), .C1(new_n874), .C2(new_n782), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n881), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n883), .A2(new_n863), .A3(new_n872), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n858), .A2(new_n862), .A3(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n867), .A2(new_n631), .A3(new_n693), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n864), .B1(new_n845), .B2(new_n844), .ZN(new_n888));
  NOR2_X1   g702(.A1(KEYINPUT114), .A2(KEYINPUT48), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(KEYINPUT114), .B2(KEYINPUT48), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n800), .B1(new_n892), .B2(new_n893), .ZN(G75));
  OR2_X1    g708(.A1(new_n283), .A2(G952), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT116), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n320), .B1(new_n839), .B2(new_n855), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT56), .B1(new_n897), .B2(new_n305), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n255), .A2(new_n257), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n288), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n901), .A2(new_n904), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(G51));
  INV_X1    g721(.A(new_n710), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n856), .A2(new_n857), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n740), .B(KEYINPUT117), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT57), .Z(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n839), .A2(new_n855), .ZN(new_n913));
  INV_X1    g727(.A(new_n768), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n319), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT118), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n897), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n896), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(KEYINPUT119), .B(new_n896), .C1(new_n912), .C2(new_n919), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(G54));
  NAND3_X1  g738(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n636), .Z(new_n926));
  INV_X1    g740(.A(new_n896), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(G60));
  XNOR2_X1  g742(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n496), .A2(new_n462), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n613), .A2(new_n617), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n909), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n909), .B2(new_n931), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n927), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n913), .A2(new_n647), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n595), .B1(new_n913), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n927), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n939), .B(new_n941), .C1(new_n942), .C2(KEYINPUT61), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT61), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n283), .B1(new_n383), .B2(new_n282), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n832), .A2(new_n818), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n283), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n902), .B1(G898), .B2(new_n283), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n948), .B(new_n949), .Z(G69));
  NOR2_X1   g764(.A1(new_n517), .A2(new_n519), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n409), .A2(new_n411), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n801), .A2(new_n728), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n683), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n961));
  INV_X1    g775(.A(new_n620), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n465), .B2(new_n640), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n379), .A2(new_n680), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n963), .A2(new_n602), .A3(new_n964), .A4(new_n776), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n778), .A2(new_n788), .A3(new_n961), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n955), .B1(new_n967), .B2(new_n283), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n774), .A2(new_n763), .A3(new_n846), .A4(new_n802), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n788), .B(new_n970), .C1(new_n775), .C2(new_n777), .ZN(new_n971));
  OR3_X1    g785(.A1(new_n748), .A2(new_n750), .A3(new_n956), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n283), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n659), .A2(G953), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n973), .A2(KEYINPUT125), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(KEYINPUT125), .B1(new_n973), .B2(new_n974), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n954), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI221_X1 g793(.A(G953), .B1(new_n323), .B2(new_n659), .C1(new_n954), .C2(KEYINPUT126), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n969), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n968), .B2(new_n978), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n967), .B2(new_n947), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n550), .A2(new_n551), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n987), .A2(new_n511), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n971), .A2(new_n972), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n986), .B1(new_n991), .B2(new_n947), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n511), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n994), .B(new_n988), .C1(new_n993), .C2(new_n992), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n913), .A2(new_n986), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n552), .A2(new_n523), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n927), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n990), .A2(new_n995), .A3(new_n998), .ZN(G57));
endmodule


