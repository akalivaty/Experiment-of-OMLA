

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U556 ( .A1(n680), .A2(n679), .ZN(n727) );
  INV_X1 U557 ( .A(n729), .ZN(n705) );
  NOR2_X1 U558 ( .A1(n811), .A2(n810), .ZN(n813) );
  XNOR2_X1 U559 ( .A(KEYINPUT29), .B(n520), .ZN(n719) );
  AND2_X1 U560 ( .A1(n718), .A2(n717), .ZN(n520) );
  XNOR2_X1 U561 ( .A(n690), .B(n689), .ZN(n735) );
  XNOR2_X1 U562 ( .A(KEYINPUT31), .B(KEYINPUT91), .ZN(n689) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n774) );
  INV_X1 U564 ( .A(KEYINPUT96), .ZN(n812) );
  NOR2_X1 U565 ( .A1(G651), .A2(n629), .ZN(n647) );
  NOR2_X1 U566 ( .A1(n530), .A2(n529), .ZN(G160) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n521), .Z(n887) );
  NAND2_X1 U569 ( .A1(n887), .A2(G137), .ZN(n524) );
  INV_X1 U570 ( .A(G2104), .ZN(n525) );
  NOR2_X2 U571 ( .A1(G2105), .A2(n525), .ZN(n894) );
  NAND2_X1 U572 ( .A1(G101), .A2(n894), .ZN(n522) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  NAND2_X1 U574 ( .A1(n524), .A2(n523), .ZN(n530) );
  INV_X1 U575 ( .A(G2105), .ZN(n526) );
  NOR2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n888) );
  NAND2_X1 U577 ( .A1(G113), .A2(n888), .ZN(n528) );
  NOR2_X1 U578 ( .A1(n526), .A2(G2104), .ZN(n889) );
  NAND2_X1 U579 ( .A1(G125), .A2(n889), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U581 ( .A1(G114), .A2(n888), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G126), .A2(n889), .ZN(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U584 ( .A(KEYINPUT80), .B(n533), .ZN(n538) );
  NAND2_X1 U585 ( .A1(G138), .A2(n887), .ZN(n535) );
  NAND2_X1 U586 ( .A1(G102), .A2(n894), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U588 ( .A(KEYINPUT81), .B(n536), .Z(n537) );
  NOR2_X1 U589 ( .A1(n538), .A2(n537), .ZN(G164) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U591 ( .A1(G135), .A2(n887), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G111), .A2(n888), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n889), .A2(G123), .ZN(n541) );
  XOR2_X1 U595 ( .A(KEYINPUT18), .B(n541), .Z(n542) );
  NOR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n894), .A2(G99), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n939) );
  XNOR2_X1 U599 ( .A(G2096), .B(n939), .ZN(n546) );
  OR2_X1 U600 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  XOR2_X1 U604 ( .A(G543), .B(KEYINPUT0), .Z(n629) );
  NAND2_X1 U605 ( .A1(G52), .A2(n647), .ZN(n549) );
  INV_X1 U606 ( .A(G651), .ZN(n550) );
  NOR2_X1 U607 ( .A1(G543), .A2(n550), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT1), .B(n547), .Z(n640) );
  NAND2_X1 U609 ( .A1(G64), .A2(n640), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n556) );
  NOR2_X1 U611 ( .A1(G543), .A2(G651), .ZN(n639) );
  NAND2_X1 U612 ( .A1(G90), .A2(n639), .ZN(n552) );
  NOR2_X1 U613 ( .A1(n629), .A2(n550), .ZN(n643) );
  NAND2_X1 U614 ( .A1(G77), .A2(n643), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT66), .B(n554), .ZN(n555) );
  NOR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  NAND2_X1 U620 ( .A1(G53), .A2(n647), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G65), .A2(n640), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G91), .A2(n639), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G78), .A2(n643), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n698) );
  INV_X1 U627 ( .A(n698), .ZN(G299) );
  NAND2_X1 U628 ( .A1(n639), .A2(G89), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G76), .A2(n643), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G51), .A2(n647), .ZN(n568) );
  NAND2_X1 U634 ( .A1(G63), .A2(n640), .ZN(n567) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U639 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n832) );
  NAND2_X1 U643 ( .A1(n832), .A2(G567), .ZN(n574) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U645 ( .A1(G56), .A2(n640), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n575), .Z(n582) );
  NAND2_X1 U647 ( .A1(n643), .A2(G68), .ZN(n576) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(n576), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n639), .A2(G81), .ZN(n577) );
  XOR2_X1 U650 ( .A(KEYINPUT12), .B(n577), .Z(n578) );
  NOR2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U652 ( .A(n580), .B(KEYINPUT13), .ZN(n581) );
  NOR2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n647), .A2(G43), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n584), .A2(n583), .ZN(n988) );
  INV_X1 U656 ( .A(n988), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n585), .A2(G860), .ZN(G153) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U659 ( .A1(n647), .A2(G54), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G79), .A2(n643), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G66), .A2(n640), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n639), .A2(G92), .ZN(n588) );
  XOR2_X1 U664 ( .A(KEYINPUT68), .B(n588), .Z(n589) );
  NOR2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U667 ( .A(KEYINPUT15), .B(n593), .Z(n993) );
  INV_X1 U668 ( .A(G868), .ZN(n659) );
  NAND2_X1 U669 ( .A1(n993), .A2(n659), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(G284) );
  NOR2_X1 U671 ( .A1(G286), .A2(n659), .ZN(n597) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n597), .A2(n596), .ZN(G297) );
  INV_X1 U674 ( .A(G559), .ZN(n598) );
  NOR2_X1 U675 ( .A1(G860), .A2(n598), .ZN(n599) );
  XNOR2_X1 U676 ( .A(KEYINPUT69), .B(n599), .ZN(n600) );
  INV_X1 U677 ( .A(n993), .ZN(n615) );
  NAND2_X1 U678 ( .A1(n600), .A2(n615), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(n993), .A2(n659), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT70), .B(n602), .Z(n603) );
  NOR2_X1 U682 ( .A1(G559), .A2(n603), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT71), .B(n604), .Z(n606) );
  NOR2_X1 U684 ( .A1(G868), .A2(n988), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U686 ( .A1(G67), .A2(n640), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT74), .ZN(n614) );
  NAND2_X1 U688 ( .A1(G93), .A2(n639), .ZN(n609) );
  NAND2_X1 U689 ( .A1(G55), .A2(n647), .ZN(n608) );
  NAND2_X1 U690 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U691 ( .A1(G80), .A2(n643), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT73), .B(n610), .ZN(n611) );
  NOR2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n660) );
  XNOR2_X1 U695 ( .A(n988), .B(KEYINPUT72), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n615), .A2(G559), .ZN(n616) );
  XNOR2_X1 U697 ( .A(n617), .B(n616), .ZN(n657) );
  NOR2_X1 U698 ( .A1(n657), .A2(G860), .ZN(n618) );
  XOR2_X1 U699 ( .A(n660), .B(n618), .Z(G145) );
  NAND2_X1 U700 ( .A1(G88), .A2(n639), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G75), .A2(n643), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U703 ( .A(KEYINPUT75), .B(n621), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n647), .A2(G50), .ZN(n623) );
  NAND2_X1 U705 ( .A1(G62), .A2(n640), .ZN(n622) );
  AND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(G303) );
  INV_X1 U708 ( .A(G303), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G49), .A2(n647), .ZN(n627) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U711 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U712 ( .A1(n640), .A2(n628), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G85), .A2(n639), .ZN(n633) );
  NAND2_X1 U716 ( .A1(G72), .A2(n643), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G60), .A2(n640), .ZN(n634) );
  XNOR2_X1 U719 ( .A(KEYINPUT65), .B(n634), .ZN(n635) );
  NOR2_X1 U720 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n647), .A2(G47), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(G290) );
  NAND2_X1 U723 ( .A1(G86), .A2(n639), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G61), .A2(n640), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n647), .A2(G48), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT77), .ZN(n651) );
  XNOR2_X1 U732 ( .A(G288), .B(KEYINPUT76), .ZN(n650) );
  XNOR2_X1 U733 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U734 ( .A(G166), .B(n652), .ZN(n654) );
  XNOR2_X1 U735 ( .A(G290), .B(n698), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n655), .B(G305), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(n660), .ZN(n906) );
  XNOR2_X1 U739 ( .A(n657), .B(n906), .ZN(n658) );
  NOR2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U741 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U742 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(KEYINPUT78), .B(n663), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U746 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U752 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(G96), .A2(n670), .ZN(n836) );
  NAND2_X1 U754 ( .A1(n836), .A2(G2106), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U756 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G108), .A2(n672), .ZN(n837) );
  NAND2_X1 U758 ( .A1(n837), .A2(G567), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n838) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n838), .A2(n675), .ZN(n676) );
  XOR2_X1 U762 ( .A(KEYINPUT79), .B(n676), .Z(n835) );
  NAND2_X1 U763 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n773) );
  INV_X1 U765 ( .A(n773), .ZN(n677) );
  NAND2_X2 U766 ( .A1(n677), .A2(n774), .ZN(n729) );
  NAND2_X1 U767 ( .A1(n729), .A2(G8), .ZN(n678) );
  OR2_X1 U768 ( .A1(n678), .A2(KEYINPUT88), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n678), .A2(KEYINPUT88), .ZN(n679) );
  NOR2_X1 U770 ( .A1(n727), .A2(G1966), .ZN(n722) );
  NOR2_X1 U771 ( .A1(G2084), .A2(n729), .ZN(n723) );
  NOR2_X1 U772 ( .A1(n722), .A2(n723), .ZN(n681) );
  NAND2_X1 U773 ( .A1(G8), .A2(n681), .ZN(n682) );
  XNOR2_X1 U774 ( .A(n682), .B(KEYINPUT30), .ZN(n683) );
  NOR2_X1 U775 ( .A1(G168), .A2(n683), .ZN(n688) );
  XOR2_X1 U776 ( .A(G2078), .B(KEYINPUT25), .Z(n966) );
  NOR2_X1 U777 ( .A1(n966), .A2(n729), .ZN(n684) );
  XNOR2_X1 U778 ( .A(n684), .B(KEYINPUT89), .ZN(n686) );
  OR2_X1 U779 ( .A1(G1961), .A2(n705), .ZN(n685) );
  NAND2_X1 U780 ( .A1(n686), .A2(n685), .ZN(n691) );
  NOR2_X1 U781 ( .A1(G171), .A2(n691), .ZN(n687) );
  NOR2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(G171), .ZN(n720) );
  NAND2_X1 U784 ( .A1(n705), .A2(G2072), .ZN(n692) );
  XNOR2_X1 U785 ( .A(n692), .B(KEYINPUT27), .ZN(n694) );
  AND2_X1 U786 ( .A1(G1956), .A2(n729), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n696) );
  XOR2_X1 U789 ( .A(KEYINPUT28), .B(KEYINPUT90), .Z(n695) );
  XNOR2_X1 U790 ( .A(n696), .B(n695), .ZN(n718) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n716) );
  XNOR2_X1 U792 ( .A(KEYINPUT64), .B(KEYINPUT26), .ZN(n706) );
  NOR2_X1 U793 ( .A1(G1996), .A2(n706), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n699), .A2(n988), .ZN(n703) );
  NAND2_X1 U795 ( .A1(G1348), .A2(n729), .ZN(n701) );
  NAND2_X1 U796 ( .A1(n705), .A2(G2067), .ZN(n700) );
  NAND2_X1 U797 ( .A1(n701), .A2(n700), .ZN(n712) );
  NAND2_X1 U798 ( .A1(n993), .A2(n712), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n711) );
  INV_X1 U800 ( .A(G1341), .ZN(n1018) );
  NAND2_X1 U801 ( .A1(n1018), .A2(n706), .ZN(n704) );
  NAND2_X1 U802 ( .A1(n704), .A2(n729), .ZN(n709) );
  AND2_X1 U803 ( .A1(n705), .A2(G1996), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n712), .A2(n993), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n733) );
  AND2_X1 U811 ( .A1(n735), .A2(n733), .ZN(n721) );
  NOR2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n725) );
  NAND2_X1 U813 ( .A1(G8), .A2(n723), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U815 ( .A(n726), .B(KEYINPUT92), .ZN(n743) );
  INV_X1 U816 ( .A(n727), .ZN(n804) );
  NOR2_X1 U817 ( .A1(n727), .A2(G1971), .ZN(n728) );
  XNOR2_X1 U818 ( .A(KEYINPUT93), .B(n728), .ZN(n732) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U820 ( .A1(G166), .A2(n730), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n736) );
  AND2_X1 U822 ( .A1(n733), .A2(n736), .ZN(n734) );
  NAND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n739) );
  INV_X1 U824 ( .A(n736), .ZN(n737) );
  OR2_X1 U825 ( .A1(n737), .A2(G286), .ZN(n738) );
  AND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U828 ( .A(n741), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n743), .A2(n742), .ZN(n803) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n750), .A2(n744), .ZN(n987) );
  NAND2_X1 U833 ( .A1(n803), .A2(n987), .ZN(n747) );
  INV_X1 U834 ( .A(n747), .ZN(n746) );
  INV_X1 U835 ( .A(KEYINPUT94), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U837 ( .A1(KEYINPUT94), .A2(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n755) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n991) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n750), .A2(n804), .ZN(n751) );
  NOR2_X1 U842 ( .A1(n757), .A2(n751), .ZN(n752) );
  XNOR2_X1 U843 ( .A(n752), .B(KEYINPUT95), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n991), .A2(n756), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n727), .A2(n753), .ZN(n754) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n760) );
  INV_X1 U847 ( .A(n756), .ZN(n758) );
  OR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  AND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n797) );
  XNOR2_X1 U850 ( .A(G1981), .B(G305), .ZN(n984) );
  XNOR2_X1 U851 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n764) );
  NAND2_X1 U852 ( .A1(G116), .A2(n888), .ZN(n762) );
  NAND2_X1 U853 ( .A1(G128), .A2(n889), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n764), .B(n763), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n887), .A2(G140), .ZN(n765) );
  XNOR2_X1 U857 ( .A(n765), .B(KEYINPUT82), .ZN(n767) );
  NAND2_X1 U858 ( .A1(G104), .A2(n894), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n768), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U862 ( .A(n771), .B(KEYINPUT36), .ZN(n772) );
  XNOR2_X1 U863 ( .A(n772), .B(KEYINPUT84), .ZN(n903) );
  XNOR2_X1 U864 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U865 ( .A1(n903), .A2(n824), .ZN(n941) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n826) );
  NAND2_X1 U867 ( .A1(n941), .A2(n826), .ZN(n775) );
  XOR2_X1 U868 ( .A(KEYINPUT85), .B(n775), .Z(n823) );
  NAND2_X1 U869 ( .A1(G141), .A2(n887), .ZN(n777) );
  NAND2_X1 U870 ( .A1(G117), .A2(n888), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n894), .A2(G105), .ZN(n778) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n889), .A2(G129), .ZN(n781) );
  NAND2_X1 U876 ( .A1(n782), .A2(n781), .ZN(n870) );
  NAND2_X1 U877 ( .A1(G1996), .A2(n870), .ZN(n783) );
  XNOR2_X1 U878 ( .A(n783), .B(KEYINPUT87), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G107), .A2(n888), .ZN(n785) );
  NAND2_X1 U880 ( .A1(G119), .A2(n889), .ZN(n784) );
  NAND2_X1 U881 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U882 ( .A(KEYINPUT86), .B(n786), .Z(n790) );
  NAND2_X1 U883 ( .A1(n894), .A2(G95), .ZN(n788) );
  NAND2_X1 U884 ( .A1(G131), .A2(n887), .ZN(n787) );
  AND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n869) );
  AND2_X1 U887 ( .A1(G1991), .A2(n869), .ZN(n791) );
  NOR2_X1 U888 ( .A1(n792), .A2(n791), .ZN(n936) );
  INV_X1 U889 ( .A(n826), .ZN(n793) );
  NOR2_X1 U890 ( .A1(n936), .A2(n793), .ZN(n818) );
  INV_X1 U891 ( .A(n818), .ZN(n794) );
  AND2_X1 U892 ( .A1(n823), .A2(n794), .ZN(n809) );
  INV_X1 U893 ( .A(n809), .ZN(n795) );
  OR2_X1 U894 ( .A1(n984), .A2(n795), .ZN(n796) );
  NOR2_X1 U895 ( .A1(n797), .A2(n796), .ZN(n811) );
  NOR2_X1 U896 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U897 ( .A1(G8), .A2(n798), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n799) );
  XOR2_X1 U899 ( .A(n799), .B(KEYINPUT24), .Z(n800) );
  OR2_X1 U900 ( .A1(n727), .A2(n800), .ZN(n805) );
  AND2_X1 U901 ( .A1(n801), .A2(n805), .ZN(n802) );
  AND2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n807) );
  AND2_X1 U903 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U904 ( .A1(n807), .A2(n806), .ZN(n808) );
  AND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U906 ( .A(n813), .B(n812), .ZN(n815) );
  XNOR2_X1 U907 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U908 ( .A1(n826), .A2(n990), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n830) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n870), .ZN(n933) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n869), .ZN(n938) );
  NOR2_X1 U913 ( .A1(n816), .A2(n938), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n933), .A2(n819), .ZN(n820) );
  XOR2_X1 U916 ( .A(n820), .B(KEYINPUT39), .Z(n821) );
  XNOR2_X1 U917 ( .A(KEYINPUT97), .B(n821), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n903), .A2(n824), .ZN(n935) );
  NAND2_X1 U920 ( .A1(n825), .A2(n935), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT98), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U924 ( .A(KEYINPUT40), .B(n831), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U927 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(G188) );
  NOR2_X1 U930 ( .A1(n837), .A2(n836), .ZN(G325) );
  XOR2_X1 U931 ( .A(KEYINPUT102), .B(G325), .Z(G261) );
  INV_X1 U932 ( .A(n838), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U934 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U937 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1976), .B(G1971), .Z(n848) );
  XNOR2_X1 U943 ( .A(G1986), .B(G1961), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n858) );
  XOR2_X1 U945 ( .A(KEYINPUT103), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1996), .B(KEYINPUT104), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(G1991), .B(G1956), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1981), .B(G1966), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U952 ( .A(KEYINPUT105), .B(G2474), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U954 ( .A(n858), .B(n857), .Z(G229) );
  NAND2_X1 U955 ( .A1(G100), .A2(n894), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G112), .A2(n888), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n868) );
  XOR2_X1 U958 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n862) );
  NAND2_X1 U959 ( .A1(G124), .A2(n889), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n865) );
  NAND2_X1 U961 ( .A1(n887), .A2(G136), .ZN(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT107), .B(n863), .ZN(n864) );
  NOR2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(KEYINPUT108), .B(n866), .Z(n867) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(G162) );
  XNOR2_X1 U966 ( .A(G160), .B(n869), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(n875) );
  XNOR2_X1 U968 ( .A(KEYINPUT109), .B(KEYINPUT113), .ZN(n873) );
  XNOR2_X1 U969 ( .A(n939), .B(KEYINPUT48), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U971 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U972 ( .A(G164), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U973 ( .A(n877), .B(n876), .ZN(n886) );
  NAND2_X1 U974 ( .A1(G118), .A2(n888), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G130), .A2(n889), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G106), .A2(n894), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G142), .A2(n887), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n882), .Z(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(n886), .B(n885), .Z(n902) );
  NAND2_X1 U983 ( .A1(G139), .A2(n887), .ZN(n899) );
  XNOR2_X1 U984 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n893) );
  NAND2_X1 U985 ( .A1(G115), .A2(n888), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G127), .A2(n889), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n897) );
  NAND2_X1 U989 ( .A1(n894), .A2(G103), .ZN(n895) );
  XOR2_X1 U990 ( .A(KEYINPUT110), .B(n895), .Z(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n900), .B(KEYINPUT112), .ZN(n948) );
  XNOR2_X1 U994 ( .A(n948), .B(G162), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U998 ( .A(G286), .B(n906), .ZN(n909) );
  XNOR2_X1 U999 ( .A(KEYINPUT114), .B(G301), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n907), .B(n993), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1002 ( .A(n910), .B(n988), .Z(n911) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n911), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2443), .B(KEYINPUT100), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2451), .B(G2427), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1007 ( .A(n914), .B(KEYINPUT101), .Z(n916) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n916), .B(n915), .ZN(n920) );
  XOR2_X1 U1010 ( .A(G2435), .B(G2438), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G2454), .B(G2430), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1013 ( .A(n920), .B(n919), .Z(n922) );
  XNOR2_X1 U1014 ( .A(G2446), .B(KEYINPUT99), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n923), .A2(G14), .ZN(n931) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n931), .ZN(n928) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G227), .A2(G229), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(n925), .B(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT115), .B(n926), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1024 ( .A1(n930), .A2(n929), .ZN(G225) );
  XNOR2_X1 U1025 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G120), .ZN(G236) );
  INV_X1 U1028 ( .A(G96), .ZN(G221) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  INV_X1 U1031 ( .A(n931), .ZN(G401) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n934), .Z(n947) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n945) );
  XOR2_X1 U1036 ( .A(G2084), .B(G160), .Z(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1040 ( .A(KEYINPUT118), .B(n943), .Z(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n953) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n950) );
  XNOR2_X1 U1044 ( .A(G2072), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1046 ( .A(KEYINPUT50), .B(n951), .Z(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n954), .ZN(n956) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n957), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1052 ( .A(G29), .B(KEYINPUT123), .ZN(n980) );
  XNOR2_X1 U1053 ( .A(G2084), .B(G34), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(n958), .B(KEYINPUT54), .ZN(n976) );
  XNOR2_X1 U1055 ( .A(G2090), .B(G35), .ZN(n973) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n959) );
  NAND2_X1 U1057 ( .A1(n959), .A2(G28), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(n960), .B(KEYINPUT119), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G32), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(G2072), .B(G33), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n970) );
  XOR2_X1 U1063 ( .A(G2067), .B(G26), .Z(n968) );
  XOR2_X1 U1064 ( .A(G27), .B(KEYINPUT120), .Z(n965) );
  XNOR2_X1 U1065 ( .A(n966), .B(n965), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(KEYINPUT121), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(KEYINPUT55), .B(n977), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT122), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n981), .A2(G11), .ZN(n1035) );
  INV_X1 U1076 ( .A(G16), .ZN(n1031) );
  XOR2_X1 U1077 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n982) );
  XNOR2_X1 U1078 ( .A(n1031), .B(n982), .ZN(n1007) );
  XOR2_X1 U1079 ( .A(G1966), .B(G168), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1081 ( .A(KEYINPUT57), .B(n985), .Z(n1005) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(n1018), .B(n988), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G299), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n992), .A2(n991), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(G301), .B(G1961), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n993), .B(G1348), .ZN(n994) );
  NOR2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(n996), .B(KEYINPUT125), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1003), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1033) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(G1986), .B(G24), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1008) );
  NOR2_X1 U1101 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(n1013), .B(n1012), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1014) );
  NOR2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1028) );
  XNOR2_X1 U1109 ( .A(G19), .B(n1018), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G1981), .B(G6), .ZN(n1020) );
  XNOR2_X1 U1111 ( .A(G1956), .B(G20), .ZN(n1019) );
  NOR2_X1 U1112 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1113 ( .A1(n1022), .A2(n1021), .ZN(n1025) );
  XOR2_X1 U1114 ( .A(KEYINPUT59), .B(G1348), .Z(n1023) );
  XNOR2_X1 U1115 ( .A(G4), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1116 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1117 ( .A(KEYINPUT60), .B(n1026), .Z(n1027) );
  NOR2_X1 U1118 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1119 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

