//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1232, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  AOI22_X1  g0008(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n217), .A2(new_n218), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n225), .B1(new_n218), .B2(new_n217), .C1(new_n213), .C2(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n215), .A2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT2), .ZN(new_n229));
  INV_X1    g0029(.A(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G1), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G274), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT66), .B(G45), .ZN(new_n246));
  INV_X1    g0046(.A(G41), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n249));
  OR2_X1    g0049(.A1(KEYINPUT67), .A2(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT67), .A2(G1), .ZN(new_n251));
  AND2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n249), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(G226), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G77), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n257), .A2(G1698), .ZN(new_n261));
  INV_X1    g0061(.A(G223), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n259), .B1(new_n260), .B2(new_n257), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI211_X1 g0063(.A(new_n248), .B(new_n256), .C1(new_n263), .C2(new_n249), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G179), .ZN(new_n265));
  INV_X1    g0065(.A(G169), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n264), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT8), .A2(G58), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT68), .B(G58), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT8), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n223), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n222), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n252), .B2(G20), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G50), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n250), .A2(G13), .A3(G20), .A4(new_n251), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n279), .B(new_n281), .C1(G50), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n267), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT69), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n283), .B(KEYINPUT9), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n264), .A2(G190), .ZN(new_n287));
  INV_X1    g0087(.A(G200), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n264), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT10), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n257), .A2(G232), .A3(new_n258), .ZN(new_n291));
  INV_X1    g0091(.A(G107), .ZN(new_n292));
  INV_X1    g0092(.A(G238), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n291), .B1(new_n292), .B2(new_n257), .C1(new_n261), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n249), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n248), .B1(new_n255), .B2(G244), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G179), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n266), .B2(new_n297), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n280), .A2(G77), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT70), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n300), .B(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT8), .B(G58), .Z(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n268), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT15), .B(G87), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(new_n223), .B2(new_n260), .C1(new_n275), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n282), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n306), .A2(new_n278), .B1(new_n260), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n299), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT71), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n309), .B(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n297), .A2(new_n288), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(G190), .B2(new_n297), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n311), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n285), .A2(new_n290), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n274), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n280), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n274), .A2(new_n307), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n219), .B1(new_n272), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G20), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n268), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT74), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n335), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n223), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n223), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT75), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n337), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT16), .B(new_n328), .C1(new_n343), .C2(new_n323), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT16), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n339), .B1(new_n257), .B2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n332), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n323), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n327), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n278), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n322), .B1(new_n344), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n248), .B1(new_n255), .B2(G232), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G226), .A2(G1698), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n262), .B2(G1698), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n357), .A2(new_n330), .A3(new_n333), .A4(new_n334), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT76), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n249), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n266), .ZN(new_n365));
  INV_X1    g0165(.A(G179), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n355), .B(new_n366), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT18), .B1(new_n354), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n364), .A2(new_n288), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n355), .B(new_n371), .C1(new_n362), .C2(new_n363), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n354), .A2(KEYINPUT17), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n335), .B2(new_n223), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n342), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n323), .B1(new_n377), .B2(new_n336), .ZN(new_n378));
  NOR3_X1   g0178(.A1(new_n378), .A2(new_n345), .A3(new_n327), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n321), .B1(new_n379), .B2(new_n352), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT18), .ZN(new_n381));
  INV_X1    g0181(.A(new_n368), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n373), .B(new_n321), .C1(new_n379), .C2(new_n352), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT17), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n369), .A2(new_n374), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n248), .B1(new_n255), .B2(G238), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n257), .A2(G226), .A3(new_n258), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n257), .A2(G232), .A3(G1698), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n249), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n388), .B2(new_n393), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n398), .A2(KEYINPUT14), .A3(new_n266), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT14), .B1(new_n398), .B2(new_n266), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n395), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n399), .B(new_n400), .C1(new_n366), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT12), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n280), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n307), .A2(KEYINPUT12), .A3(new_n323), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(KEYINPUT12), .C2(new_n307), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n268), .A2(G50), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n223), .B2(G68), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n275), .A2(new_n260), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n278), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT73), .B(KEYINPUT11), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n403), .A2(new_n371), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n415), .B1(new_n398), .B2(new_n288), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n317), .A2(new_n387), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n278), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT23), .B1(new_n223), .B2(G107), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT23), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(new_n292), .A3(G20), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G116), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n425), .B(new_n427), .C1(G20), .C2(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n330), .A2(new_n333), .A3(new_n223), .A4(new_n334), .ZN(new_n432));
  INV_X1    g0232(.A(G87), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT22), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT85), .B(KEYINPUT22), .Z(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(new_n223), .A3(G87), .A4(new_n257), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n430), .A2(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n424), .B1(new_n437), .B2(KEYINPUT24), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(KEYINPUT24), .B2(new_n437), .ZN(new_n439));
  INV_X1    g0239(.A(G250), .ZN(new_n440));
  INV_X1    g0240(.A(G257), .ZN(new_n441));
  MUX2_X1   g0241(.A(new_n440), .B(new_n441), .S(G1698), .Z(new_n442));
  INV_X1    g0242(.A(G294), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n335), .A2(new_n442), .B1(new_n329), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n249), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT67), .B(G1), .ZN(new_n447));
  OAI21_X1  g0247(.A(G45), .B1(new_n247), .B2(KEYINPUT5), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n253), .B1(new_n450), .B2(G41), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT77), .A3(new_n250), .A4(new_n251), .ZN(new_n452));
  OAI21_X1  g0252(.A(G274), .B1(new_n450), .B2(G41), .ZN(new_n453));
  INV_X1    g0253(.A(new_n222), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G41), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G264), .ZN(new_n458));
  INV_X1    g0258(.A(new_n249), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n450), .A2(G41), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n250), .A2(new_n460), .A3(G45), .A4(new_n251), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n450), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n445), .B(new_n457), .C1(new_n458), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n288), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G190), .B2(new_n464), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n282), .B(new_n424), .C1(new_n329), .C2(new_n447), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n292), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n282), .A2(KEYINPUT25), .A3(G107), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT25), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n307), .B2(new_n292), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n468), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n439), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n463), .A2(new_n458), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n249), .B2(new_n444), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G179), .A3(new_n457), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n464), .A2(G169), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n439), .A2(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT87), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n439), .A2(new_n472), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT87), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n439), .A2(new_n466), .A3(new_n472), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n293), .A2(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n330), .A2(new_n333), .A3(new_n334), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT81), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n330), .A2(new_n333), .A3(G244), .A4(new_n334), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n258), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n428), .B1(new_n488), .B2(KEYINPUT81), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n249), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n447), .A2(new_n253), .A3(G274), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n447), .A2(new_n253), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n494), .B(new_n459), .C1(G250), .C2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n366), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n223), .B1(new_n391), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G87), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n292), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n223), .A2(G33), .A3(G97), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n501), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n323), .B2(new_n432), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n278), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n307), .A2(new_n305), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n305), .B(KEYINPUT82), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n506), .C1(new_n467), .C2(new_n507), .ZN(new_n508));
  AND4_X1   g0308(.A1(G244), .A2(new_n330), .A3(new_n333), .A4(new_n334), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(G1698), .B1(KEYINPUT81), .B2(new_n488), .ZN(new_n510));
  INV_X1    g0310(.A(new_n492), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n459), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n496), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n497), .B(new_n508), .C1(new_n514), .C2(G169), .ZN(new_n515));
  OAI21_X1  g0315(.A(G200), .B1(new_n512), .B2(new_n513), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n493), .A2(G190), .A3(new_n496), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n505), .A2(new_n506), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n467), .A2(new_n433), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n459), .B(G257), .C1(new_n461), .C2(new_n462), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n457), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n523), .B1(new_n457), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT79), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n457), .A2(new_n524), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT78), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT79), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n457), .A2(new_n523), .A3(new_n524), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT4), .B1(new_n509), .B2(new_n258), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n249), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n527), .A2(new_n532), .A3(new_n366), .A4(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G97), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n282), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(G97), .B2(new_n467), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT7), .B1(new_n348), .B2(new_n223), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n339), .B(G20), .C1(new_n347), .C2(new_n334), .ZN(new_n544));
  OAI21_X1  g0344(.A(G107), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n292), .A2(KEYINPUT6), .A3(G97), .ZN(new_n546));
  AND2_X1   g0346(.A1(G97), .A2(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(KEYINPUT6), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n545), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n542), .B1(new_n552), .B2(new_n278), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n529), .A2(new_n538), .A3(new_n531), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(new_n266), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n539), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n522), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n527), .A2(new_n532), .A3(new_n538), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(G200), .ZN(new_n559));
  INV_X1    g0359(.A(new_n553), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n529), .A2(new_n538), .A3(new_n531), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(G190), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT80), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n559), .A2(new_n562), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT80), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n557), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n329), .A2(G97), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(new_n569), .B2(new_n536), .ZN(new_n570));
  INV_X1    g0370(.A(G116), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n223), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n278), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT20), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n307), .A2(new_n571), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n467), .B2(new_n571), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  MUX2_X1   g0377(.A(new_n441), .B(new_n458), .S(G1698), .Z(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n335), .A2(new_n578), .B1(new_n579), .B2(new_n257), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n249), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n459), .B(G270), .C1(new_n461), .C2(new_n462), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(G179), .A3(new_n457), .A4(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n568), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n576), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  XNOR2_X1  g0386(.A(new_n573), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n583), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT83), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(new_n457), .A3(new_n582), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n288), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G190), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n577), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(G169), .A3(new_n592), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n266), .B1(new_n585), .B2(new_n587), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(KEYINPUT21), .A3(new_n592), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n591), .A2(new_n595), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n599), .A2(KEYINPUT21), .A3(new_n592), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT21), .B1(new_n599), .B2(new_n592), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n591), .A4(new_n595), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n423), .A2(new_n486), .A3(new_n567), .A4(new_n608), .ZN(G372));
  INV_X1    g0409(.A(new_n515), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n515), .A2(new_n521), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n611), .A2(new_n556), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n613), .B2(KEYINPUT26), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT26), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n539), .A2(new_n555), .A3(KEYINPUT88), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT88), .B1(new_n539), .B2(new_n555), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n615), .B(new_n522), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n539), .A2(new_n555), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n563), .B1(new_n559), .B2(new_n562), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n591), .A2(new_n600), .A3(new_n598), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n484), .B1(new_n624), .B2(new_n478), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n614), .B(new_n618), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n423), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n285), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n369), .A2(new_n383), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n421), .A2(new_n311), .B1(new_n404), .B2(new_n416), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n374), .A2(new_n386), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n633), .B2(new_n290), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n627), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(G13), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(G20), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n252), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n577), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n608), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n624), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(KEYINPUT89), .B(G330), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n480), .A2(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n486), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT90), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT90), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n478), .A2(new_n643), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n647), .A2(new_n643), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n657), .A2(new_n662), .B1(new_n478), .B2(new_n644), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n216), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G1), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n500), .A2(new_n292), .A3(new_n571), .ZN(new_n669));
  OAI22_X1  g0469(.A1(new_n668), .A2(new_n669), .B1(new_n220), .B2(new_n667), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n514), .A2(new_n475), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT92), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT92), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n475), .A2(new_n493), .A3(new_n674), .A4(new_n496), .ZN(new_n675));
  NOR2_X1   g0475(.A1(KEYINPUT93), .A2(KEYINPUT30), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n554), .A2(new_n583), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(KEYINPUT93), .A2(KEYINPUT30), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n673), .A2(new_n675), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n583), .A2(new_n676), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n675), .A2(new_n561), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n674), .B1(new_n514), .B2(new_n475), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n464), .A2(new_n366), .A3(new_n592), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n558), .B(new_n685), .C1(new_n512), .C2(new_n513), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n680), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(KEYINPUT91), .B(KEYINPUT31), .Z(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n643), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n643), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n692), .B2(KEYINPUT31), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n567), .A2(new_n486), .A3(new_n608), .A4(new_n644), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n650), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n626), .A2(new_n644), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI211_X1 g0500(.A(KEYINPUT94), .B(KEYINPUT29), .C1(new_n626), .C2(new_n644), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n522), .B1(new_n616), .B2(new_n617), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT26), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n610), .B1(new_n612), .B2(new_n615), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n704), .B(new_n705), .C1(new_n623), .C2(new_n625), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n644), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n696), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n671), .B1(new_n708), .B2(G1), .ZN(G364));
  AOI21_X1  g0509(.A(new_n668), .B1(G45), .B2(new_n637), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n652), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n649), .A2(new_n651), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n636), .A2(new_n329), .A3(KEYINPUT96), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT96), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(G13), .B2(G33), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n223), .ZN(new_n719));
  XOR2_X1   g0519(.A(new_n719), .B(KEYINPUT97), .Z(new_n720));
  NOR2_X1   g0520(.A1(new_n649), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n720), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n222), .B1(G20), .B2(new_n266), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n246), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n220), .ZN(new_n726));
  INV_X1    g0526(.A(new_n335), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n665), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n726), .B(new_n729), .C1(new_n239), .C2(G45), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n665), .A2(new_n348), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n571), .B2(new_n665), .ZN(new_n732));
  XOR2_X1   g0532(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  OAI21_X1  g0533(.A(new_n724), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n223), .A2(G190), .ZN(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT99), .Z(new_n736));
  NOR3_X1   g0536(.A1(new_n736), .A2(G179), .A3(new_n288), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G107), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n736), .A2(G179), .A3(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G159), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT32), .Z(new_n745));
  NOR2_X1   g0545(.A1(new_n223), .A2(new_n371), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n366), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n272), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n366), .A2(new_n288), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n735), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n735), .A2(new_n747), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n323), .B1(new_n758), .B2(new_n260), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n223), .B1(new_n760), .B2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n746), .A2(new_n756), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n257), .B1(new_n761), .B2(new_n540), .C1(new_n762), .C2(new_n202), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n746), .A2(new_n366), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n759), .B(new_n763), .C1(G87), .C2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n742), .A2(new_n745), .A3(new_n755), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n741), .A2(G283), .ZN(new_n768));
  INV_X1    g0568(.A(new_n757), .ZN(new_n769));
  NOR2_X1   g0569(.A1(KEYINPUT33), .A2(G317), .ZN(new_n770));
  AND2_X1   g0570(.A1(KEYINPUT33), .A2(G317), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n579), .B2(new_n764), .ZN(new_n773));
  INV_X1    g0573(.A(new_n762), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(G326), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n761), .A2(new_n443), .ZN(new_n776));
  INV_X1    g0576(.A(new_n758), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n257), .B(new_n776), .C1(G311), .C2(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G322), .A2(new_n753), .B1(new_n743), .B2(G329), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n768), .A2(new_n775), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n767), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n723), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n734), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n710), .B1(new_n721), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n714), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n313), .A2(new_n315), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n309), .A2(new_n643), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT103), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n310), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n311), .A2(new_n644), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n698), .B(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n710), .B1(new_n794), .B2(new_n696), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n696), .B2(new_n794), .ZN(new_n796));
  INV_X1    g0596(.A(new_n718), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n782), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n710), .B1(G77), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n764), .A2(new_n292), .B1(new_n757), .B2(new_n800), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n348), .B1(new_n761), .B2(new_n540), .C1(new_n762), .C2(new_n579), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n801), .B(new_n802), .C1(G116), .C2(new_n777), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G294), .A2(new_n753), .B1(new_n743), .B2(G311), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(new_n740), .C2(new_n433), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G137), .A2(new_n774), .B1(new_n777), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G150), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n807), .B2(new_n757), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G143), .B2(new_n753), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT102), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n811));
  XNOR2_X1  g0611(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n741), .A2(G68), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n743), .A2(G132), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n727), .B1(new_n202), .B2(new_n764), .ZN(new_n815));
  INV_X1    g0615(.A(new_n761), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n754), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n805), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n799), .B1(new_n819), .B2(new_n723), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n793), .B2(new_n797), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n796), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(G384));
  OAI211_X1 g0623(.A(G116), .B(new_n224), .C1(new_n550), .C2(KEYINPUT35), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(KEYINPUT35), .B2(new_n550), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT36), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n221), .B(G77), .C1(new_n323), .C2(new_n272), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n202), .A2(G68), .ZN(new_n828));
  AOI211_X1 g0628(.A(G13), .B(new_n252), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT109), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT31), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n691), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n687), .A2(KEYINPUT109), .A3(KEYINPUT31), .A4(new_n643), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n695), .A2(new_n689), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n835), .B1(new_n836), .B2(new_n691), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n384), .B1(new_n354), .B2(new_n641), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n377), .A2(new_n336), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n327), .B1(new_n841), .B2(G68), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n352), .B1(new_n842), .B2(KEYINPUT16), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n382), .B1(new_n843), .B2(new_n322), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT37), .B1(new_n844), .B2(KEYINPUT106), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT106), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n382), .C1(new_n843), .C2(new_n322), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n840), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n641), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n380), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(new_n844), .A3(new_n384), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  INV_X1    g0652(.A(new_n850), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n848), .A2(new_n852), .B1(new_n387), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT108), .B1(new_n854), .B2(KEYINPUT38), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT108), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT38), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n847), .A2(new_n850), .A3(new_n384), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n859), .A2(new_n845), .B1(KEYINPUT37), .B2(new_n851), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n850), .B1(new_n629), .B2(new_n631), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n856), .B(new_n857), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(KEYINPUT105), .A2(KEYINPUT16), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n328), .B(new_n864), .C1(new_n343), .C2(new_n323), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n378), .B2(new_n327), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n278), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n641), .B1(new_n867), .B2(new_n321), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n387), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  INV_X1    g0670(.A(new_n384), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n368), .B1(new_n867), .B2(new_n321), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n870), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n344), .A2(new_n353), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n368), .B1(new_n876), .B2(new_n321), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n870), .B1(new_n877), .B2(new_n846), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n878), .A2(new_n858), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT38), .B(new_n869), .C1(new_n875), .C2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n855), .A2(new_n862), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n791), .A2(new_n792), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n417), .B(new_n421), .C1(new_n415), .C2(new_n644), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n416), .B(new_n643), .C1(new_n404), .C2(new_n420), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n838), .A2(new_n881), .A3(KEYINPUT40), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n692), .B1(new_n695), .B2(new_n689), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n835), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT107), .ZN(new_n889));
  INV_X1    g0689(.A(new_n880), .ZN(new_n890));
  NOR3_X1   g0690(.A1(new_n873), .A2(new_n868), .A3(new_n871), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n891), .A2(new_n870), .B1(new_n878), .B2(new_n858), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n892), .B2(new_n869), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n889), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n875), .A2(new_n879), .ZN(new_n895));
  INV_X1    g0695(.A(new_n869), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n857), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(KEYINPUT107), .A3(new_n880), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n888), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n886), .B1(new_n899), .B2(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n838), .A2(new_n423), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(new_n650), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n883), .A2(new_n884), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n626), .A2(new_n793), .A3(new_n644), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n792), .B(KEYINPUT104), .Z(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n890), .A2(new_n893), .A3(new_n889), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT107), .B1(new_n897), .B2(new_n880), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n629), .A2(new_n849), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n417), .A2(new_n643), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT39), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n855), .A2(new_n862), .A3(new_n916), .A4(new_n880), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT39), .B1(new_n890), .B2(new_n893), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n423), .B(new_n707), .C1(new_n700), .C2(new_n701), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n634), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n903), .A2(new_n923), .B1(new_n252), .B2(new_n637), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n903), .A2(new_n923), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n830), .B1(new_n924), .B2(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n658), .A2(new_n659), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT42), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n556), .B1(new_n553), .B2(new_n644), .C1(new_n621), .C2(new_n622), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n619), .A2(new_n643), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n662), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n927), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n556), .B1(new_n929), .B2(new_n482), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n644), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n928), .B1(new_n927), .B2(new_n934), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n643), .B1(new_n518), .B2(new_n519), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n515), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT110), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n522), .A2(new_n942), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n944), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT111), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n941), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n661), .A2(new_n932), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n941), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n953), .B(new_n954), .C1(new_n938), .C2(new_n939), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n951), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n952), .B1(new_n951), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n666), .B(KEYINPUT41), .Z(new_n959));
  INV_X1    g0759(.A(KEYINPUT113), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n660), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n931), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT45), .B1(new_n663), .B2(new_n931), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT112), .B(KEYINPUT44), .Z(new_n967));
  OR3_X1    g0767(.A1(new_n663), .A2(new_n931), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n663), .B2(new_n931), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n965), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n963), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n973), .A2(new_n968), .A3(new_n969), .A4(new_n961), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n658), .A2(new_n652), .A3(new_n659), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n661), .A2(new_n662), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n975), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n933), .B1(new_n977), .B2(new_n660), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n971), .A2(new_n974), .A3(new_n708), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n959), .B1(new_n980), .B2(new_n708), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n244), .B1(new_n637), .B2(G45), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n958), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n724), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n729), .A2(new_n235), .B1(new_n216), .B2(new_n305), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n711), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n741), .A2(G97), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n777), .A2(G283), .ZN(new_n990));
  XNOR2_X1  g0790(.A(KEYINPUT114), .B(G311), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n443), .B2(new_n757), .C1(new_n762), .C2(new_n991), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n727), .B(new_n992), .C1(G107), .C2(new_n816), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT115), .B1(new_n764), .B2(new_n571), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n743), .A2(G317), .B1(KEYINPUT46), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT46), .ZN(new_n996));
  INV_X1    g0796(.A(new_n994), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n753), .A2(G303), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n989), .A2(new_n993), .A3(new_n995), .A4(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n740), .A2(new_n260), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G150), .A2(new_n753), .B1(new_n743), .B2(G137), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n761), .A2(new_n323), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n348), .B(new_n1002), .C1(G143), .C2(new_n774), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n764), .A2(new_n272), .B1(new_n758), .B2(new_n202), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G159), .B2(new_n769), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n999), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT47), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n723), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .C1(new_n949), .C2(new_n720), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT116), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n984), .A2(new_n1012), .ZN(G387));
  NAND3_X1  g0813(.A1(new_n976), .A2(new_n978), .A3(new_n708), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(new_n666), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n708), .B2(new_n979), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n658), .A2(new_n659), .A3(new_n722), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n729), .B1(new_n232), .B2(new_n725), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n669), .B2(new_n731), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n303), .A2(new_n202), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n253), .B1(new_n323), .B2(new_n260), .ZN(new_n1022));
  NOR3_X1   g0822(.A1(new_n1021), .A2(new_n669), .A3(new_n1022), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n1019), .A2(new_n1023), .B1(G107), .B2(new_n216), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1024), .A2(new_n724), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n764), .A2(new_n260), .B1(new_n758), .B2(new_n323), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n335), .B(new_n1026), .C1(G159), .C2(new_n774), .ZN(new_n1027));
  XOR2_X1   g0827(.A(KEYINPUT117), .B(G150), .Z(new_n1028));
  INV_X1    g0828(.A(new_n507), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n743), .A2(new_n1028), .B1(new_n1029), .B2(new_n816), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n753), .A2(G50), .B1(new_n318), .B2(new_n769), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n989), .A2(new_n1027), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n727), .B1(new_n743), .B2(G326), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n764), .A2(new_n443), .B1(new_n761), .B2(new_n800), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n774), .A2(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n579), .B2(new_n758), .C1(new_n757), .C2(new_n991), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G317), .B2(new_n753), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1034), .B1(new_n1037), .B2(KEYINPUT48), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(KEYINPUT48), .B2(new_n1037), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1033), .B1(new_n571), .B2(new_n740), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1032), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n711), .B(new_n1025), .C1(new_n723), .C2(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n979), .A2(new_n983), .B1(new_n1017), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1016), .A2(new_n1045), .ZN(G393));
  OAI21_X1  g0846(.A(new_n661), .B1(new_n966), .B2(new_n970), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n973), .A2(new_n660), .A3(new_n968), .A4(new_n969), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n1014), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n980), .A2(new_n666), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n932), .A2(new_n722), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT118), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n242), .A2(new_n728), .B1(G97), .B2(new_n665), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n711), .B1(new_n724), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n753), .A2(G311), .B1(G317), .B2(new_n774), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n743), .A2(G322), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n816), .A2(G116), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n257), .B1(new_n765), .B2(G283), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n769), .B1(new_n777), .B2(G294), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n741), .B2(G107), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n743), .A2(G143), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n769), .A2(G50), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n765), .A2(G68), .B1(new_n777), .B2(new_n303), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n761), .A2(new_n260), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n335), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n741), .B2(G87), .ZN(new_n1069));
  INV_X1    g0869(.A(G159), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n752), .A2(new_n1070), .B1(new_n807), .B2(new_n762), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n1056), .A2(new_n1062), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1054), .B1(new_n1073), .B2(new_n782), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1052), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1075), .B1(new_n1076), .B2(new_n983), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1050), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  OAI211_X1 g0879(.A(new_n917), .B(new_n918), .C1(new_n907), .C2(new_n914), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n696), .A2(new_n885), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n706), .A2(new_n644), .A3(new_n791), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT119), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n792), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1082), .B2(new_n792), .ZN(new_n1086));
  NOR3_X1   g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n904), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n881), .A2(new_n915), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1080), .B(new_n1081), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n917), .A2(new_n918), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n905), .A2(new_n906), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n883), .A2(new_n884), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n915), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1082), .A2(new_n792), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n1093), .A3(new_n1084), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n867), .A2(new_n321), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n849), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n874), .A2(new_n1101), .A3(new_n384), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT37), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1103), .A2(new_n848), .B1(new_n387), .B2(new_n868), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1099), .A2(KEYINPUT108), .B1(new_n1104), .B2(KEYINPUT38), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n914), .B1(new_n1105), .B2(new_n862), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1091), .A2(new_n1095), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  AND3_X1   g0907(.A1(new_n791), .A2(G330), .A3(new_n792), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1093), .B(new_n1108), .C1(new_n887), .C2(new_n835), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1089), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1108), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n904), .B1(new_n837), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n1081), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n695), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n651), .B(new_n793), .C1(new_n1114), .C2(new_n693), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n904), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n1092), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n838), .A2(G330), .A3(new_n423), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n921), .A2(new_n1120), .A3(new_n634), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n667), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1110), .A2(new_n982), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n710), .B1(new_n318), .B2(new_n798), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n757), .A2(new_n292), .B1(new_n758), .B2(new_n540), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1066), .B(new_n1127), .C1(G283), .C2(new_n774), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n257), .B1(new_n765), .B2(G87), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n753), .A2(G116), .B1(KEYINPUT120), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(KEYINPUT120), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(new_n743), .B2(G294), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n813), .A2(new_n1128), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n740), .A2(new_n202), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n765), .A2(new_n1028), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G125), .B2(new_n743), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n257), .B1(new_n762), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G137), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n757), .A2(new_n1140), .B1(new_n758), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(G159), .C2(new_n816), .ZN(new_n1143));
  INV_X1    g0943(.A(G132), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1137), .B(new_n1143), .C1(new_n1144), .C2(new_n752), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1133), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1126), .B1(new_n1146), .B2(new_n723), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1090), .B2(new_n797), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1124), .A2(new_n1125), .A3(new_n1148), .ZN(G378));
  OAI211_X1 g0949(.A(G330), .B(new_n886), .C1(new_n899), .C2(KEYINPUT40), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1090), .A2(new_n914), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n283), .A2(new_n849), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n290), .A2(new_n284), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1153), .B1(new_n290), .B2(new_n284), .ZN(new_n1156));
  XOR2_X1   g0956(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1157));
  OR3_X1    g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AND4_X1   g0961(.A1(new_n1152), .A2(new_n912), .A3(new_n910), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n894), .A2(new_n898), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n911), .B1(new_n1163), .B2(new_n907), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1161), .B1(new_n1164), .B2(new_n1152), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1151), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1160), .B1(new_n913), .B2(new_n919), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n1152), .A3(new_n1161), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1150), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1121), .B1(new_n1110), .B2(new_n1122), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1172), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n666), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n710), .B1(G50), .B2(new_n798), .ZN(new_n1176));
  INV_X1    g0976(.A(G125), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n762), .A2(new_n1177), .B1(new_n758), .B2(new_n1140), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n764), .A2(new_n1141), .B1(new_n757), .B2(new_n1144), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G150), .C2(new_n816), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1138), .B2(new_n752), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1182));
  XNOR2_X1  g0982(.A(new_n1181), .B(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n741), .A2(G159), .ZN(new_n1184));
  AOI211_X1 g0984(.A(G33), .B(G41), .C1(new_n743), .C2(G124), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n741), .A2(new_n754), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n762), .A2(new_n571), .B1(new_n757), .B2(new_n540), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n247), .B1(new_n764), .B2(new_n260), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1188), .A2(new_n1189), .A3(new_n727), .A4(new_n1002), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n743), .A2(G283), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n753), .A2(G107), .B1(new_n1029), .B2(new_n777), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1187), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT58), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1183), .A2(new_n1186), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(G41), .B1(new_n727), .B2(G33), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1195), .B1(new_n1194), .B2(new_n1193), .C1(G50), .C2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1176), .B1(new_n1197), .B2(new_n723), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(new_n1160), .B2(new_n797), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT122), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1170), .B2(new_n983), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1175), .A2(new_n1201), .ZN(G375));
  AND2_X1   g1002(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n921), .A2(new_n1120), .A3(new_n634), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n959), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(new_n1122), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n904), .A2(new_n718), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n710), .B1(G68), .B2(new_n798), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n753), .A2(G137), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n762), .A2(new_n1144), .B1(new_n757), .B2(new_n1141), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(G150), .B2(new_n777), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n335), .B1(G50), .B2(new_n816), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1187), .A2(new_n1210), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n743), .A2(G128), .B1(G159), .B2(new_n765), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT123), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n348), .B1(new_n757), .B2(new_n571), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n764), .A2(new_n540), .B1(new_n762), .B2(new_n443), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1217), .B(new_n1218), .C1(G107), .C2(new_n777), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n753), .A2(G283), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n743), .A2(G303), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1029), .A2(new_n816), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1214), .A2(new_n1216), .B1(new_n1000), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1209), .B1(new_n1224), .B2(new_n723), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1119), .A2(new_n983), .B1(new_n1208), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1207), .A2(new_n1226), .ZN(G381));
  NOR2_X1   g1027(.A1(G375), .A2(G378), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n984), .A2(new_n1078), .A3(new_n1012), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(G393), .A2(G396), .A3(G384), .A4(G381), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(G407));
  INV_X1    g1031(.A(new_n1228), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G407), .B(G213), .C1(G343), .C2(new_n1232), .ZN(G409));
  NAND3_X1  g1033(.A1(new_n1175), .A2(G378), .A3(new_n1201), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1124), .A2(new_n1125), .A3(new_n1148), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1170), .A2(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT124), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1166), .A2(new_n1169), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n982), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1170), .A2(new_n1171), .A3(new_n1206), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1199), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1234), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n642), .A2(G213), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1122), .A2(new_n666), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1205), .A2(KEYINPUT60), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1119), .A2(new_n1121), .A3(KEYINPUT60), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1226), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n822), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1248), .A2(new_n822), .A3(new_n1249), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1243), .A2(new_n1244), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT125), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1244), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1234), .B2(new_n1242), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT125), .A3(new_n1253), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT62), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1261));
  OR3_X1    g1061(.A1(new_n1248), .A2(new_n822), .A3(new_n1249), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(G2897), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1262), .A2(new_n1250), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1262), .B2(new_n1250), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1254), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT126), .B1(new_n1260), .B2(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n785), .B1(new_n1016), .B2(new_n1045), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1078), .B1(new_n984), .B2(new_n1012), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1229), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G387), .A2(G390), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1273), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n984), .A2(new_n1078), .A3(new_n1012), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT62), .ZN(new_n1281));
  AND4_X1   g1081(.A1(KEYINPUT125), .A2(new_n1243), .A3(new_n1244), .A4(new_n1253), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT125), .B1(new_n1258), .B2(new_n1253), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT61), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G2897), .B(new_n1257), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1262), .A2(new_n1250), .A3(new_n1263), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1286), .B1(new_n1289), .B2(new_n1258), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1281), .B1(new_n1258), .B2(new_n1253), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1284), .A2(new_n1285), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1270), .A2(new_n1280), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1256), .A2(new_n1295), .A3(new_n1259), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1253), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1275), .A2(new_n1279), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1267), .A4(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1299), .ZN(G405));
  AOI21_X1  g1100(.A(new_n1235), .B1(new_n1175), .B2(new_n1201), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1232), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1280), .B(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1253), .A2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1304), .B(new_n1306), .ZN(G402));
endmodule


