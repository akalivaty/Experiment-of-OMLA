//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n644, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1255, new_n1256,
    new_n1257;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  AND2_X1   g018(.A1(G2072), .A2(G2078), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g044(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n463), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n463), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n480));
  OAI221_X1 g055(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n463), .B1(new_n484), .B2(new_n485), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n483), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n463), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n484), .B2(new_n485), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n463), .A2(G114), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n488), .B2(G126), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT69), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT69), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT6), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n517), .A2(new_n525), .A3(G62), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n508), .A2(new_n509), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n519), .B1(new_n528), .B2(new_n530), .ZN(G166));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT69), .A2(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n534), .B1(new_n540), .B2(new_n511), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n510), .A2(KEYINPUT71), .A3(new_n512), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(G543), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n532), .B(new_n533), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT7), .Z(new_n547));
  AOI21_X1  g122(.A(new_n522), .B1(new_n510), .B2(new_n512), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(G89), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n551), .B1(new_n513), .B2(new_n534), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n552), .A2(G51), .A3(new_n542), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n532), .B1(new_n553), .B2(new_n533), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n550), .A2(new_n554), .ZN(G168));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n522), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(new_n530), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT73), .Z(new_n560));
  INV_X1    g135(.A(G90), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n513), .A2(new_n517), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n543), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n564), .A2(G52), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(G171));
  NAND3_X1  g141(.A1(new_n552), .A2(G43), .A3(new_n542), .ZN(new_n567));
  NAND2_X1  g142(.A1(G68), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G56), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n522), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n548), .A2(G81), .B1(new_n570), .B2(new_n530), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  NAND4_X1  g153(.A1(new_n541), .A2(G53), .A3(G543), .A4(new_n542), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n552), .A2(new_n581), .A3(G53), .A4(new_n542), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n522), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  INV_X1    g162(.A(G91), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n562), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n583), .A2(new_n590), .ZN(G299));
  INV_X1    g166(.A(G171), .ZN(G301));
  INV_X1    g167(.A(G168), .ZN(G286));
  NAND2_X1  g168(.A1(new_n528), .A2(new_n530), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n518), .B2(new_n514), .ZN(G303));
  INV_X1    g170(.A(G49), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n543), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT74), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n552), .A2(new_n598), .A3(G49), .A4(new_n542), .ZN(new_n599));
  INV_X1    g174(.A(G74), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n537), .B1(new_n522), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n548), .B2(G87), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(G288));
  INV_X1    g178(.A(G73), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT75), .B1(new_n604), .B2(new_n551), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n606), .A2(G73), .A3(G543), .ZN(new_n607));
  INV_X1    g182(.A(G61), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n605), .B(new_n607), .C1(new_n522), .C2(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(G48), .A2(G543), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n609), .A2(new_n530), .B1(new_n513), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n513), .A2(G86), .A3(new_n517), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(G305));
  AOI22_X1  g188(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(new_n529), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n548), .A2(G85), .ZN(new_n616));
  INV_X1    g191(.A(G47), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n543), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n619));
  AND2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(G290));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  INV_X1    g198(.A(G92), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n562), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n548), .A2(KEYINPUT10), .A3(G92), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G66), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G66), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n517), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G79), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n551), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n625), .A2(new_n626), .B1(G651), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n564), .A2(G54), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G171), .B2(new_n636), .ZN(G284));
  OAI21_X1  g213(.A(new_n637), .B1(G171), .B2(new_n636), .ZN(G321));
  NAND2_X1  g214(.A1(G299), .A2(new_n636), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G168), .B2(new_n636), .ZN(G297));
  XNOR2_X1  g216(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g217(.A(new_n635), .ZN(new_n643));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(G860), .ZN(G148));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G868), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n494), .A2(new_n474), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n488), .A2(G123), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT79), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n486), .A2(G135), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n463), .A2(G111), .ZN(new_n657));
  OAI21_X1  g232(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(G2096), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(G2096), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n660), .A3(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT82), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2427), .B(G2430), .Z(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1341), .B(G1348), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2443), .B(G2446), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2451), .B(G2454), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(G14), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G401));
  XOR2_X1   g257(.A(G2084), .B(G2090), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT84), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(KEYINPUT17), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  AOI21_X1  g263(.A(KEYINPUT18), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2100), .ZN(new_n690));
  NOR2_X1   g265(.A1(G2072), .A2(G2078), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n444), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n686), .B2(KEYINPUT18), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G2096), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1961), .B(G1966), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT19), .ZN(new_n699));
  XOR2_X1   g274(.A(G1956), .B(G2474), .Z(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n697), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(KEYINPUT87), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(new_n700), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n705), .A2(new_n699), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n704), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g286(.A(G1991), .B(G1996), .Z(new_n712));
  OR3_X1    g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n710), .B2(new_n711), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1981), .B(G1986), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n716), .A3(new_n714), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(G229));
  NAND2_X1  g294(.A1(new_n573), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G16), .B2(G19), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT93), .B(G1341), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(G162), .A2(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G29), .B2(G35), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT29), .B(G2090), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(G160), .A2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G34), .Z(new_n733));
  OAI21_X1  g308(.A(new_n731), .B1(G29), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n730), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n724), .A2(new_n725), .A3(new_n729), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G33), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  OR3_X1    g315(.A1(new_n740), .A2(KEYINPUT95), .A3(new_n463), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT95), .B1(new_n740), .B2(new_n463), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT25), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G139), .B2(new_n486), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(G29), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT96), .B(G2072), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT30), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n753));
  OR2_X1    g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n752), .A2(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n659), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n735), .B2(new_n734), .ZN(new_n759));
  NOR2_X1   g334(.A1(G27), .A2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G164), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2078), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n750), .A2(new_n759), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n757), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n486), .A2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n488), .A2(G128), .ZN(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n766), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(G2067), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n738), .A2(new_n764), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G16), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n780), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n780), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n757), .A2(G32), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G105), .B2(new_n474), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n486), .A2(G141), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n488), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT98), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n785), .B1(new_n795), .B2(new_n757), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT27), .B(G1996), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n780), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n643), .B2(new_n780), .ZN(new_n800));
  INV_X1    g375(.A(G1348), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n779), .A2(new_n784), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n780), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT23), .ZN(new_n805));
  INV_X1    g380(.A(G299), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n780), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT99), .B(G1956), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n780), .A2(G21), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G168), .B2(new_n780), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(G1966), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(G1966), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n803), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n780), .A2(G23), .ZN(new_n817));
  AND3_X1   g392(.A1(new_n597), .A2(new_n599), .A3(new_n602), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n780), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT91), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n819), .B(new_n820), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n780), .A2(G6), .ZN(new_n827));
  INV_X1    g402(.A(G305), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n780), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT32), .B(G1981), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT90), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n829), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(G166), .A2(G16), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G16), .B2(G22), .ZN(new_n834));
  INV_X1    g409(.A(G1971), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n823), .A2(new_n826), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n486), .A2(G131), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n488), .A2(G119), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n463), .A2(G107), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  MUX2_X1   g422(.A(G25), .B(new_n847), .S(G29), .Z(new_n848));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G1991), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(G290), .B(KEYINPUT88), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n851), .A2(new_n780), .ZN(new_n852));
  NOR2_X1   g427(.A1(G16), .A2(G24), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT89), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT89), .ZN(new_n855));
  INV_X1    g430(.A(new_n853), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n855), .B(new_n856), .C1(new_n851), .C2(new_n780), .ZN(new_n857));
  INV_X1    g432(.A(G1986), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n854), .B2(new_n857), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n842), .B(new_n850), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT92), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n840), .B2(new_n841), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n823), .A2(new_n826), .A3(new_n839), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(KEYINPUT92), .A3(KEYINPUT34), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT36), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n850), .B1(new_n865), .B2(KEYINPUT34), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n854), .A2(new_n857), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G1986), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(new_n859), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT36), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n864), .A2(new_n866), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n816), .B1(new_n868), .B2(new_n875), .ZN(G311));
  AND3_X1   g451(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n872), .B2(new_n874), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n815), .B1(new_n877), .B2(new_n878), .ZN(G150));
  NAND2_X1  g454(.A1(new_n643), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g456(.A1(G80), .A2(G543), .ZN(new_n882));
  INV_X1    g457(.A(G67), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n522), .B2(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n548), .A2(G93), .B1(new_n884), .B2(new_n530), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n541), .A2(G55), .A3(G543), .A4(new_n542), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n572), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n567), .A2(new_n571), .A3(new_n886), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n881), .B(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(KEYINPUT39), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(KEYINPUT39), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(G860), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(G860), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT37), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n895), .A2(new_n897), .ZN(G145));
  XNOR2_X1  g473(.A(G160), .B(new_n490), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n659), .Z(new_n900));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n495), .A2(G2105), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n470), .B2(new_n471), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n904), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n496), .ZN(new_n905));
  OAI211_X1 g480(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n502), .A2(new_n503), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n902), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n501), .A2(new_n505), .A3(KEYINPUT100), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n775), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n774), .A3(new_n773), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n901), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n914), .A3(new_n901), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n794), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n795), .B1(new_n919), .B2(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n747), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n912), .A2(new_n914), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT102), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n912), .A2(new_n914), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n793), .ZN(new_n928));
  INV_X1    g503(.A(new_n793), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n746), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n651), .B(new_n847), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n486), .A2(G142), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT103), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n488), .A2(G130), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n463), .A2(G118), .ZN(new_n936));
  OAI21_X1  g511(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n932), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT104), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n922), .A2(new_n931), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n922), .B2(new_n931), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n900), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n922), .A2(new_n931), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n939), .ZN(new_n946));
  INV_X1    g521(.A(new_n900), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT105), .B(G37), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n944), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g526(.A1(G290), .A2(new_n828), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  NOR2_X1   g528(.A1(G303), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(G166), .A2(KEYINPUT107), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G288), .ZN(new_n957));
  OAI211_X1 g532(.A(G305), .B(new_n615), .C1(new_n620), .C2(new_n621), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n818), .B1(new_n954), .B2(new_n955), .ZN(new_n959));
  AND4_X1   g534(.A1(new_n952), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n952), .A2(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT42), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  NAND2_X1  g539(.A1(G299), .A2(new_n635), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n583), .A2(new_n633), .A3(new_n590), .A4(new_n634), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(KEYINPUT41), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT41), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n965), .B2(new_n966), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n969), .A3(new_n966), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n973), .B2(new_n964), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n646), .B(new_n891), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n967), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(new_n975), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n963), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n963), .A2(new_n978), .ZN(new_n980));
  OAI21_X1  g555(.A(G868), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n887), .A2(new_n636), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(G295));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n982), .ZN(G331));
  INV_X1    g559(.A(new_n962), .ZN(new_n985));
  NAND2_X1  g560(.A1(G168), .A2(new_n890), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n888), .B(new_n889), .C1(new_n550), .C2(new_n554), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(G301), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(G171), .A3(new_n987), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n972), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n964), .B1(new_n992), .B2(new_n970), .ZN(new_n993));
  INV_X1    g568(.A(new_n968), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n967), .B1(new_n989), .B2(new_n990), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  INV_X1    g573(.A(G37), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n991), .A2(new_n977), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n962), .B(new_n1000), .C1(new_n974), .C2(new_n991), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n993), .A2(new_n994), .ZN(new_n1004));
  INV_X1    g579(.A(new_n991), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n996), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G37), .B1(new_n1006), .B2(new_n962), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n998), .A4(new_n997), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n991), .B1(new_n971), .B2(new_n972), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n985), .B1(new_n1012), .B2(new_n996), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(new_n949), .A3(new_n1001), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1011), .B1(new_n1014), .B2(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n998), .B1(new_n1007), .B2(new_n997), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(G397));
  INV_X1    g596(.A(KEYINPUT125), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n1023));
  OAI211_X1 g598(.A(G303), .B(G8), .C1(new_n1023), .C2(KEYINPUT55), .ZN(new_n1024));
  XOR2_X1   g599(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(G166), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G125), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1029), .B1(new_n493), .B2(new_n464), .ZN(new_n1030));
  INV_X1    g605(.A(new_n468), .ZN(new_n1031));
  OAI21_X1  g606(.A(G2105), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(G40), .A3(new_n472), .A4(new_n475), .ZN(new_n1033));
  INV_X1    g608(.A(G1384), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n905), .B2(new_n908), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(G1384), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n909), .A2(new_n910), .A3(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1037), .A2(KEYINPUT111), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT111), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1040), .A2(new_n1041), .A3(G1971), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1033), .B1(new_n1035), .B2(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n1034), .C1(new_n905), .C2(new_n908), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G2090), .ZN(new_n1047));
  OAI211_X1 g622(.A(G8), .B(new_n1028), .C1(new_n1042), .C2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n597), .A2(G1976), .A3(new_n599), .A4(new_n602), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(new_n1026), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(KEYINPUT52), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G40), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n469), .A2(new_n476), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1384), .B1(new_n501), .B2(new_n505), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n513), .A2(new_n610), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n605), .A2(new_n607), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n608), .B1(new_n515), .B2(new_n516), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n530), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n612), .A2(new_n1064), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n611), .A2(KEYINPUT114), .A3(new_n1068), .A4(new_n612), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G305), .A2(G1981), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1063), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1071), .A2(new_n1072), .B1(G1981), .B2(G305), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT49), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(G288), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1077), .A2(new_n1079), .B1(new_n1052), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1048), .A2(new_n1058), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT111), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n909), .A2(new_n910), .A3(new_n1038), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1060), .B1(new_n1061), .B2(KEYINPUT45), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1037), .A2(new_n1039), .A3(KEYINPUT111), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n835), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1061), .A2(new_n1090), .A3(new_n1044), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1045), .A2(KEYINPUT116), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1043), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1089), .B1(G2090), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1028), .B1(new_n1094), .B2(G8), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1022), .B1(new_n1083), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1056), .B1(new_n1055), .B2(KEYINPUT52), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT113), .B(new_n1053), .C1(new_n1049), .C2(new_n1051), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1052), .A2(new_n1081), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1079), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1051), .B1(new_n1078), .B2(KEYINPUT49), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1093), .A2(G2090), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n1042), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1028), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(KEYINPUT125), .A4(new_n1048), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1096), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1348), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1062), .A2(G2067), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n643), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n1117));
  INV_X1    g692(.A(G1996), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1037), .A2(new_n1039), .A3(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1062), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1122), .B2(new_n573), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n572), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1112), .A2(new_n635), .A3(new_n1115), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n643), .B1(new_n1114), .B2(new_n1111), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1113), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(G299), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n583), .A2(new_n590), .A3(new_n1131), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1131), .B1(new_n583), .B2(new_n590), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1132), .B(new_n589), .C1(new_n580), .C2(new_n582), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1136), .A2(new_n1137), .A3(KEYINPUT120), .ZN(new_n1138));
  INV_X1    g713(.A(G1956), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1093), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1135), .A2(new_n1138), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1141), .A2(new_n1142), .B1(new_n1093), .B2(new_n1139), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1144), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1145), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1129), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1144), .A2(new_n1127), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1150), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1046), .A2(new_n783), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1038), .B1(new_n905), .B2(new_n908), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1159), .B(new_n1060), .C1(new_n1061), .C2(KEYINPUT45), .ZN(new_n1160));
  OAI21_X1  g735(.A(KEYINPUT124), .B1(new_n1160), .B2(G2078), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1037), .A2(new_n1162), .A3(new_n762), .A4(new_n1159), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(KEYINPUT53), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(G2078), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1158), .B(new_n1164), .C1(new_n1165), .C2(KEYINPUT53), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1157), .B1(new_n1167), .B2(G301), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1036), .B1(new_n911), .B2(G1384), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n762), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1169), .A2(new_n1039), .A3(new_n1170), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1158), .B(new_n1171), .C1(new_n1165), .C2(KEYINPUT53), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(G171), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1153), .A2(new_n1156), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1060), .B1(new_n1061), .B2(new_n1044), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1045), .A2(new_n735), .ZN(new_n1177));
  OAI21_X1  g752(.A(KEYINPUT117), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(G1966), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1160), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT117), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1043), .A2(new_n1181), .A3(new_n735), .A4(new_n1045), .ZN(new_n1182));
  NAND4_X1  g757(.A1(G168), .A2(new_n1178), .A3(new_n1180), .A4(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT51), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1026), .B1(KEYINPUT121), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(KEYINPUT121), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1183), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1178), .A2(new_n1182), .A3(new_n1180), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1189), .A2(G286), .A3(G8), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1187), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1175), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1192), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(KEYINPUT122), .A3(new_n1190), .A4(new_n1188), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1197));
  NOR2_X1   g772(.A1(new_n1167), .A2(G301), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1172), .A2(G171), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1110), .A2(new_n1174), .A3(new_n1196), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1196), .A2(KEYINPUT62), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1193), .A2(new_n1195), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1110), .A2(new_n1202), .A3(new_n1204), .A4(new_n1198), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT118), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1189), .A2(G8), .A3(G168), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1048), .A2(new_n1058), .A3(new_n1082), .A4(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1208), .B2(new_n1095), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1208), .A2(new_n1206), .A3(new_n1095), .ZN(new_n1212));
  OAI21_X1  g787(.A(G8), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n1107), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1214), .A2(KEYINPUT63), .ZN(new_n1215));
  OAI22_X1  g790(.A1(new_n1211), .A2(new_n1212), .B1(new_n1208), .B2(new_n1215), .ZN(new_n1216));
  NOR3_X1   g791(.A1(new_n1048), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1217));
  OAI211_X1 g792(.A(new_n1080), .B(new_n818), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1073), .ZN(new_n1219));
  XNOR2_X1  g794(.A(new_n1051), .B(KEYINPUT115), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1217), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1201), .A2(new_n1205), .A3(new_n1216), .A4(new_n1221), .ZN(new_n1222));
  INV_X1    g797(.A(G290), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1169), .A2(new_n1033), .ZN(new_n1224));
  NAND3_X1  g799(.A1(new_n1223), .A2(new_n858), .A3(new_n1224), .ZN(new_n1225));
  NAND3_X1  g800(.A1(G290), .A2(G1986), .A3(new_n1224), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g802(.A(new_n1227), .B(KEYINPUT110), .Z(new_n1228));
  XNOR2_X1  g803(.A(new_n775), .B(new_n777), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n793), .A2(G1996), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1229), .B(new_n1230), .C1(G1996), .C2(new_n794), .ZN(new_n1231));
  INV_X1    g806(.A(new_n849), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n847), .B(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1224), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  AND2_X1   g809(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1222), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1229), .A2(new_n929), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT46), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1224), .A2(new_n1118), .ZN(new_n1239));
  AOI22_X1  g814(.A1(new_n1237), .A2(new_n1224), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g815(.A1(new_n1239), .A2(new_n1238), .ZN(new_n1241));
  AND2_X1   g816(.A1(new_n1241), .A2(KEYINPUT126), .ZN(new_n1242));
  NOR2_X1   g817(.A1(new_n1241), .A2(KEYINPUT126), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1240), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g819(.A(new_n1244), .B(KEYINPUT47), .Z(new_n1245));
  OR2_X1    g820(.A1(new_n847), .A2(new_n1232), .ZN(new_n1246));
  OAI22_X1  g821(.A1(new_n1231), .A2(new_n1246), .B1(G2067), .B2(new_n775), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1247), .A2(new_n1224), .ZN(new_n1248));
  XNOR2_X1  g823(.A(new_n1234), .B(KEYINPUT127), .ZN(new_n1249));
  XOR2_X1   g824(.A(new_n1225), .B(KEYINPUT48), .Z(new_n1250));
  OAI21_X1  g825(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NOR2_X1   g826(.A1(new_n1245), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1236), .A2(new_n1252), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g828(.A1(G227), .A2(new_n461), .ZN(new_n1255));
  NAND2_X1  g829(.A1(new_n681), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g830(.A(new_n1256), .B1(new_n717), .B2(new_n718), .ZN(new_n1257));
  OAI211_X1 g831(.A(new_n950), .B(new_n1257), .C1(new_n1018), .C2(new_n1019), .ZN(G225));
  INV_X1    g832(.A(G225), .ZN(G308));
endmodule


