//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G113), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n196), .ZN(new_n198));
  XNOR2_X1  g012(.A(G116), .B(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n200), .A3(KEYINPUT67), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT67), .B1(new_n197), .B2(new_n200), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT30), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(new_n207), .B2(G143), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n205), .A3(G146), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n207), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n205), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G134), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(G134), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n222), .B1(new_n220), .B2(new_n221), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT11), .A2(G134), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G137), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n222), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n219), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n225), .A2(new_n224), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT65), .A2(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT65), .A2(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(G137), .A3(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n233), .A2(new_n219), .A3(new_n231), .A4(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n218), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G143), .B(G146), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G128), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n214), .B2(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n211), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(G137), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n222), .A2(G134), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n237), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n204), .B1(new_n239), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n231), .B(new_n236), .C1(new_n246), .C2(KEYINPUT11), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n217), .B1(new_n252), .B2(new_n237), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n237), .A2(new_n245), .A3(new_n248), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT30), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n203), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n203), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n239), .A2(new_n257), .A3(new_n249), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G101), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n253), .A2(new_n254), .A3(new_n203), .ZN(new_n267));
  INV_X1    g081(.A(new_n264), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n256), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n256), .A2(new_n269), .A3(KEYINPUT31), .A4(new_n265), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n203), .B1(new_n253), .B2(new_n254), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n258), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n267), .A2(KEYINPUT28), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(KEYINPUT70), .B(new_n268), .C1(new_n277), .C2(new_n278), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n187), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT32), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n267), .A2(new_n266), .A3(new_n268), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n258), .B2(new_n264), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT31), .B1(new_n288), .B2(new_n256), .ZN(new_n289));
  INV_X1    g103(.A(new_n273), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n281), .B(new_n282), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n292), .A3(new_n187), .ZN(new_n293));
  INV_X1    g107(.A(new_n256), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n268), .B1(new_n294), .B2(new_n267), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n257), .B1(new_n239), .B2(new_n249), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT28), .B1(new_n297), .B2(new_n267), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n258), .A2(new_n275), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n264), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n301), .B(new_n302), .C1(new_n296), .C2(new_n300), .ZN(new_n303));
  AOI22_X1  g117(.A1(new_n285), .A2(new_n293), .B1(G472), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G217), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(G234), .B2(new_n302), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT22), .B(G137), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n308), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n188), .A2(G128), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n188), .A2(G128), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G110), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT24), .B(G110), .Z(new_n317));
  XNOR2_X1  g131(.A(G119), .B(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G125), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT71), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n324), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G125), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT71), .B(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n207), .B(new_n329), .C1(new_n333), .C2(KEYINPUT16), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT16), .B1(new_n335), .B2(new_n330), .ZN(new_n336));
  INV_X1    g150(.A(new_n329), .ZN(new_n337));
  AOI21_X1  g151(.A(G146), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n321), .B1(new_n334), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT72), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n341), .B(new_n321), .C1(new_n334), .C2(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(G146), .A3(new_n337), .ZN(new_n344));
  XNOR2_X1  g158(.A(G125), .B(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n207), .ZN(new_n346));
  OAI22_X1  g160(.A1(new_n315), .A2(G110), .B1(new_n317), .B2(new_n318), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n311), .B1(new_n343), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  INV_X1    g164(.A(new_n311), .ZN(new_n351));
  AOI211_X1 g165(.A(new_n350), .B(new_n351), .C1(new_n340), .C2(new_n342), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n307), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT25), .B1(new_n353), .B2(new_n302), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n327), .A2(G125), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n325), .A2(KEYINPUT71), .ZN(new_n359));
  OAI21_X1  g173(.A(G140), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n322), .B1(new_n360), .B2(new_n331), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n207), .B1(new_n361), .B2(new_n329), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n344), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n341), .B1(new_n363), .B2(new_n321), .ZN(new_n364));
  AOI211_X1 g178(.A(KEYINPUT72), .B(new_n320), .C1(new_n362), .C2(new_n344), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n348), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n351), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n343), .A2(new_n348), .A3(new_n311), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(KEYINPUT25), .A3(new_n302), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n306), .B1(new_n357), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n356), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT74), .B1(new_n304), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n303), .A2(G472), .ZN(new_n374));
  INV_X1    g188(.A(new_n187), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n298), .A2(new_n299), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT70), .B1(new_n376), .B2(new_n268), .ZN(new_n377));
  INV_X1    g191(.A(new_n282), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n272), .A2(new_n273), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT32), .B(new_n375), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n292), .B1(new_n291), .B2(new_n187), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n374), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT74), .ZN(new_n384));
  INV_X1    g198(.A(new_n372), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G221), .B1(new_n390), .B2(G902), .ZN(new_n391));
  OAI21_X1  g205(.A(G214), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  AOI22_X1  g209(.A1(KEYINPUT76), .A2(new_n394), .B1(new_n395), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  AND4_X1   g212(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT3), .A4(G104), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n397), .A2(KEYINPUT3), .B1(new_n398), .B2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G101), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(G101), .ZN(new_n404));
  INV_X1    g218(.A(G101), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n396), .C1(new_n399), .C2(new_n400), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(KEYINPUT4), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n203), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n193), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n199), .A2(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n412), .A2(new_n200), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n398), .A2(G104), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n395), .A2(G107), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n405), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI22_X1  g230(.A1(new_n397), .A2(KEYINPUT3), .B1(new_n398), .B2(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n414), .B1(KEYINPUT76), .B2(new_n394), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT3), .A4(G104), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n416), .B1(new_n420), .B2(new_n405), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n408), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n408), .A2(new_n424), .A3(new_n422), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n245), .A2(new_n332), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n332), .B2(new_n217), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n309), .A2(G224), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n428), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(KEYINPUT7), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n436), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n431), .B(new_n438), .C1(new_n332), .C2(new_n217), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(new_n427), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n424), .B(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT80), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n411), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n410), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n411), .A2(new_n444), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n421), .B(new_n200), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  OAI22_X1  g262(.A1(new_n448), .A2(KEYINPUT81), .B1(new_n421), .B2(new_n413), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n443), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(G902), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n435), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT82), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n435), .A2(new_n452), .A3(new_n454), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n393), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT78), .ZN(new_n459));
  OAI21_X1  g273(.A(G128), .B1(new_n206), .B2(new_n241), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(new_n216), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT77), .B1(new_n244), .B2(new_n240), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n463), .A3(new_n242), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n421), .ZN(new_n465));
  INV_X1    g279(.A(new_n416), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n406), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n211), .A2(new_n244), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n242), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n252), .A2(new_n237), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n470), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT12), .B1(new_n470), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n471), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(KEYINPUT12), .A3(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT10), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n465), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n407), .A2(new_n218), .A3(new_n403), .ZN(new_n482));
  INV_X1    g296(.A(new_n471), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n245), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G140), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n309), .A2(G227), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n486), .B(new_n487), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n474), .A2(new_n479), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n471), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n485), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n302), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n302), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n477), .A2(new_n478), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n485), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n488), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(new_n485), .A3(new_n489), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(G469), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT85), .ZN(new_n509));
  XNOR2_X1  g323(.A(G128), .B(G143), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT13), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n243), .A2(KEYINPUT13), .A3(G143), .ZN(new_n512));
  INV_X1    g326(.A(G134), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n220), .A2(new_n221), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n510), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n190), .B2(G122), .ZN(new_n519));
  INV_X1    g333(.A(G122), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT84), .A3(G116), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n190), .A2(G122), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n398), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n398), .B1(new_n522), .B2(new_n523), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n515), .B(new_n517), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n516), .B(new_n510), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(KEYINPUT14), .ZN(new_n529));
  OR3_X1    g343(.A1(new_n520), .A2(KEYINPUT14), .A3(G116), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G107), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n532), .A3(new_n524), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n309), .A2(G217), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n390), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n527), .B2(new_n533), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n302), .B(new_n509), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n527), .A2(new_n533), .ZN(new_n540));
  INV_X1    g354(.A(new_n535), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n538), .B(new_n539), .C1(new_n544), .C2(new_n508), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(KEYINPUT86), .A3(new_n509), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  INV_X1    g362(.A(G237), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n309), .A3(G214), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n205), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(KEYINPUT17), .A3(G131), .ZN(new_n554));
  INV_X1    g368(.A(new_n552), .ZN(new_n555));
  AOI21_X1  g369(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n551), .A2(new_n219), .A3(new_n552), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n362), .A2(new_n344), .A3(new_n554), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G113), .B(G122), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(new_n395), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n346), .B1(new_n333), .B2(new_n207), .ZN(new_n564));
  NAND2_X1  g378(.A1(KEYINPUT18), .A2(G131), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n552), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n553), .A2(KEYINPUT18), .A3(G131), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n557), .A2(new_n559), .ZN(new_n570));
  OAI211_X1 g384(.A(KEYINPUT19), .B(new_n331), .C1(new_n332), .C2(new_n323), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n345), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n571), .A2(new_n207), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n344), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n568), .ZN(new_n576));
  INV_X1    g390(.A(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(G475), .A2(G902), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n580), .B(KEYINPUT83), .Z(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n548), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  AOI211_X1 g397(.A(KEYINPUT20), .B(new_n581), .C1(new_n569), .C2(new_n578), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n568), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n586), .B2(new_n569), .ZN(new_n587));
  INV_X1    g401(.A(G475), .ZN(new_n588));
  OAI22_X1  g402(.A1(new_n583), .A2(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n309), .A2(G952), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(G234), .B2(G237), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n302), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT21), .B(G898), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n547), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n391), .A2(new_n458), .A3(new_n506), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n387), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n291), .A2(new_n302), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(G472), .B1(new_n187), .B2(new_n291), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n506), .A2(new_n391), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n385), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(KEYINPUT87), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(KEYINPUT87), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n435), .A2(new_n452), .A3(new_n454), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n454), .B1(new_n435), .B2(new_n452), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n392), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n603), .A2(new_n604), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n544), .A2(new_n507), .ZN(new_n609));
  NAND2_X1  g423(.A1(G478), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n542), .B2(KEYINPUT88), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n542), .A2(new_n543), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n609), .B(new_n610), .C1(new_n614), .C2(new_n507), .ZN(new_n615));
  INV_X1    g429(.A(new_n589), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n594), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(KEYINPUT89), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n583), .B2(new_n584), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n563), .B1(new_n575), .B2(new_n568), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n334), .A2(new_n338), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n560), .A2(new_n554), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n625), .B1(new_n629), .B2(new_n563), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT20), .B1(new_n630), .B2(new_n581), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n579), .A2(new_n548), .A3(new_n582), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(KEYINPUT89), .A3(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n545), .B(new_n546), .C1(new_n588), .C2(new_n587), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n594), .B(KEYINPUT90), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n608), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G107), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  AOI21_X1  g455(.A(new_n350), .B1(new_n340), .B2(new_n342), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n642), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n307), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT91), .B1(new_n371), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n306), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n367), .A2(new_n302), .A3(new_n368), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT25), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n648), .B1(new_n651), .B2(new_n369), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT91), .ZN(new_n653));
  INV_X1    g467(.A(new_n646), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n596), .A2(new_n656), .A3(new_n600), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT92), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT37), .B(G110), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND3_X1  g474(.A1(new_n371), .A2(KEYINPUT91), .A3(new_n646), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n285), .A2(new_n293), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n374), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT94), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT93), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n591), .B1(new_n592), .B2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n634), .A2(new_n667), .A3(new_n636), .A4(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n624), .A2(new_n633), .A3(new_n670), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT93), .B1(new_n672), .B2(new_n635), .ZN(new_n673));
  INV_X1    g487(.A(new_n454), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n453), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n393), .B1(new_n675), .B2(new_n457), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n671), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n665), .A2(new_n666), .A3(new_n601), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n383), .A2(new_n656), .A3(new_n677), .A4(new_n601), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT94), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XOR2_X1   g496(.A(new_n669), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n601), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n652), .A2(new_n654), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n264), .B1(new_n258), .B2(new_n276), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT95), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n270), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n692), .B2(G902), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n664), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n455), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n435), .B2(new_n452), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n605), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT38), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT38), .B1(new_n605), .B2(new_n696), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n545), .A2(new_n546), .A3(new_n392), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n616), .A2(new_n702), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n689), .A2(new_n694), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n687), .A2(new_n688), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT97), .B(G143), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G45));
  AND3_X1   g521(.A1(new_n383), .A2(new_n601), .A3(new_n656), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n615), .A2(new_n616), .A3(new_n669), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n709), .A2(new_n676), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  NAND2_X1  g526(.A1(new_n496), .A2(new_n302), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n391), .A3(new_n498), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n607), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n383), .A2(new_n385), .A3(new_n619), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT98), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n715), .A2(new_n618), .A3(new_n594), .A4(new_n607), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n385), .A4(new_n383), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n383), .A2(new_n385), .A3(new_n638), .A4(new_n716), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n383), .A2(new_n656), .A3(new_n595), .A4(new_n716), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT99), .B(G119), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G21));
  INV_X1    g543(.A(G472), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n730), .B1(new_n291), .B2(new_n302), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n375), .B1(new_n380), .B2(new_n279), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n703), .B(new_n637), .C1(new_n605), .C2(new_n606), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n715), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n735), .A3(new_n385), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT100), .B(G122), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G24));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n599), .A2(G472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n371), .A2(new_n646), .ZN(new_n742));
  INV_X1    g556(.A(new_n732), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n741), .A2(new_n709), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n736), .A2(new_n676), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n740), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n731), .A2(new_n689), .A3(new_n732), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n747), .A2(KEYINPUT101), .A3(new_n709), .A4(new_n716), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  AOI21_X1  g564(.A(new_n489), .B1(new_n501), .B2(new_n485), .ZN(new_n751));
  INV_X1    g565(.A(new_n504), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT102), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT102), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n504), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n498), .A3(new_n500), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n605), .A2(new_n696), .A3(new_n393), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n757), .A2(new_n391), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n383), .A2(new_n385), .A3(new_n759), .A4(new_n709), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT103), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n372), .B1(new_n664), .B2(new_n374), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT42), .A3(new_n709), .A4(new_n759), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n760), .A2(new_n761), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT103), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  INV_X1    g585(.A(KEYINPUT104), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n671), .A2(new_n673), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n765), .A2(new_n772), .A3(new_n773), .A4(new_n759), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n383), .A2(new_n385), .A3(new_n759), .A4(new_n773), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n600), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT107), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n781));
  OR3_X1    g595(.A1(new_n615), .A2(new_n589), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n783));
  OAI22_X1  g597(.A1(new_n615), .A2(new_n589), .B1(new_n783), .B2(new_n781), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n689), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT44), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n503), .A2(new_n504), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n497), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n753), .A2(KEYINPUT45), .A3(new_n755), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n499), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n498), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT105), .B1(new_n795), .B2(KEYINPUT46), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT106), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT105), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT106), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n498), .A4(new_n796), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n795), .A2(KEYINPUT46), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n806), .A2(new_n391), .A3(new_n683), .ZN(new_n807));
  INV_X1    g621(.A(new_n758), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n787), .B2(KEYINPUT44), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n790), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT109), .B(G137), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G39));
  AND3_X1   g626(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n391), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n806), .B2(new_n391), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n372), .A2(new_n709), .A3(new_n758), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n383), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n323), .ZN(G42));
  NAND2_X1  g632(.A1(new_n714), .A2(new_n498), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT110), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT49), .Z(new_n821));
  INV_X1    g635(.A(new_n391), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n615), .A2(new_n822), .A3(new_n393), .A4(new_n589), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n385), .A2(new_n823), .ZN(new_n824));
  OR4_X1    g638(.A1(new_n694), .A2(new_n821), .A3(new_n701), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n587), .A2(new_n588), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n672), .A2(new_n826), .A3(new_n547), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n383), .A2(new_n656), .A3(new_n601), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n757), .A2(new_n391), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n747), .A2(new_n709), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n758), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n777), .A2(KEYINPUT112), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT112), .B1(new_n777), .B2(new_n832), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n387), .A2(new_n596), .B1(new_n718), .B2(new_n721), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n725), .A2(new_n727), .A3(new_n657), .A4(new_n737), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n458), .A2(new_n637), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n616), .A2(new_n547), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n838), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n840), .A2(KEYINPUT111), .B1(new_n841), .B2(new_n617), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT111), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n602), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n764), .A2(new_n836), .A3(new_n846), .A4(new_n769), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n835), .A2(KEYINPUT53), .A3(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n708), .A2(new_n710), .B1(new_n746), .B2(new_n748), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n702), .B(new_n616), .C1(new_n457), .C2(new_n675), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n742), .A2(new_n669), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n694), .A2(new_n850), .A3(new_n829), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n681), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n853), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT113), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n854), .B1(new_n856), .B2(KEYINPUT52), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  AOI211_X1 g672(.A(KEYINPUT113), .B(new_n858), .C1(new_n853), .C2(new_n855), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n848), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n836), .A2(new_n846), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n770), .B(new_n861), .C1(new_n834), .C2(new_n833), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n853), .A2(KEYINPUT52), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n849), .A2(new_n681), .A3(new_n858), .A4(new_n852), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT53), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n860), .A2(KEYINPUT54), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n766), .B2(new_n767), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n836), .A2(new_n846), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n835), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n857), .B2(new_n859), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n868), .B1(new_n862), .B2(new_n865), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n694), .ZN(new_n876));
  INV_X1    g690(.A(new_n591), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n715), .A2(new_n808), .A3(new_n372), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n617), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n590), .B(KEYINPUT118), .Z(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n782), .B2(new_n784), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n733), .A3(new_n385), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n879), .B(new_n880), .C1(new_n745), .C2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n808), .A2(new_n715), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT116), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT116), .B1(new_n881), .B2(new_n884), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n765), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n887), .A2(KEYINPUT48), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT48), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n882), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n758), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n820), .A2(new_n822), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n815), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT50), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n701), .A2(new_n392), .A3(new_n715), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n898), .B2(new_n882), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n892), .A2(KEYINPUT50), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n747), .B1(new_n885), .B2(new_n886), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n876), .A2(new_n878), .A3(new_n616), .A4(new_n615), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT117), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n901), .A2(new_n906), .A3(new_n902), .A4(new_n903), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(KEYINPUT51), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n891), .B1(new_n895), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n806), .A2(new_n391), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT47), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n806), .A2(KEYINPUT47), .A3(new_n391), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n894), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n758), .A3(new_n892), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n902), .A2(new_n903), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n901), .A2(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT51), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n867), .A2(new_n875), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n867), .A2(new_n875), .A3(new_n921), .A4(KEYINPUT119), .ZN(new_n925));
  OR2_X1    g739(.A1(G952), .A2(G953), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n825), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT120), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n930), .B(new_n825), .C1(new_n924), .C2(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G75));
  NOR2_X1   g746(.A1(new_n309), .A2(G952), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n428), .A2(new_n430), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n434), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n302), .B1(new_n872), .B2(new_n874), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(G210), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n455), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n936), .A2(new_n939), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n933), .B(new_n940), .C1(new_n941), .C2(new_n942), .ZN(G51));
  NAND2_X1  g757(.A1(new_n872), .A2(new_n874), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n875), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(new_n499), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n496), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n937), .A2(new_n794), .A3(new_n793), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n933), .B1(new_n950), .B2(new_n951), .ZN(G54));
  INV_X1    g766(.A(new_n933), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n937), .A2(KEYINPUT58), .A3(G475), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n579), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n579), .B2(new_n954), .ZN(G60));
  XOR2_X1   g770(.A(new_n610), .B(KEYINPUT59), .Z(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n867), .B2(new_n875), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n953), .B1(new_n958), .B2(new_n614), .ZN(new_n959));
  INV_X1    g773(.A(new_n614), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT122), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G63));
  NAND2_X1  g779(.A1(G217), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  NAND2_X1  g781(.A1(new_n944), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n354), .A2(new_n355), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n933), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n944), .A2(new_n645), .A3(new_n967), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT61), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT124), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT124), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n970), .A2(new_n975), .A3(KEYINPUT61), .A4(new_n972), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n972), .B(KEYINPUT123), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n978), .B1(new_n979), .B2(new_n971), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n977), .A2(new_n980), .ZN(G66));
  NOR2_X1   g795(.A1(new_n861), .A2(G953), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  INV_X1    g797(.A(G224), .ZN(new_n984));
  OAI21_X1  g798(.A(G953), .B1(new_n593), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n934), .B1(G898), .B2(new_n309), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(G69));
  NAND2_X1  g802(.A1(G900), .A2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n770), .A2(new_n777), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT127), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n810), .A2(new_n817), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n849), .A2(new_n681), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n807), .A2(new_n765), .A3(new_n850), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n991), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n989), .B1(new_n995), .B2(G953), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n250), .A2(new_n255), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n571), .A2(new_n573), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT126), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n705), .A2(new_n993), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT62), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n808), .B1(new_n618), .B2(new_n839), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n387), .A2(new_n601), .A3(new_n683), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1002), .A2(new_n992), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1000), .A2(G953), .ZN(new_n1006));
  AOI22_X1  g820(.A1(new_n996), .A2(new_n1000), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  INV_X1    g825(.A(new_n861), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n294), .A2(new_n267), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1014), .A2(new_n268), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n933), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1011), .B1(new_n995), .B2(new_n1012), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1017), .A2(new_n268), .A3(new_n1014), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n295), .A2(new_n270), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n860), .A2(new_n866), .A3(new_n1011), .A4(new_n1019), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n1016), .A2(new_n1018), .A3(new_n1020), .ZN(G57));
endmodule


