//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND3_X1  g0009(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n209), .B1(new_n210), .B2(new_n212), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G58), .B(G77), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n236), .B(new_n237), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  OAI211_X1 g0046(.A(G1), .B(G13), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G45), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n247), .A2(G274), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n250), .B1(new_n253), .B2(new_n215), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(G33), .B2(G41), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n228), .A2(G1698), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n257), .B(new_n258), .C1(G226), .C2(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n254), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g0062(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n263));
  XNOR2_X1  g0063(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G200), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT72), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n264), .A2(KEYINPUT72), .A3(G200), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n255), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G20), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n273), .A2(new_n202), .B1(new_n274), .B2(G68), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n245), .A2(new_n216), .A3(G20), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT11), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G68), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n282), .B(KEYINPUT12), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n271), .B1(new_n251), .B2(G20), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(G68), .B2(new_n284), .ZN(new_n285));
  AND3_X1   g0085(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n262), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n263), .B2(new_n262), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G190), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n269), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n264), .A2(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT14), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(G179), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT14), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n264), .A2(new_n295), .A3(G169), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n286), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT74), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT3), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(G33), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n245), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(G33), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G223), .B2(G1698), .ZN(new_n309));
  INV_X1    g0109(.A(G87), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n306), .A2(new_n309), .B1(new_n245), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n256), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n250), .B1(new_n253), .B2(new_n228), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G190), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n256), .B2(new_n311), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT8), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G58), .ZN(new_n326));
  INV_X1    g0126(.A(G58), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(KEYINPUT8), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT68), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n281), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n330), .B2(new_n284), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n327), .A2(new_n214), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n272), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n306), .A2(new_n338), .A3(new_n274), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G68), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n338), .B1(new_n306), .B2(new_n274), .ZN(new_n341));
  OAI211_X1 g0141(.A(KEYINPUT16), .B(new_n337), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT7), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n257), .B2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n305), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n345), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n350), .A3(new_n274), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n214), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n343), .B1(new_n352), .B2(new_n336), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n342), .A2(new_n353), .A3(new_n271), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n321), .A2(new_n332), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT17), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(new_n332), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n315), .A2(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n318), .A2(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT18), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(new_n364), .A3(new_n361), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n321), .A2(KEYINPUT17), .A3(new_n332), .A4(new_n354), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n357), .A2(new_n363), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G223), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n347), .A2(new_n305), .A3(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT67), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n257), .A2(KEYINPUT67), .A3(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n257), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G222), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n375), .A2(new_n376), .B1(new_n216), .B2(new_n257), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n256), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n250), .B1(new_n253), .B2(new_n307), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G169), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n245), .A2(G20), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n324), .A2(new_n329), .A3(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n272), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n271), .ZN(new_n388));
  OAI21_X1  g0188(.A(G50), .B1(new_n274), .B2(G1), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n389), .B(KEYINPUT69), .Z(new_n390));
  AND3_X1   g0190(.A1(new_n281), .A2(new_n255), .A3(new_n270), .ZN(new_n391));
  INV_X1    g0191(.A(new_n281), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n390), .A2(new_n391), .B1(new_n202), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n378), .A2(new_n395), .A3(new_n380), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n383), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT67), .B1(new_n257), .B2(G1698), .ZN(new_n399));
  AND4_X1   g0199(.A1(KEYINPUT67), .A2(new_n347), .A3(new_n305), .A4(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(G223), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n348), .A2(G1698), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(G222), .B1(G77), .B2(new_n348), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n247), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G200), .B1(new_n404), .B2(new_n379), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT9), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n388), .B2(new_n393), .ZN(new_n407));
  INV_X1    g0207(.A(new_n271), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n385), .B2(new_n386), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n389), .B(KEYINPUT69), .ZN(new_n410));
  INV_X1    g0210(.A(new_n391), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n410), .A2(new_n411), .B1(G50), .B2(new_n281), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT9), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n405), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT70), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n381), .B2(new_n316), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n414), .A2(KEYINPUT10), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n388), .A2(new_n393), .A3(new_n406), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT9), .B1(new_n409), .B2(new_n412), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n419), .A2(new_n420), .B1(new_n381), .B2(G200), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n404), .A2(new_n379), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT70), .B1(new_n422), .B2(G190), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n418), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n398), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n322), .A2(new_n273), .B1(new_n274), .B2(new_n216), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n426), .B1(new_n384), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(new_n408), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n284), .A2(G77), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(G77), .B2(new_n281), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(G238), .B1(new_n399), .B2(new_n400), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n402), .A2(G232), .B1(G107), .B2(new_n348), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n247), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n250), .B1(new_n253), .B2(new_n217), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n439), .B2(G190), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n319), .B2(new_n439), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n395), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n382), .B1(new_n437), .B2(new_n438), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n434), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n300), .A2(new_n367), .A3(new_n425), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G97), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n392), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n251), .A2(G33), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n281), .A2(new_n449), .A3(new_n255), .A4(new_n270), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n450), .B2(new_n447), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT78), .ZN(new_n453));
  AND2_X1   g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G97), .A2(G107), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n454), .A2(new_n455), .B1(KEYINPUT77), .B2(KEYINPUT6), .ZN(new_n456));
  NOR2_X1   g0256(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(KEYINPUT6), .B2(new_n447), .ZN(new_n458));
  XNOR2_X1  g0258(.A(G97), .B(G107), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n456), .B(G20), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n272), .A2(KEYINPUT76), .A3(G77), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT76), .B1(new_n272), .B2(G77), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n346), .A2(new_n351), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n453), .B1(new_n467), .B2(new_n271), .ZN(new_n468));
  INV_X1    g0268(.A(G107), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n346), .B2(new_n351), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n460), .A2(new_n463), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n453), .B(new_n271), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n452), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT79), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n251), .B(G45), .C1(new_n246), .C2(KEYINPUT5), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT80), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n248), .A2(G1), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT80), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT81), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G274), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n256), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n477), .A2(new_n478), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT81), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n480), .A2(KEYINPUT80), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n484), .A2(new_n486), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n489), .A3(new_n491), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G257), .A3(new_n247), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n217), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n257), .A2(new_n374), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n217), .A2(G1698), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n497), .B1(new_n306), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n247), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n319), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n504), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n256), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n316), .A3(new_n492), .A4(new_n494), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n271), .B1(new_n470), .B2(new_n471), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n472), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT79), .A3(new_n452), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n476), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n493), .A2(G264), .A3(new_n247), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n493), .A2(KEYINPUT87), .A3(G264), .A4(new_n247), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G250), .B2(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n306), .A2(new_n524), .B1(new_n245), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n526), .A2(new_n256), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  AND4_X1   g0328(.A1(new_n395), .A2(new_n521), .A3(new_n492), .A4(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n527), .B1(new_n519), .B2(new_n520), .ZN(new_n530));
  AOI21_X1  g0330(.A(G169), .B1(new_n530), .B2(new_n492), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n303), .A2(new_n304), .A3(new_n274), .A4(new_n305), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT22), .B1(new_n533), .B2(new_n310), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n310), .A2(KEYINPUT22), .A3(G20), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n257), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT86), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT86), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n257), .A2(new_n538), .A3(new_n535), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(G116), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n245), .A2(new_n542), .A3(G20), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n274), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n469), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n541), .B1(new_n540), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n271), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n392), .A2(KEYINPUT25), .A3(new_n469), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT25), .B1(new_n392), .B2(new_n469), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n553), .A2(new_n554), .B1(new_n469), .B2(new_n450), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n532), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(G169), .B1(new_n495), .B2(new_n505), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n509), .A2(G179), .A3(new_n492), .A4(new_n494), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n474), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n516), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n392), .A2(new_n542), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n450), .B2(new_n542), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(G20), .B1(G33), .B2(G283), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n245), .A2(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT85), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n270), .A2(new_n255), .B1(G20), .B2(new_n542), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT20), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT85), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT85), .B1(new_n567), .B2(new_n568), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT20), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n566), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n302), .A2(G33), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n582));
  OAI21_X1  g0382(.A(G303), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n522), .A2(new_n374), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(G264), .B2(new_n374), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n306), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n256), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n493), .A2(G270), .A3(new_n247), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n490), .A2(new_n486), .A3(new_n491), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n587), .B(new_n588), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n580), .A2(new_n591), .A3(G169), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n580), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n492), .A2(G190), .A3(new_n587), .A4(new_n588), .ZN(new_n596));
  INV_X1    g0396(.A(new_n591), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n319), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(G179), .A3(new_n580), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n580), .A2(new_n591), .A3(KEYINPUT21), .A4(G169), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n594), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n530), .A2(new_n316), .A3(new_n492), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n521), .A2(new_n492), .A3(new_n528), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(G200), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n540), .A2(new_n547), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT24), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n548), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n555), .B1(new_n607), .B2(new_n271), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n217), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(G238), .B2(G1698), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n306), .A2(new_n611), .B1(new_n245), .B2(new_n542), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT83), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI221_X1 g0414(.A(KEYINPUT83), .B1(new_n245), .B2(new_n542), .C1(new_n306), .C2(new_n611), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n256), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(KEYINPUT82), .A2(G250), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n480), .A2(new_n485), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(G250), .ZN(new_n619));
  OAI22_X1  g0419(.A1(KEYINPUT82), .A2(new_n619), .B1(new_n248), .B2(G1), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n247), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT19), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n310), .A2(new_n447), .A3(new_n469), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n260), .A2(new_n274), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n623), .A2(new_n274), .A3(G33), .A4(G97), .ZN(new_n627));
  OAI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n533), .B2(new_n214), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n628), .A2(new_n271), .B1(new_n392), .B2(new_n427), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n391), .A2(new_n428), .A3(new_n449), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n622), .A2(new_n382), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n395), .A3(new_n621), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n533), .A2(new_n214), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n624), .A2(new_n625), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n627), .B1(new_n634), .B2(KEYINPUT19), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n271), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n391), .A2(KEYINPUT84), .A3(G87), .A4(new_n449), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n450), .B2(new_n310), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n427), .A2(new_n392), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n621), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n247), .B1(new_n612), .B2(new_n613), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n643), .B1(new_n644), .B2(new_n615), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n645), .B2(G190), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n622), .A2(G200), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n631), .A2(new_n632), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n601), .A2(new_n609), .A3(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n563), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n446), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT88), .Z(G372));
  NAND2_X1  g0452(.A1(new_n629), .A2(new_n630), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n632), .B(new_n653), .C1(G169), .C2(new_n645), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n616), .A2(G190), .A3(new_n621), .ZN(new_n655));
  INV_X1    g0455(.A(new_n642), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n655), .B(new_n656), .C1(new_n319), .C2(new_n645), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n608), .B2(new_n604), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n599), .A2(new_n600), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n530), .A2(new_n395), .A3(new_n492), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n603), .B2(G169), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n594), .B(new_n660), .C1(new_n662), .C2(new_n608), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n516), .A2(new_n562), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(KEYINPUT89), .B(KEYINPUT26), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n562), .A2(new_n658), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n476), .A2(new_n515), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n561), .A3(new_n648), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n446), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT90), .Z(new_n675));
  AND2_X1   g0475(.A1(new_n363), .A2(new_n365), .ZN(new_n676));
  INV_X1    g0476(.A(new_n444), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n291), .A2(new_n677), .B1(new_n298), .B2(new_n297), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n357), .A2(new_n366), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT10), .B1(new_n414), .B2(new_n416), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n421), .A2(new_n423), .A3(new_n418), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n397), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n675), .A2(new_n685), .ZN(G369));
  NAND3_X1  g0486(.A1(new_n251), .A2(new_n274), .A3(G13), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(G213), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n557), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n558), .A2(new_n609), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n693), .A2(new_n662), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT91), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT91), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n693), .A2(new_n697), .A3(new_n662), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n701));
  INV_X1    g0501(.A(new_n692), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n595), .A2(new_n702), .ZN(new_n703));
  MUX2_X1   g0503(.A(new_n601), .B(new_n701), .S(new_n703), .Z(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G330), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n558), .A2(new_n692), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n692), .B1(new_n660), .B2(new_n594), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(new_n699), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(G399));
  NOR2_X1   g0511(.A1(new_n624), .A2(G116), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n207), .A2(new_n246), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(G1), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n212), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT28), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT29), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n702), .C1(new_n666), .C2(new_n672), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT93), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT79), .B1(new_n514), .B2(new_n452), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n475), .B(new_n451), .C1(new_n513), .C2(new_n472), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n506), .A2(new_n510), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n562), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n719), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n701), .B1(new_n557), .B2(new_n532), .ZN(new_n726));
  AND4_X1   g0526(.A1(new_n316), .A2(new_n521), .A3(new_n492), .A4(new_n528), .ZN(new_n727));
  AOI21_X1  g0527(.A(G200), .B1(new_n530), .B2(new_n492), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n648), .B1(new_n729), .B2(new_n557), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n516), .A2(KEYINPUT93), .A3(new_n562), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n725), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n654), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n670), .A2(KEYINPUT26), .A3(new_n561), .A4(new_n648), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n667), .B1(new_n562), .B2(new_n658), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n692), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n718), .B1(new_n738), .B2(new_n717), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n560), .A2(new_n622), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .A3(new_n530), .A4(new_n597), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  INV_X1    g0544(.A(new_n495), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n745), .A2(new_n645), .A3(G179), .A4(new_n509), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n597), .A2(new_n530), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n745), .B2(new_n509), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n530), .A2(new_n492), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n591), .A4(new_n622), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n743), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n692), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n650), .A2(new_n702), .B1(new_n741), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT92), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n740), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n739), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n716), .B1(new_n760), .B2(G1), .ZN(G364));
  INV_X1    g0561(.A(new_n705), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n274), .A2(G13), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n251), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n713), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n704), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n257), .A2(new_n207), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n207), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n238), .A2(new_n248), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n306), .A2(new_n207), .ZN(new_n774));
  INV_X1    g0574(.A(new_n212), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(new_n248), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n772), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n255), .B1(G20), .B2(new_n382), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n767), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n274), .A2(new_n395), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR3_X1   g0586(.A1(new_n786), .A2(new_n316), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n316), .A2(new_n319), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n785), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n788), .A2(new_n327), .B1(new_n790), .B2(new_n202), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n447), .ZN(new_n796));
  NOR4_X1   g0596(.A1(new_n274), .A2(new_n319), .A3(G179), .A4(G190), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n469), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n791), .A2(new_n796), .A3(new_n348), .A4(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n786), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n789), .A2(G20), .A3(new_n395), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n216), .B1(new_n310), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n786), .A2(new_n319), .A3(G190), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G68), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n792), .A2(G20), .A3(new_n316), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(KEYINPUT94), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(KEYINPUT94), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT32), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n810), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n800), .A2(new_n806), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n803), .B(KEYINPUT95), .Z(new_n815));
  AOI21_X1  g0615(.A(new_n257), .B1(new_n815), .B2(G303), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT96), .Z(new_n817));
  INV_X1    g0617(.A(G283), .ZN(new_n818));
  INV_X1    g0618(.A(G326), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n798), .A2(new_n818), .B1(new_n819), .B2(new_n790), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n802), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G322), .C2(new_n787), .ZN(new_n823));
  INV_X1    g0623(.A(new_n810), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G329), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n794), .A2(G294), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT33), .B(G317), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT97), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n805), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n823), .A2(new_n825), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n814), .B1(new_n817), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n784), .B1(new_n832), .B2(new_n781), .ZN(new_n833));
  INV_X1    g0633(.A(new_n780), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n704), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n769), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n673), .A2(new_n702), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n434), .A2(new_n692), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n441), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n444), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n444), .A2(new_n692), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n838), .B(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n758), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n767), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n257), .B(new_n796), .C1(G294), .C2(new_n787), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n815), .A2(G107), .B1(new_n824), .B2(G311), .ZN(new_n850));
  AOI22_X1  g0650(.A1(G116), .A2(new_n801), .B1(new_n805), .B2(G283), .ZN(new_n851));
  INV_X1    g0651(.A(new_n790), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G303), .B1(G87), .B2(new_n797), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n805), .A2(G150), .B1(new_n852), .B2(G137), .ZN(new_n855));
  INV_X1    g0655(.A(G143), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n855), .B1(new_n856), .B2(new_n788), .C1(new_n811), .C2(new_n802), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  NOR2_X1   g0658(.A1(new_n798), .A2(new_n214), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n306), .B(new_n859), .C1(G58), .C2(new_n794), .ZN(new_n860));
  INV_X1    g0660(.A(new_n815), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n860), .B1(new_n202), .B2(new_n861), .C1(new_n862), .C2(new_n810), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n854), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n781), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n781), .A2(new_n778), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n766), .B(new_n765), .C1(new_n216), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n677), .B1(new_n441), .B2(new_n839), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n868), .A2(new_n842), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n865), .B(new_n867), .C1(new_n869), .C2(new_n779), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n848), .A2(new_n870), .ZN(G384));
  NAND2_X1  g0671(.A1(new_n286), .A2(new_n290), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n267), .B2(new_n268), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n298), .B(new_n692), .C1(new_n873), .C2(new_n297), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n298), .A2(new_n692), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n291), .A2(new_n299), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n844), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n665), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n601), .A2(new_n609), .A3(new_n648), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n558), .A4(new_n702), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n753), .A2(new_n741), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(new_n881), .A3(new_n755), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(new_n690), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n358), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n355), .A2(new_n362), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n358), .A2(new_n317), .A3(new_n320), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n408), .B1(new_n891), .B2(new_n343), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT98), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n342), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI211_X1 g0694(.A(KEYINPUT98), .B(new_n408), .C1(new_n891), .C2(new_n343), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n332), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(new_n361), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n886), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n889), .B1(new_n899), .B2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n367), .A2(new_n886), .A3(new_n896), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n885), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT99), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n897), .B2(new_n898), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT38), .B(new_n901), .C1(new_n906), .C2(new_n889), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n904), .B1(new_n903), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n884), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n887), .B1(new_n679), .B2(new_n676), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n888), .B(new_n905), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n885), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n907), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n877), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n911), .A2(new_n912), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n882), .A2(new_n446), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n921), .A3(new_n740), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n874), .A2(new_n876), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n702), .B(new_n869), .C1(new_n666), .C2(new_n672), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n843), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n923), .B(new_n925), .C1(new_n909), .C2(new_n910), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n903), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n297), .A2(new_n298), .A3(new_n702), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n676), .A2(new_n886), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n926), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n739), .A2(new_n446), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n685), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n922), .A2(new_n937), .B1(new_n251), .B2(new_n763), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n922), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n210), .A2(new_n542), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT35), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT36), .ZN(new_n945));
  OR3_X1    g0745(.A1(new_n212), .A2(new_n216), .A3(new_n333), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n202), .A2(G68), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n251), .B(G13), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n939), .A2(new_n945), .A3(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n656), .A2(new_n702), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT100), .B1(new_n734), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n658), .B2(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n734), .A2(KEYINPUT100), .A3(new_n950), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(KEYINPUT43), .A3(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT103), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n723), .A2(new_n719), .A3(new_n724), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT93), .B1(new_n516), .B2(new_n562), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n702), .B1(new_n476), .B2(new_n515), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n670), .A2(new_n561), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n692), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n699), .A2(new_n709), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n956), .B1(new_n968), .B2(KEYINPUT42), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT42), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n965), .A2(new_n967), .A3(KEYINPUT103), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n959), .A2(new_n961), .B1(new_n963), .B2(new_n692), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n562), .B1(new_n973), .B2(new_n558), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n974), .A2(new_n702), .B1(new_n968), .B2(KEYINPUT42), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n955), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT102), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n952), .A2(new_n953), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT101), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(KEYINPUT101), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n976), .A2(new_n977), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n978), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n976), .A2(new_n977), .ZN(new_n987));
  AOI211_X1 g0787(.A(KEYINPUT102), .B(new_n955), .C1(new_n972), .C2(new_n975), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n707), .A2(new_n973), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT104), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n989), .ZN(new_n993));
  INV_X1    g0793(.A(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT104), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n986), .A2(new_n989), .A3(new_n996), .A4(new_n990), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n699), .B(new_n709), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(new_n762), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n760), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n710), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n973), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n965), .A2(new_n710), .A3(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n973), .A3(KEYINPUT44), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n965), .B2(new_n710), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n706), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1006), .A2(new_n1010), .A3(new_n707), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1001), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n760), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n713), .B(KEYINPUT41), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n764), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n992), .A2(new_n995), .A3(new_n997), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n805), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n1020), .A2(new_n811), .B1(new_n790), .B2(new_n856), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n348), .B(new_n1021), .C1(G50), .C2(new_n801), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n795), .A2(new_n214), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n824), .A2(G137), .ZN(new_n1025));
  INV_X1    g0825(.A(G150), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n788), .A2(new_n1026), .B1(new_n216), .B2(new_n798), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n803), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1027), .B1(G58), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(G303), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n788), .A2(new_n1031), .B1(new_n790), .B2(new_n821), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT105), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n815), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(KEYINPUT105), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n1020), .A2(new_n525), .B1(new_n447), .B2(new_n798), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G283), .B2(new_n801), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT46), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n803), .B2(new_n542), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G107), .B2(new_n794), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n824), .A2(G317), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1030), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT47), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n781), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n979), .A2(new_n780), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n782), .B1(new_n207), .B2(new_n427), .C1(new_n234), .C2(new_n774), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1047), .A2(new_n767), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1019), .A2(new_n1050), .ZN(G387));
  OR2_X1    g0851(.A1(new_n760), .A2(new_n999), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1052), .A2(new_n766), .A3(new_n1000), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n700), .A2(new_n780), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n770), .A2(new_n712), .B1(G107), .B2(new_n207), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n231), .A2(new_n248), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n712), .ZN(new_n1057));
  AOI211_X1 g0857(.A(G45), .B(new_n1057), .C1(G68), .C2(G77), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n322), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n774), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1055), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n767), .B1(new_n1062), .B2(new_n783), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n802), .A2(new_n214), .B1(new_n447), .B2(new_n798), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n306), .B(new_n1064), .C1(new_n428), .C2(new_n794), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n330), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n805), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n824), .A2(G150), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n790), .A2(new_n811), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n803), .A2(new_n216), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G50), .C2(new_n787), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1041), .B1(G116), .B2(new_n797), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n805), .A2(G311), .B1(new_n852), .B2(G322), .ZN(new_n1074));
  INV_X1    g0874(.A(G317), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1031), .B2(new_n802), .C1(new_n1075), .C2(new_n788), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT106), .Z(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1028), .A2(G294), .B1(new_n794), .B2(G283), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT49), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1073), .B1(new_n819), .B2(new_n810), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1072), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1063), .B1(new_n1086), .B2(new_n781), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n999), .A2(new_n765), .B1(new_n1054), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1053), .A2(new_n1088), .ZN(G393));
  INV_X1    g0889(.A(KEYINPUT107), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n1013), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1091), .B1(new_n1092), .B2(KEYINPUT107), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n766), .B(new_n1014), .C1(new_n1093), .C2(new_n1001), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n765), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n243), .A2(new_n774), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n782), .B1(new_n447), .B2(new_n207), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n767), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n802), .A2(new_n322), .B1(new_n310), .B2(new_n798), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n1020), .A2(new_n202), .B1(new_n214), .B2(new_n803), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n795), .A2(new_n216), .ZN(new_n1101));
  OR4_X1    g0901(.A1(new_n306), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n787), .A2(G159), .B1(new_n852), .B2(G150), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n856), .B2(new_n810), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n257), .B(new_n799), .C1(G116), .C2(new_n794), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G294), .A2(new_n801), .B1(new_n805), .B2(G303), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n818), .C2(new_n803), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n788), .A2(new_n821), .B1(new_n790), .B2(new_n1075), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1110), .A2(new_n1112), .B1(new_n824), .B2(G322), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n1102), .A2(new_n1106), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1098), .B1(new_n1115), .B2(new_n781), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n965), .B2(new_n834), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1094), .A2(new_n1095), .A3(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(KEYINPUT110), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n692), .B(new_n868), .C1(new_n733), .C2(new_n737), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n842), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n733), .A2(new_n737), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1122), .A2(new_n702), .A3(new_n841), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1123), .A2(KEYINPUT110), .A3(new_n843), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1121), .A2(new_n923), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n916), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n931), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n925), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n923), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n930), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n928), .A2(new_n929), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n758), .A2(new_n869), .A3(new_n923), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1128), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1125), .A2(new_n1127), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n877), .A2(new_n882), .A3(G330), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n446), .A2(new_n882), .A3(G330), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n935), .A2(new_n1140), .A3(new_n685), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n882), .A2(G330), .A3(new_n869), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n1130), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1120), .A2(new_n1119), .A3(new_n842), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT110), .B1(new_n1123), .B2(new_n843), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1134), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n923), .B1(new_n758), .B2(new_n869), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n925), .B1(new_n1147), .B2(new_n1137), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1141), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1139), .A2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1135), .B(new_n1149), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n766), .A3(new_n1152), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1139), .A2(new_n764), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n866), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n767), .B1(new_n1066), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1101), .B1(G116), .B2(new_n787), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT111), .Z(new_n1158));
  OAI22_X1  g0958(.A1(new_n1020), .A2(new_n469), .B1(new_n802), .B2(new_n447), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G283), .B2(new_n852), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n859), .A2(new_n257), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n815), .A2(G87), .B1(new_n824), .B2(G294), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI22_X1  g0964(.A1(new_n1164), .A2(new_n801), .B1(new_n787), .B2(G132), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n257), .B1(new_n790), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G159), .B2(new_n794), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n805), .A2(G137), .B1(G50), .B2(new_n797), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1165), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n803), .A2(new_n1026), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  INV_X1    g0972(.A(G125), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n810), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1158), .A2(new_n1163), .B1(new_n1170), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1156), .B1(new_n1175), .B2(new_n781), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1132), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n779), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1153), .A2(new_n1154), .A3(new_n1178), .ZN(G378));
  OAI21_X1  g0979(.A(new_n767), .B1(new_n1155), .B2(G50), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT114), .Z(new_n1181));
  NAND2_X1  g0981(.A1(new_n797), .A2(G58), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT112), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n787), .A2(G107), .B1(new_n852), .B2(G116), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n428), .A2(new_n801), .B1(new_n805), .B2(G97), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1023), .A2(new_n1070), .A3(G41), .A4(new_n1041), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n818), .C2(new_n810), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT113), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n824), .A2(G124), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n245), .B(new_n246), .C1(new_n798), .C2(new_n811), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n788), .A2(new_n1166), .B1(new_n790), .B2(new_n1173), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G137), .B2(new_n801), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n805), .A2(G132), .B1(new_n1028), .B2(new_n1164), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(new_n1197), .C1(new_n1026), .C2(new_n795), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1193), .B(new_n1194), .C1(new_n1198), .C2(KEYINPUT59), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n246), .B1(new_n306), .B2(new_n245), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1199), .A2(new_n1200), .B1(new_n202), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1191), .A2(new_n1192), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1181), .B1(new_n1203), .B2(new_n781), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n690), .B1(new_n388), .B2(new_n393), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n684), .B2(new_n398), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n397), .B(new_n1207), .C1(new_n682), .C2(new_n683), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(new_n1210), .A3(KEYINPUT115), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT115), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n425), .A2(new_n1207), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n684), .A2(new_n398), .A3(new_n1208), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1206), .B1(new_n1211), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(KEYINPUT115), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1205), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1216), .A2(KEYINPUT116), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT116), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1204), .B1(new_n1222), .B2(new_n779), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT117), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n740), .B1(new_n917), .B2(new_n916), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n889), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n896), .A2(new_n361), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n898), .A2(new_n1227), .A3(new_n355), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1226), .B1(new_n1228), .B2(new_n905), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT38), .B1(new_n1229), .B2(new_n901), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n907), .ZN(new_n1231));
  OAI21_X1  g1031(.A(KEYINPUT99), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n883), .B1(new_n1232), .B2(new_n908), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1222), .B(new_n1225), .C1(new_n1233), .C2(KEYINPUT40), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n877), .A2(new_n882), .A3(KEYINPUT40), .ZN(new_n1235));
  OAI21_X1  g1035(.A(G330), .B1(new_n1235), .B2(new_n1126), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(new_n911), .B2(new_n912), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1234), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n934), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT118), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT118), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1239), .A2(new_n1240), .A3(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n934), .B(new_n1234), .C1(new_n1238), .C2(new_n1237), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT119), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1242), .B(new_n1244), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1224), .B1(new_n1249), .B2(new_n765), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT120), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1141), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1152), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .A4(KEYINPUT57), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT57), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1152), .B2(new_n1252), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1251), .B1(new_n1257), .B2(new_n1254), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n766), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1253), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1250), .B1(new_n1259), .B2(new_n1260), .ZN(G375));
  NAND2_X1  g1061(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1141), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1016), .A3(new_n1150), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1130), .A2(new_n778), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n861), .A2(new_n447), .B1(new_n1031), .B2(new_n810), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n788), .A2(new_n818), .B1(new_n802), .B2(new_n469), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1020), .A2(new_n542), .B1(new_n790), .B2(new_n525), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n348), .B1(new_n798), .B2(new_n216), .C1(new_n427), .C2(new_n795), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n861), .A2(new_n811), .B1(new_n1166), .B2(new_n810), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1164), .A2(new_n805), .B1(new_n787), .B2(G137), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n306), .B1(G50), .B2(new_n794), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n1026), .C2(new_n802), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n790), .A2(new_n862), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT121), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1183), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1272), .A2(new_n1275), .A3(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n781), .B1(new_n1271), .B2(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1280), .B(new_n767), .C1(G68), .C2(new_n1155), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT122), .Z(new_n1282));
  AOI22_X1  g1082(.A1(new_n1262), .A2(new_n765), .B1(new_n1266), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1265), .A2(new_n1283), .ZN(G381));
  NAND3_X1  g1084(.A1(new_n1053), .A2(new_n836), .A3(new_n1088), .ZN(new_n1285));
  OR4_X1    g1085(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1285), .ZN(new_n1286));
  OR4_X1    g1086(.A1(G387), .A2(new_n1286), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  INV_X1    g1088(.A(G213), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1289), .A2(G343), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  OAI211_X1 g1092(.A(G378), .B(new_n1250), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1249), .A2(new_n1016), .A3(new_n1253), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1224), .B1(new_n1254), .B2(new_n765), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1288), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1290), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1264), .B1(new_n1300), .B2(new_n1149), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1263), .A2(KEYINPUT60), .A3(new_n1141), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n766), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1283), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n848), .A3(new_n870), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(G384), .A3(new_n1283), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(new_n1299), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT123), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1290), .B1(new_n1293), .B2(new_n1297), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT123), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n1308), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1310), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT124), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1310), .A2(new_n1317), .A3(new_n1311), .A4(new_n1314), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G393), .A2(G396), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(G390), .A2(new_n1285), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1285), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1321), .A2(new_n1094), .A3(new_n1095), .A4(new_n1117), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G387), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1019), .A2(new_n1320), .A3(new_n1322), .A4(new_n1050), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1290), .A2(G2897), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1307), .B(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1327), .B1(new_n1330), .B2(new_n1312), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1312), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1308), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1316), .A2(new_n1318), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1338), .B(new_n1339), .C1(new_n1312), .C2(new_n1330), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT62), .B1(new_n1310), .B2(new_n1314), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1337), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1336), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT127), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1336), .A2(KEYINPUT127), .A3(new_n1342), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1288), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1293), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1308), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(new_n1337), .ZN(G402));
endmodule


