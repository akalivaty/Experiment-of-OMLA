//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n474), .B2(new_n461), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(KEYINPUT65), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n469), .B1(new_n475), .B2(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT67), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n481));
  INV_X1    g056(.A(new_n467), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OAI21_X1  g058(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  XNOR2_X1  g063(.A(KEYINPUT68), .B(G114), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n461), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G126), .ZN(new_n492));
  OAI22_X1  g067(.A1(new_n490), .A2(new_n491), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n493), .A2(new_n494), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n471), .A2(new_n461), .ZN(new_n500));
  INV_X1    g075(.A(G138), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n496), .A2(new_n497), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT71), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n508), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  AOI211_X1 g089(.A(KEYINPUT71), .B(new_n514), .C1(new_n509), .C2(new_n511), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n506), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n514), .B2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT70), .B(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(new_n514), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n512), .A2(new_n523), .A3(KEYINPUT5), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G88), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n522), .A2(new_n507), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n529), .B1(G50), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n519), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G89), .Z(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n526), .A2(new_n527), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n530), .A2(G51), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT74), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n516), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT75), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT75), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n548), .B(new_n544), .C1(new_n516), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(G651), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n528), .A2(G90), .B1(G52), .B2(new_n530), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n528), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n530), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n516), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n560));
  INV_X1    g135(.A(G651), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n559), .B2(KEYINPUT76), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n556), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n530), .A2(G53), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n571), .A2(new_n572), .B1(G91), .B2(new_n528), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT78), .B1(new_n513), .B2(new_n515), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n526), .A2(new_n527), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g151(.A(KEYINPUT79), .B(G65), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT80), .B1(new_n580), .B2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  AOI211_X1 g157(.A(new_n582), .B(new_n561), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n573), .B1(new_n581), .B2(new_n583), .ZN(G299));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n542), .B(new_n585), .ZN(G286));
  OAI21_X1  g161(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n528), .A2(G87), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n530), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT81), .Z(G288));
  AOI22_X1  g166(.A1(new_n536), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n561), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n530), .A2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT82), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n530), .A2(new_n596), .A3(G48), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n595), .A2(new_n597), .B1(new_n528), .B2(G86), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n528), .A2(G85), .B1(G47), .B2(new_n530), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n561), .B2(new_n601), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT83), .Z(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n530), .A2(G54), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n528), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT10), .B1(new_n528), .B2(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT85), .B(G66), .Z(new_n609));
  NAND3_X1  g184(.A1(new_n574), .A2(new_n576), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(G79), .A2(G543), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT84), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n561), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n604), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n604), .B1(G868), .B2(new_n614), .ZN(G321));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G286), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(G297));
  XNOR2_X1  g196(.A(new_n620), .B(KEYINPUT86), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(new_n563), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n618), .ZN(new_n626));
  INV_X1    g201(.A(new_n614), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n626), .B1(new_n628), .B2(new_n618), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n485), .A2(G123), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT87), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n482), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n461), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n500), .A2(G2104), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT12), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT12), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n500), .A2(new_n640), .A3(G2104), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n637), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT90), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT89), .B(KEYINPUT14), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2451), .B(G2454), .Z(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT91), .ZN(new_n662));
  INV_X1    g237(.A(G14), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT92), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n668), .A2(new_n669), .ZN(new_n672));
  AOI21_X1  g247(.A(KEYINPUT18), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G2100), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n670), .B2(KEYINPUT18), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(G2096), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n674), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1971), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n697), .A2(G23), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n590), .B(KEYINPUT93), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G16), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n700), .A2(new_n701), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n701), .B2(new_n700), .ZN(new_n707));
  MUX2_X1   g282(.A(G6), .B(G305), .S(G16), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(new_n702), .B2(new_n705), .ZN(new_n711));
  OR3_X1    g286(.A1(new_n707), .A2(KEYINPUT34), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT34), .B1(new_n707), .B2(new_n711), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n697), .A2(G24), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G290), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n716), .A2(G1986), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(G1986), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n485), .A2(G119), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n461), .A2(G107), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G25), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n717), .A2(new_n718), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n712), .A2(new_n713), .A3(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT36), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n697), .A2(G4), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n614), .B2(new_n697), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT95), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G1348), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n697), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n563), .B2(new_n697), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1341), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n733), .A2(G1348), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G32), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n741));
  INV_X1    g316(.A(G129), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n484), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NOR2_X1   g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT99), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  OR4_X1    g326(.A1(new_n734), .A2(new_n737), .A3(new_n738), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT31), .B(G11), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT101), .ZN(new_n754));
  INV_X1    g329(.A(G28), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT30), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT30), .B2(new_n755), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n757), .C1(new_n636), .C2(new_n739), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT24), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G160), .B2(new_n739), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(G2084), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n739), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n739), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT29), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n765), .B1(G2090), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n739), .A2(G33), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(new_n461), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT97), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n776));
  NAND2_X1  g351(.A1(G103), .A2(G2104), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n482), .A2(G139), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n774), .A2(new_n775), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n771), .B1(new_n781), .B2(G29), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n782), .A2(new_n442), .B1(new_n764), .B2(G2084), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n770), .B(new_n783), .C1(new_n442), .C2(new_n782), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n739), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n485), .A2(G128), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n482), .A2(G140), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n461), .A2(G116), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G29), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(KEYINPUT96), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n697), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n697), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n769), .A2(G2090), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT102), .ZN(new_n801));
  OAI221_X1 g376(.A(new_n797), .B1(G1966), .B2(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n739), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n739), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n443), .ZN(new_n805));
  INV_X1    g380(.A(new_n800), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(KEYINPUT102), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n784), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n697), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n617), .B2(new_n697), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n799), .A2(G1966), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n697), .A2(G5), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G171), .B2(new_n697), .ZN(new_n817));
  INV_X1    g392(.A(G1961), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n808), .A2(new_n813), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n730), .A2(new_n752), .A3(new_n820), .ZN(G311));
  OR3_X1    g396(.A1(new_n730), .A2(new_n752), .A3(new_n820), .ZN(G150));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n526), .B2(new_n527), .ZN(new_n824));
  AND2_X1   g399(.A1(G80), .A2(G543), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n824), .A2(KEYINPUT103), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT103), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(G651), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n528), .A2(G93), .B1(G55), .B2(new_n530), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n625), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n563), .A2(new_n828), .A3(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NOR2_X1   g411(.A1(new_n627), .A2(new_n623), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(new_n830), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT104), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n847), .ZN(G145));
  NAND2_X1  g423(.A1(new_n482), .A2(G142), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n485), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n461), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n642), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n723), .ZN(new_n855));
  AOI22_X1  g430(.A1(new_n500), .A2(new_n502), .B1(KEYINPUT4), .B2(new_n498), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(new_n493), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n855), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n791), .B(KEYINPUT105), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n781), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n747), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n859), .A2(new_n862), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(G162), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n636), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g446(.A(new_n835), .B(new_n628), .ZN(new_n872));
  NAND2_X1  g447(.A1(G299), .A2(new_n627), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n614), .B(new_n573), .C1(new_n581), .C2(new_n583), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n876), .A3(new_n874), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(KEYINPUT106), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n873), .A2(new_n876), .A3(new_n874), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n881), .B2(KEYINPUT106), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n875), .B1(new_n883), .B2(new_n872), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(G303), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n704), .B(G305), .Z(new_n888));
  XOR2_X1   g463(.A(new_n887), .B(new_n888), .Z(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n884), .A2(new_n885), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n886), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n886), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n845), .A2(new_n618), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(G295));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n895), .ZN(G331));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  NAND3_X1  g473(.A1(G168), .A2(new_n550), .A3(new_n551), .ZN(new_n899));
  NAND2_X1  g474(.A1(G286), .A2(G301), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n563), .B1(new_n843), .B2(new_n844), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n625), .A2(new_n842), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n833), .A2(new_n834), .A3(new_n900), .A4(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n898), .B1(new_n882), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n561), .B1(new_n578), .B2(new_n579), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT80), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n614), .B1(new_n909), .B2(new_n573), .ZN(new_n910));
  NOR2_X1   g485(.A1(G299), .A2(new_n627), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n877), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n877), .A2(KEYINPUT106), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n913), .A2(new_n914), .A3(new_n898), .A4(new_n906), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n904), .A2(new_n905), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n873), .A3(new_n874), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n890), .B1(new_n907), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n906), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT107), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n921), .A2(new_n889), .A3(new_n917), .A4(new_n915), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n869), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT43), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n917), .B1(new_n881), .B2(new_n916), .ZN(new_n927));
  AOI21_X1  g502(.A(G37), .B1(new_n890), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n921), .A2(new_n917), .A3(new_n915), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n933), .B2(new_n890), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n922), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n932), .B1(new_n939), .B2(new_n940), .ZN(G397));
  AND2_X1   g516(.A1(G160), .A2(G40), .ZN(new_n942));
  XOR2_X1   g517(.A(KEYINPUT109), .B(G1384), .Z(new_n943));
  NAND3_X1  g518(.A1(new_n858), .A2(KEYINPUT45), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT45), .B1(new_n504), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(KEYINPUT56), .B(G2072), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT50), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n504), .A2(new_n951), .A3(new_n946), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n857), .A2(G1384), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT50), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(new_n955), .A3(new_n942), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT119), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n956), .A2(new_n957), .A3(new_n812), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n957), .B1(new_n956), .B2(new_n812), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT57), .ZN(new_n961));
  XNOR2_X1  g536(.A(G299), .B(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G160), .A2(G40), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(new_n951), .B2(new_n953), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n504), .A2(new_n946), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1348), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n965), .A2(new_n954), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n969), .A2(new_n970), .B1(new_n796), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n964), .B1(new_n627), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n956), .A2(new_n812), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT119), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n956), .A2(new_n957), .A3(new_n812), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(new_n962), .A3(new_n950), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n964), .A2(new_n978), .A3(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT120), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n971), .A2(new_n796), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n966), .A2(new_n968), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n982), .B(KEYINPUT60), .C1(new_n983), .C2(G1348), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT121), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n627), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n972), .A2(KEYINPUT60), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n614), .B(KEYINPUT121), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n984), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT122), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n964), .A2(new_n978), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT61), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n990), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT122), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n986), .A4(new_n987), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n945), .A2(new_n948), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G1996), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT58), .B(G1341), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n971), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n563), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT59), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n991), .A2(new_n994), .A3(new_n997), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n979), .B1(new_n981), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n998), .B2(G2078), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n969), .A2(new_n818), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n942), .B(KEYINPUT116), .C1(KEYINPUT45), .C2(new_n953), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n953), .A2(KEYINPUT45), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n965), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1006), .A2(G2078), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1007), .A2(new_n1008), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G171), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT124), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT124), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1019), .A3(G171), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n858), .A2(new_n943), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1014), .A2(G40), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n476), .A2(new_n469), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n944), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n942), .A2(new_n944), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1026), .A2(new_n947), .A3(G2078), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1008), .B(new_n1025), .C1(KEYINPUT53), .C2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1028), .A2(G171), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1018), .A2(new_n1020), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1026), .B2(new_n947), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n969), .B2(G2090), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G166), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT111), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1035), .A2(new_n1043), .A3(G8), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1034), .B1(G2090), .B2(new_n956), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(G8), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n598), .A2(KEYINPUT112), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n598), .A2(KEYINPUT112), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n593), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(G1981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT114), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT113), .B1(G305), .B2(G1981), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1050), .B2(G1981), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT49), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1054), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(G1981), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT49), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(KEYINPUT114), .A3(new_n1060), .A4(new_n1052), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n971), .A2(new_n1036), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n1064));
  INV_X1    g639(.A(new_n704), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(new_n1062), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1066), .A2(new_n1062), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1047), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1031), .B1(new_n1028), .B2(G171), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1007), .A2(G301), .A3(new_n1008), .A4(new_n1015), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1009), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1078));
  INV_X1    g653(.A(G1966), .ZN(new_n1079));
  INV_X1    g654(.A(G2084), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1078), .A2(new_n1079), .B1(new_n983), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1077), .B1(new_n1081), .B2(new_n1036), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT51), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n983), .A2(new_n1080), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(G8), .B1(new_n1086), .B2(G286), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1083), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1081), .A2(G168), .ZN(new_n1090));
  OAI211_X1 g665(.A(KEYINPUT51), .B(new_n1082), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1032), .A2(new_n1076), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1005), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1063), .A2(new_n1071), .A3(new_n1044), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G305), .A2(G1981), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G288), .A2(G1976), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1097), .B1(new_n1063), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1062), .B1(new_n1099), .B2(KEYINPUT115), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1036), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1035), .A2(new_n1043), .A3(G8), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT63), .A4(G168), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1035), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1043), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1063), .A2(new_n1071), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n1109), .B2(KEYINPUT117), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1063), .A2(new_n1071), .A3(new_n1108), .A4(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1081), .A2(new_n1036), .A3(G286), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1047), .A2(new_n1063), .A3(new_n1071), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1110), .A2(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1095), .B1(new_n1102), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1109), .A2(KEYINPUT117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1105), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1112), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1099), .A2(KEYINPUT115), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1062), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1122), .A2(new_n1125), .A3(KEYINPUT118), .A4(new_n1096), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1092), .A2(KEYINPUT62), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1089), .A2(new_n1091), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1072), .B1(new_n1020), .B2(new_n1018), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1094), .A2(new_n1117), .A3(new_n1126), .A4(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1022), .A2(new_n965), .ZN(new_n1133));
  INV_X1    g708(.A(G1996), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n747), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n791), .B(new_n796), .ZN(new_n1136));
  OAI21_X1  g711(.A(G1996), .B1(new_n743), .B2(new_n746), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(new_n1139), .B(KEYINPUT110), .Z(new_n1140));
  INV_X1    g715(.A(new_n1133), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n723), .B(new_n725), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(G290), .B(G1986), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1133), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1132), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n723), .A2(new_n726), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1140), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n791), .A2(G2067), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1141), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  XOR2_X1   g725(.A(new_n1150), .B(KEYINPUT125), .Z(new_n1151));
  NAND2_X1  g726(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT46), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT126), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1136), .A2(new_n747), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1152), .A2(new_n1153), .B1(new_n1133), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1141), .A2(G290), .A3(G1986), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT48), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1159), .B1(new_n1143), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1151), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1146), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n1166));
  INV_X1    g740(.A(G319), .ZN(new_n1167));
  NOR3_X1   g741(.A1(G229), .A2(new_n1167), .A3(G227), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n870), .A2(new_n1168), .A3(new_n665), .ZN(new_n1169));
  INV_X1    g743(.A(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n930), .B2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g745(.A(KEYINPUT127), .B(new_n1169), .C1(new_n924), .C2(new_n929), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1171), .A2(new_n1172), .ZN(G308));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n1170), .ZN(G225));
endmodule


