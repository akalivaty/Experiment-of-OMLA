//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n202), .A2(new_n203), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n214), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n213), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n214), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT64), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n222), .B(new_n226), .C1(KEYINPUT1), .C2(new_n221), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G68), .B(G77), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G50), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G58), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(new_n203), .A2(G20), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n211), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g0047(.A(KEYINPUT70), .B1(new_n246), .B2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT70), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(new_n211), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI221_X1 g0052(.A(new_n245), .B1(new_n201), .B2(new_n247), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n214), .B2(new_n246), .ZN(new_n255));
  NAND4_X1  g0055(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n255), .A2(new_n210), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT11), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n245), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT12), .Z(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n257), .B1(new_n265), .B2(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n259), .B(new_n264), .C1(new_n203), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n210), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G41), .A2(G45), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G238), .ZN(new_n276));
  OAI21_X1  g0076(.A(KEYINPUT67), .B1(new_n273), .B2(G1), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n278), .B(new_n265), .C1(G41), .C2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(G274), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n269), .B2(new_n270), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(new_n280), .B2(new_n283), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n276), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT75), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT13), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n276), .B(new_n289), .C1(new_n284), .C2(new_n285), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  OAI211_X1 g0092(.A(G232), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  OAI211_X1 g0094(.A(G226), .B(new_n294), .C1(new_n291), .C2(new_n292), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G97), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n272), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT74), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT74), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(new_n300), .A3(new_n272), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n287), .A2(new_n288), .A3(new_n290), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT76), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n286), .A2(KEYINPUT75), .B1(new_n299), .B2(new_n301), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n306), .A2(KEYINPUT76), .A3(new_n288), .A4(new_n290), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n287), .A2(new_n290), .A3(new_n302), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT13), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(G169), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT77), .ZN(new_n313));
  AND4_X1   g0113(.A1(new_n313), .A2(new_n287), .A3(new_n290), .A4(new_n302), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n306), .B2(new_n290), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT13), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n303), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n311), .B1(new_n310), .B2(G169), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n268), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n268), .B1(new_n310), .B2(G200), .ZN(new_n324));
  INV_X1    g0124(.A(G190), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n316), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(new_n316), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G20), .A2(G33), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(KEYINPUT8), .B(G58), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n251), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n257), .ZN(new_n337));
  XOR2_X1   g0137(.A(new_n337), .B(KEYINPUT71), .Z(new_n338));
  NAND2_X1  g0138(.A1(new_n261), .A2(G20), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G50), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n266), .B2(G50), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n285), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(G226), .B2(new_n275), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n246), .ZN(new_n347));
  NAND2_X1  g0147(.A1(KEYINPUT3), .A2(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n294), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G223), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  INV_X1    g0151(.A(G222), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n294), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n350), .B1(new_n252), .B2(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n272), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n345), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n356), .A2(new_n318), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n345), .B2(new_n355), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n342), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g0160(.A(new_n360), .B(KEYINPUT72), .Z(new_n361));
  INV_X1    g0161(.A(KEYINPUT9), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n342), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n345), .B2(new_n355), .ZN(new_n365));
  INV_X1    g0165(.A(new_n356), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(G190), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n338), .A2(KEYINPUT9), .A3(new_n341), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n363), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT10), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n363), .A2(new_n371), .A3(new_n367), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n343), .A2(new_n344), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n275), .A2(G244), .ZN(new_n375));
  INV_X1    g0175(.A(G232), .ZN(new_n376));
  INV_X1    g0176(.A(G107), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n353), .A2(new_n376), .B1(new_n377), .B2(new_n351), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(G238), .B2(new_n349), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n374), .B(new_n375), .C1(new_n379), .C2(new_n271), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n364), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(G190), .B2(new_n380), .ZN(new_n382));
  INV_X1    g0182(.A(new_n335), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n387), .B1(new_n211), .B2(new_n252), .C1(new_n251), .C2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(new_n257), .ZN(new_n390));
  INV_X1    g0190(.A(new_n339), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n252), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n267), .B2(new_n252), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n394), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n380), .A2(G169), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n380), .A2(new_n318), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n361), .A2(new_n373), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n339), .A2(new_n335), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n266), .B2(new_n335), .ZN(new_n404));
  INV_X1    g0204(.A(new_n257), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n351), .B2(G20), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n291), .A2(new_n292), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n203), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT79), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n207), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G20), .ZN(new_n416));
  INV_X1    g0216(.A(G159), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT80), .B1(new_n247), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT80), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n333), .A2(new_n419), .A3(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT16), .B1(new_n410), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT7), .B1(new_n408), .B2(new_n211), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n291), .A2(new_n292), .A3(new_n406), .A4(G20), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT16), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n415), .A2(G20), .B1(new_n418), .B2(new_n420), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n405), .B1(new_n423), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n404), .B1(new_n430), .B2(KEYINPUT81), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n410), .A2(new_n422), .A3(KEYINPUT16), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n257), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT81), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G223), .B(new_n294), .C1(new_n291), .C2(new_n292), .ZN(new_n438));
  OAI211_X1 g0238(.A(G226), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n439));
  INV_X1    g0239(.A(G87), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n438), .B(new_n439), .C1(new_n246), .C2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT82), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n272), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n441), .B2(new_n272), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n343), .A2(new_n344), .B1(G232), .B2(new_n275), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(KEYINPUT83), .A3(new_n318), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n441), .A2(new_n272), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n443), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n275), .A2(G232), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n318), .C1(new_n284), .C2(new_n285), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n449), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n450), .B(new_n453), .C1(new_n284), .C2(new_n285), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n358), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT18), .B1(new_n437), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n456), .A2(new_n364), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n447), .A2(new_n325), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n452), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n462), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n448), .A2(new_n455), .A3(new_n457), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n434), .A2(new_n435), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n404), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT18), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n404), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT17), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n459), .A2(new_n463), .A3(new_n469), .A4(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n402), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n332), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT91), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n294), .C1(new_n291), .C2(new_n292), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n347), .A2(G303), .A3(new_n348), .ZN(new_n478));
  OAI211_X1 g0278(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT90), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT90), .B1(new_n349), .B2(G264), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n272), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n271), .ZN(new_n489));
  INV_X1    g0289(.A(G270), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT89), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT89), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(G270), .A4(new_n271), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n283), .A2(new_n485), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND4_X1   g0296(.A1(new_n476), .A2(new_n483), .A3(new_n491), .A4(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n494), .A2(new_n485), .B1(new_n269), .B2(new_n270), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n492), .B1(new_n498), .B2(G270), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(new_n495), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n476), .B1(new_n501), .B2(new_n483), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n497), .A2(new_n502), .A3(new_n358), .ZN(new_n503));
  INV_X1    g0303(.A(G283), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n246), .A2(new_n504), .ZN(new_n505));
  AOI211_X1 g0305(.A(G20), .B(new_n505), .C1(new_n246), .C2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n257), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT92), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT92), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n257), .A2(new_n511), .A3(new_n508), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n506), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT20), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n515), .B(new_n506), .C1(new_n510), .C2(new_n512), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n391), .A2(G116), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n339), .B1(G1), .B2(new_n246), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n257), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n507), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n514), .A2(new_n516), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT21), .B1(new_n503), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n325), .B1(new_n497), .B2(new_n502), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n479), .A2(new_n480), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n477), .A2(new_n478), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n482), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n271), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n491), .A2(new_n495), .A3(new_n493), .ZN(new_n529));
  OAI21_X1  g0329(.A(KEYINPUT91), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n501), .A2(new_n476), .A3(new_n483), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n364), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n521), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n520), .A2(new_n517), .ZN(new_n534));
  INV_X1    g0334(.A(new_n506), .ZN(new_n535));
  INV_X1    g0335(.A(new_n512), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n511), .B1(new_n257), .B2(new_n508), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n530), .A2(KEYINPUT21), .A3(G169), .A4(new_n531), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n483), .A2(G179), .A3(new_n496), .A4(new_n491), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n522), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n505), .B1(new_n349), .B2(G250), .ZN(new_n546));
  OAI211_X1 g0346(.A(G244), .B(new_n294), .C1(new_n291), .C2(new_n292), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT4), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(KEYINPUT4), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n547), .B2(new_n549), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n272), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n498), .A2(G257), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n495), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  INV_X1    g0359(.A(G97), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n559), .A2(new_n560), .A3(G107), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n563), .A2(new_n211), .B1(new_n252), .B2(new_n247), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n377), .B1(new_n407), .B2(new_n409), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n257), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n339), .A2(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(new_n519), .B2(G97), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n558), .A2(new_n358), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n554), .A2(KEYINPUT85), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(new_n272), .C1(new_n552), .C2(new_n553), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n570), .A2(new_n318), .A3(new_n572), .A4(new_n557), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n556), .B1(new_n554), .B2(KEYINPUT85), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n364), .B1(new_n576), .B2(new_n572), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n566), .B(new_n568), .C1(new_n558), .C2(new_n325), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT86), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n577), .B2(new_n579), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n575), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n498), .A2(G264), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT94), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G33), .A2(G294), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G250), .B(new_n294), .C1(new_n291), .C2(new_n292), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n590), .A2(new_n587), .A3(new_n586), .A4(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n272), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n495), .B(new_n585), .C1(new_n591), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n364), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G190), .B2(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n519), .A2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n261), .A2(G20), .A3(new_n377), .ZN(new_n598));
  XOR2_X1   g0398(.A(new_n598), .B(KEYINPUT25), .Z(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n351), .A2(new_n211), .A3(G87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT22), .ZN(new_n602));
  AOI21_X1  g0402(.A(G20), .B1(new_n347), .B2(new_n348), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT93), .B1(new_n377), .B2(G20), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G116), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n607), .A2(KEYINPUT23), .B1(G20), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(KEYINPUT23), .B2(new_n607), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(KEYINPUT24), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n611), .A2(new_n257), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n610), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT24), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n600), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n596), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT95), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n596), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT19), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n248), .A2(new_n250), .A3(G97), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n622), .A2(new_n623), .B1(new_n603), .B2(G68), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G87), .A2(G97), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n377), .ZN(new_n626));
  NAND3_X1  g0426(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n627), .A2(new_n628), .A3(new_n211), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n628), .B1(new_n627), .B2(new_n211), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n405), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n388), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n339), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT88), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n623), .A2(new_n622), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n603), .A2(G68), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n257), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  INV_X1    g0440(.A(new_n634), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n519), .A2(new_n633), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(G250), .B1(new_n484), .B2(G1), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n485), .A2(G274), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n272), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n351), .A2(G244), .A3(G1698), .ZN(new_n649));
  INV_X1    g0449(.A(G238), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(new_n608), .C1(new_n353), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n651), .B2(new_n272), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(new_n358), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(G179), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n325), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(G200), .B2(new_n652), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n519), .A2(G87), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n643), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n594), .A2(G169), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n594), .A2(new_n318), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n616), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n545), .A2(new_n584), .A3(new_n621), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n475), .A2(new_n666), .ZN(G372));
  INV_X1    g0467(.A(new_n475), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n643), .A2(new_n644), .B1(new_n653), .B2(new_n654), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n640), .B1(new_n639), .B2(new_n641), .ZN(new_n670));
  AOI211_X1 g0470(.A(KEYINPUT88), .B(new_n634), .C1(new_n638), .C2(new_n257), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n659), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT96), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n643), .A2(KEYINPUT96), .A3(new_n659), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n669), .B1(new_n676), .B2(new_n658), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n542), .A2(new_n543), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n521), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT21), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n530), .A2(G169), .A3(new_n531), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n680), .B1(new_n681), .B2(new_n541), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n663), .A2(new_n662), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n612), .A2(new_n615), .ZN(new_n684));
  INV_X1    g0484(.A(new_n600), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n679), .A2(new_n682), .A3(new_n687), .ZN(new_n688));
  AND4_X1   g0488(.A1(new_n584), .A2(new_n677), .A3(new_n688), .A4(new_n621), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n575), .A2(new_n656), .A3(new_n660), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n669), .B1(new_n690), .B2(KEYINPUT26), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n574), .A2(KEYINPUT97), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT97), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n569), .A2(new_n573), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT26), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT96), .B1(new_n643), .B2(new_n659), .ZN(new_n697));
  INV_X1    g0497(.A(new_n659), .ZN(new_n698));
  AOI211_X1 g0498(.A(new_n673), .B(new_n698), .C1(new_n635), .C2(new_n642), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n658), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(new_n700), .A4(new_n656), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n691), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n668), .B1(new_n689), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n361), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n459), .A2(new_n469), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n380), .A2(new_n318), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n394), .B1(new_n706), .B2(new_n397), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n310), .A2(G169), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT14), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n312), .A3(new_n320), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n330), .A2(new_n707), .B1(new_n710), .B2(new_n268), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n463), .A2(new_n472), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n705), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n704), .B1(new_n714), .B2(new_n373), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n703), .A2(new_n715), .ZN(G369));
  OR3_X1    g0516(.A1(new_n262), .A2(KEYINPUT27), .A3(G20), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT27), .B1(new_n262), .B2(G20), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G213), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G343), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n664), .A2(new_n721), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n618), .A2(new_n620), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n723), .B1(new_n686), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n722), .B1(new_n725), .B2(new_n664), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n679), .A2(new_n682), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n521), .ZN(new_n728));
  MUX2_X1   g0528(.A(new_n727), .B(new_n545), .S(new_n728), .Z(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n725), .A2(new_n727), .A3(new_n687), .A4(new_n721), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(new_n722), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n223), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n625), .A2(new_n377), .A3(new_n507), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n208), .B2(new_n738), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g0543(.A(new_n583), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n574), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n723), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n545), .A3(new_n665), .A4(new_n721), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT30), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n554), .A2(new_n652), .A3(new_n557), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n585), .B1(new_n591), .B2(new_n593), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n750), .A2(new_n543), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n752), .B2(KEYINPUT99), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT99), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n543), .A2(new_n751), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n754), .B(KEYINPUT30), .C1(new_n755), .C2(new_n750), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n576), .A2(new_n572), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n652), .A2(G179), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n530), .A2(new_n594), .A3(new_n531), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n721), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT31), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT100), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(new_n764), .B2(KEYINPUT31), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT31), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n762), .B1(new_n753), .B2(new_n756), .ZN(new_n769));
  OAI211_X1 g0569(.A(KEYINPUT100), .B(new_n768), .C1(new_n769), .C2(new_n721), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n748), .A2(new_n765), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  AND2_X1   g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n688), .A2(new_n677), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT103), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n746), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n584), .A2(KEYINPUT103), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n773), .A2(new_n775), .A3(new_n621), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n696), .B1(new_n677), .B2(new_n695), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n656), .B1(new_n690), .B2(KEYINPUT26), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT102), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n700), .A2(new_n656), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n692), .A2(new_n694), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT26), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n661), .A2(new_n574), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n669), .B1(new_n784), .B2(new_n696), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT102), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n777), .A2(new_n780), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(KEYINPUT29), .A3(new_n721), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n721), .B1(new_n689), .B2(new_n702), .ZN(new_n790));
  NOR2_X1   g0590(.A1(KEYINPUT101), .A2(KEYINPUT29), .ZN(new_n791));
  AND2_X1   g0591(.A1(KEYINPUT101), .A2(KEYINPUT29), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n772), .B1(new_n789), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n743), .B1(new_n794), .B2(G1), .ZN(G364));
  NOR2_X1   g0595(.A1(new_n260), .A2(G20), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G45), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n738), .A2(G1), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n730), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n729), .A2(G330), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n729), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n798), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n211), .A2(G190), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n808), .A2(G179), .A3(new_n364), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n211), .A2(new_n325), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n318), .A2(G200), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n809), .A2(G283), .B1(new_n813), .B2(G322), .ZN(new_n814));
  INV_X1    g0614(.A(G326), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n318), .A2(new_n364), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n810), .A2(new_n318), .A3(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n811), .A2(new_n807), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n820), .A2(G303), .B1(new_n822), .B2(G311), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n816), .A2(new_n807), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n351), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G294), .ZN(new_n828));
  NOR2_X1   g0628(.A1(G179), .A2(G200), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G190), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(G20), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n823), .B(new_n827), .C1(new_n828), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n807), .A2(new_n829), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT106), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(KEYINPUT106), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n818), .B(new_n833), .C1(G329), .C2(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n812), .A2(new_n202), .B1(new_n821), .B2(new_n252), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n841), .A2(KEYINPUT104), .B1(new_n201), .B2(new_n817), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(KEYINPUT104), .B2(new_n841), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT105), .Z(new_n844));
  NOR2_X1   g0644(.A1(new_n834), .A2(new_n417), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT32), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n831), .A2(G97), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n819), .A2(new_n440), .ZN(new_n849));
  INV_X1    g0649(.A(new_n809), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n850), .A2(new_n377), .B1(new_n203), .B2(new_n824), .ZN(new_n851));
  NOR4_X1   g0651(.A1(new_n848), .A2(new_n408), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n840), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n210), .B1(G20), .B2(new_n358), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n351), .A2(new_n223), .ZN(new_n856));
  INV_X1    g0656(.A(G355), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n856), .A2(new_n857), .B1(G116), .B2(new_n223), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n208), .A2(new_n484), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n240), .B2(new_n484), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n736), .A2(new_n351), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n803), .A2(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n806), .B1(new_n853), .B2(new_n855), .C1(new_n862), .C2(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n799), .A2(new_n800), .B1(new_n805), .B2(new_n865), .ZN(G396));
  OAI211_X1 g0666(.A(new_n395), .B(new_n400), .C1(new_n394), .C2(new_n721), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n707), .A2(KEYINPUT107), .A3(new_n724), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT107), .B1(new_n707), .B2(new_n724), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n790), .B(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n772), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n806), .B1(new_n772), .B2(new_n871), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n839), .A2(G311), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n850), .A2(new_n440), .ZN(new_n876));
  OAI22_X1  g0676(.A1(new_n819), .A2(new_n377), .B1(new_n821), .B2(new_n507), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n876), .A2(new_n351), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(G303), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n817), .A2(new_n879), .B1(new_n824), .B2(new_n504), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(G294), .B2(new_n813), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n875), .A2(new_n878), .A3(new_n847), .A4(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n817), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(G137), .B1(new_n822), .B2(G159), .ZN(new_n884));
  INV_X1    g0684(.A(G143), .ZN(new_n885));
  INV_X1    g0685(.A(G150), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n884), .B1(new_n885), .B2(new_n812), .C1(new_n886), .C2(new_n824), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT34), .Z(new_n888));
  OAI21_X1  g0688(.A(new_n351), .B1(new_n819), .B2(new_n201), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(G68), .B2(new_n809), .ZN(new_n890));
  INV_X1    g0690(.A(G132), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n890), .B1(new_n202), .B2(new_n832), .C1(new_n891), .C2(new_n838), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n882), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n854), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n854), .A2(new_n801), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n798), .B1(new_n252), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n870), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n801), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n874), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(G384));
  NOR2_X1   g0701(.A1(new_n796), .A2(new_n265), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n268), .A2(new_n724), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n331), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n323), .A2(new_n330), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n768), .B1(new_n769), .B2(new_n721), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n765), .B(new_n908), .C1(new_n666), .C2(new_n724), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n907), .A2(new_n870), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n720), .B1(new_n431), .B2(new_n436), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n912), .B(new_n470), .C1(new_n437), .C2(new_n458), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT111), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n913), .B(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n473), .A2(new_n467), .A3(new_n720), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n434), .A2(new_n404), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n720), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n473), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n470), .A2(new_n921), .ZN(new_n924));
  AND4_X1   g0724(.A1(new_n455), .A2(new_n920), .A3(new_n448), .A4(new_n457), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n464), .A2(new_n467), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n927), .A2(new_n914), .A3(new_n470), .A4(new_n912), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g0729(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n919), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT40), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n923), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n923), .A2(new_n929), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n923), .A2(KEYINPUT110), .A3(new_n929), .A4(KEYINPUT38), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n933), .B1(new_n942), .B2(new_n910), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n932), .A2(new_n943), .A3(G330), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n332), .A2(new_n474), .A3(new_n909), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(G330), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n932), .A2(new_n943), .A3(new_n945), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n936), .A2(new_n939), .A3(KEYINPUT39), .A4(new_n940), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n919), .B2(new_n930), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n710), .A2(new_n268), .A3(new_n721), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n705), .A2(new_n720), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n870), .B(new_n721), .C1(new_n689), .C2(new_n702), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT109), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n707), .A2(new_n721), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT108), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n961), .B1(new_n960), .B2(new_n963), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n941), .B(new_n907), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n959), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n789), .A2(new_n668), .A3(new_n793), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n715), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n902), .B1(new_n951), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n951), .B2(new_n970), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n209), .A2(G77), .A3(new_n413), .A4(new_n414), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(G50), .B2(new_n203), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n974), .A2(G1), .A3(new_n260), .ZN(new_n975));
  INV_X1    g0775(.A(new_n563), .ZN(new_n976));
  OAI211_X1 g0776(.A(G116), .B(new_n212), .C1(new_n976), .C2(KEYINPUT35), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n977), .B1(KEYINPUT35), .B2(new_n976), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT36), .Z(new_n979));
  NAND3_X1  g0779(.A1(new_n972), .A2(new_n975), .A3(new_n979), .ZN(G367));
  XOR2_X1   g0780(.A(new_n737), .B(KEYINPUT41), .Z(new_n981));
  NAND2_X1  g0781(.A1(new_n566), .A2(new_n568), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n724), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n775), .A2(new_n776), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n575), .A2(new_n724), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT45), .B1(new_n734), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n733), .A2(new_n722), .ZN(new_n988));
  INV_X1    g0788(.A(new_n986), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT45), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT44), .B1(new_n734), .B2(new_n986), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT44), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n988), .A2(new_n994), .A3(new_n989), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n996), .A3(new_n732), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n987), .A2(new_n991), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n993), .A2(new_n995), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n731), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n727), .A2(new_n721), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n726), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n733), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(new_n730), .Z(new_n1004));
  NAND4_X1  g0804(.A1(new_n997), .A2(new_n1000), .A3(new_n794), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n981), .B1(new_n1005), .B2(new_n794), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n797), .A2(G1), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT113), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n989), .A2(new_n733), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT42), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n984), .A2(new_n687), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n724), .B1(new_n1014), .B2(new_n574), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n676), .A2(new_n721), .ZN(new_n1018));
  MUX2_X1   g0818(.A(new_n781), .B(new_n656), .S(new_n1018), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1016), .A2(new_n1017), .B1(KEYINPUT43), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n731), .A2(new_n986), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1021), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1010), .A2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n235), .A2(new_n736), .A3(new_n351), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n864), .B1(new_n736), .B2(new_n633), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n798), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n809), .A2(G77), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1031), .B1(new_n1032), .B2(new_n834), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n408), .B(new_n1033), .C1(G58), .C2(new_n820), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G159), .A2(new_n825), .B1(new_n822), .B2(G50), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G143), .A2(new_n883), .B1(new_n813), .B2(G150), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n831), .A2(G68), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n408), .B1(new_n834), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n828), .A2(new_n824), .B1(new_n812), .B2(new_n879), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G107), .C2(new_n831), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n820), .A2(G116), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT46), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n809), .A2(G97), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n883), .A2(G311), .B1(new_n822), .B2(G283), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT47), .B1(new_n1038), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1038), .A2(KEYINPUT47), .A3(new_n1047), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n854), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1030), .B1(new_n1048), .B2(new_n1050), .C1(new_n1020), .C2(new_n804), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1026), .A2(new_n1051), .ZN(G387));
  NAND2_X1  g0852(.A1(new_n232), .A2(G45), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n383), .A2(new_n201), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n740), .B(new_n484), .C1(new_n203), .C2(new_n252), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1053), .B(new_n861), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n856), .A2(new_n740), .B1(G107), .B2(new_n223), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n798), .B1(new_n1060), .B2(new_n863), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT115), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G50), .A2(new_n813), .B1(new_n835), .B2(G150), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n351), .A3(new_n1045), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n824), .A2(new_n335), .B1(new_n821), .B2(new_n203), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n819), .A2(new_n252), .B1(new_n817), .B2(new_n417), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n832), .A2(new_n388), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G311), .A2(new_n825), .B1(new_n813), .B2(G317), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n883), .A2(G322), .B1(new_n822), .B2(G303), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT48), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT48), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n820), .A2(G294), .B1(G283), .B2(new_n831), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n408), .B1(new_n815), .B2(new_n834), .C1(new_n850), .C2(new_n507), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1068), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1062), .B1(new_n855), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n726), .B2(new_n803), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1004), .A2(new_n794), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n737), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1004), .A2(new_n794), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n997), .A2(new_n1000), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n737), .A3(new_n1005), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n997), .A2(new_n1000), .A3(new_n1008), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(G317), .A2(new_n883), .B1(new_n813), .B2(G311), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT52), .Z(new_n1094));
  OAI21_X1  g0894(.A(new_n408), .B1(new_n850), .B2(new_n377), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G116), .B2(new_n831), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n825), .A2(G303), .B1(new_n835), .B2(G322), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n820), .A2(G283), .B1(new_n822), .B2(G294), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT118), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n824), .A2(new_n201), .B1(new_n821), .B2(new_n335), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT117), .Z(new_n1102));
  OAI22_X1  g0902(.A1(new_n819), .A2(new_n203), .B1(new_n834), .B2(new_n885), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n876), .A2(new_n408), .A3(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n817), .A2(new_n886), .B1(new_n812), .B2(new_n417), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n832), .A2(new_n252), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n855), .B1(new_n1100), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n863), .B1(new_n560), .B2(new_n223), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n243), .B2(new_n861), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1110), .A2(new_n798), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n986), .B2(new_n804), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1091), .A2(new_n1092), .A3(new_n1114), .ZN(G390));
  NAND2_X1  g0915(.A1(new_n952), .A2(new_n954), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n801), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n798), .B1(new_n335), .B2(new_n895), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n351), .B1(new_n201), .B2(new_n850), .C1(new_n838), .C2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT119), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G132), .A2(new_n813), .B1(new_n825), .B2(G137), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n820), .A2(G150), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT53), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1123), .A2(KEYINPUT53), .B1(new_n831), .B2(G159), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n883), .A2(G128), .B1(new_n822), .B2(new_n1127), .ZN(new_n1128));
  AND4_X1   g0928(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .A4(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n850), .A2(new_n203), .B1(new_n504), .B2(new_n817), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1130), .A2(new_n351), .A3(new_n849), .A4(new_n1107), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G107), .A2(new_n825), .B1(new_n822), .B2(G97), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n507), .B2(new_n812), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G294), .B2(new_n839), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1121), .A2(new_n1129), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n854), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1117), .B(new_n1118), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n323), .A2(new_n330), .A3(new_n903), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n903), .B1(new_n323), .B2(new_n330), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n960), .A2(new_n963), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT109), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1116), .B1(new_n1146), .B2(new_n956), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n788), .A2(new_n721), .A3(new_n870), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n963), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n907), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1150), .A2(new_n931), .A3(new_n955), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n870), .A2(G330), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n909), .B(new_n1153), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n907), .A2(new_n771), .A3(G330), .A4(new_n870), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1147), .A2(new_n1151), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1008), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1139), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n909), .A2(new_n1153), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n906), .A3(new_n905), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1163), .A2(new_n963), .A3(new_n1148), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n765), .B1(new_n666), .B2(new_n724), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n767), .A2(new_n770), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G330), .B(new_n870), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n1142), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1154), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1164), .A2(new_n1157), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n968), .A2(new_n946), .A3(new_n715), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1156), .A2(new_n1158), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1173), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n738), .B1(new_n1159), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1161), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(G378));
  INV_X1    g0978(.A(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1174), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n932), .A2(new_n943), .A3(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n373), .A2(new_n360), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n342), .A2(new_n720), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1183), .B(new_n1184), .ZN(new_n1185));
  XOR2_X1   g0985(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n959), .B2(new_n966), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n966), .A2(new_n958), .A3(new_n957), .A4(new_n1187), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1182), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1187), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n966), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n957), .A2(new_n958), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1195), .A2(new_n944), .A3(new_n1189), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1180), .A2(new_n1181), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1181), .B1(new_n1180), .B2(new_n1197), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n737), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1187), .A2(new_n801), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n895), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n806), .B1(G50), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n351), .A2(G41), .ZN(new_n1204));
  INV_X1    g1004(.A(G41), .ZN(new_n1205));
  AOI211_X1 g1005(.A(G50), .B(new_n1204), .C1(new_n246), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n839), .A2(G283), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G58), .A2(new_n809), .B1(new_n820), .B2(G77), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n883), .A2(G116), .B1(new_n822), .B2(new_n633), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1208), .A2(new_n1037), .A3(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G97), .A2(new_n825), .B1(new_n813), .B2(G107), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1207), .A2(new_n1210), .A3(new_n1204), .A4(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1206), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n824), .A2(new_n891), .B1(new_n821), .B2(new_n1032), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT121), .Z(new_n1216));
  NOR2_X1   g1016(.A1(new_n832), .A2(new_n886), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n819), .A2(new_n1126), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n817), .A2(new_n1119), .B1(new_n812), .B2(new_n1219), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n246), .B(new_n1205), .C1(new_n850), .C2(new_n417), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G124), .B2(new_n835), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1214), .B1(new_n1213), .B2(new_n1212), .C1(new_n1223), .C2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1203), .B1(new_n1228), .B2(new_n854), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1201), .A2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT122), .Z(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1197), .B2(new_n1008), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1200), .A2(new_n1232), .ZN(G375));
  INV_X1    g1033(.A(new_n981), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1157), .A2(new_n963), .A3(new_n1148), .A4(new_n1163), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1172), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1175), .A2(new_n1234), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1142), .A2(new_n801), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n806), .B1(G68), .B2(new_n1202), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G132), .A2(new_n883), .B1(new_n813), .B2(G137), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n408), .B1(new_n809), .B2(G58), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(new_n201), .C2(new_n832), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n820), .A2(G159), .B1(new_n825), .B2(new_n1127), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n886), .B2(new_n821), .C1(new_n838), .C2(new_n1219), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n820), .A2(G97), .B1(new_n822), .B2(G107), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n828), .B2(new_n817), .C1(new_n838), .C2(new_n879), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1067), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G116), .A2(new_n825), .B1(new_n813), .B2(G283), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n408), .A4(new_n1031), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1244), .A2(new_n1246), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1241), .B1(new_n1252), .B2(new_n854), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1239), .A2(new_n1008), .B1(new_n1240), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1238), .A2(new_n1254), .ZN(G381));
  NOR2_X1   g1055(.A1(G375), .A2(G378), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1025), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1051), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(G390), .A3(new_n1259), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1256), .A2(new_n1260), .A3(new_n1261), .ZN(G407));
  INV_X1    g1062(.A(G213), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1263), .A2(G343), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1256), .A2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G407), .A2(G213), .A3(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1067(.A(new_n1264), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n737), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1237), .A2(KEYINPUT60), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1171), .A2(new_n1271), .A3(new_n1172), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1269), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1254), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n900), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n738), .B1(new_n1239), .B2(new_n1179), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1271), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1277));
  AND4_X1   g1077(.A1(new_n1271), .A2(new_n1172), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(G384), .A3(new_n1254), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1180), .A2(new_n1234), .A3(new_n1197), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1230), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1195), .A2(new_n944), .A3(new_n1189), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n944), .B1(new_n1195), .B2(new_n1189), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT124), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1191), .A2(new_n1289), .A3(new_n1196), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1285), .B1(new_n1291), .B2(new_n1008), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1284), .B1(new_n1292), .B2(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT125), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1160), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1295), .B2(new_n1285), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G378), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1200), .A2(G378), .A3(new_n1232), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1268), .B(new_n1282), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT62), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1268), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT126), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1302), .B1(new_n1275), .B2(new_n1280), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1264), .A2(G2897), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1282), .A2(new_n1302), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1279), .A2(G384), .A3(new_n1254), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G384), .B1(new_n1279), .B2(new_n1254), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT126), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1304), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1306), .A2(new_n1307), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1307), .B1(new_n1306), .B2(new_n1312), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1301), .A2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT61), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1286), .A2(new_n1287), .A3(KEYINPUT124), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1289), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1008), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(KEYINPUT125), .A3(new_n1230), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1296), .A2(new_n1321), .A3(new_n1283), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1177), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1200), .A2(G378), .A3(new_n1232), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1325), .A2(new_n1326), .A3(new_n1268), .A4(new_n1282), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1300), .A2(new_n1316), .A3(new_n1317), .A4(new_n1327), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(G393), .B(G396), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(G390), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1331), .B1(new_n1026), .B2(new_n1051), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1332), .B2(new_n1260), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1026), .A2(new_n1051), .A3(new_n1331), .ZN(new_n1334));
  OAI21_X1  g1134(.A(G390), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1329), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1328), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1264), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1307), .ZN(new_n1340));
  NOR3_X1   g1140(.A1(new_n1303), .A2(KEYINPUT127), .A3(new_n1305), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1311), .B1(new_n1310), .B2(new_n1304), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1306), .A2(new_n1312), .A3(new_n1307), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT63), .B1(new_n1339), .B2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1299), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1333), .A2(new_n1317), .A3(new_n1336), .ZN(new_n1348));
  AOI211_X1 g1148(.A(new_n1264), .B(new_n1281), .C1(new_n1323), .C2(new_n1324), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1349), .B2(KEYINPUT63), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1347), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1338), .A2(new_n1351), .ZN(G405));
  NAND2_X1  g1152(.A1(new_n1337), .A2(new_n1281), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1333), .A2(new_n1336), .A3(new_n1282), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1177), .B1(new_n1200), .B2(new_n1232), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1355), .B1(new_n1256), .B2(new_n1356), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1256), .A2(new_n1356), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1353), .A2(new_n1358), .A3(new_n1354), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1357), .A2(new_n1359), .ZN(G402));
endmodule


