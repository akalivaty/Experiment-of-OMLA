//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n542, new_n543, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G219), .A3(G220), .A4(G218), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(new_n466), .ZN(G160));
  OR2_X1    g042(.A1(G100), .A2(G2105), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n468), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n460), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n477), .A3(new_n459), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n477), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(G124), .B2(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n484), .A2(KEYINPUT4), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n485), .A2(new_n471), .A3(new_n473), .A4(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(G102), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n459), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n471), .A2(new_n473), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n459), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT69), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT69), .A2(G651), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT6), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G651), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n498), .A2(G50), .A3(G543), .A4(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n496), .A2(new_n497), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G88), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n507));
  OAI221_X1 g082(.A(new_n501), .B1(new_n503), .B2(new_n505), .C1(new_n506), .C2(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  NAND2_X1  g084(.A1(new_n498), .A2(new_n500), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G51), .ZN(new_n513));
  INV_X1    g088(.A(new_n507), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n502), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n513), .A2(new_n515), .A3(new_n516), .A4(new_n518), .ZN(G286));
  INV_X1    g094(.A(G286), .ZN(G168));
  AOI22_X1  g095(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n505), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n498), .A2(G52), .A3(G543), .A4(new_n500), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n498), .A2(G90), .A3(new_n500), .A4(new_n502), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n525), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n530), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G171));
  NAND2_X1  g107(.A1(new_n512), .A2(G43), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n514), .A2(G81), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n505), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  NAND4_X1  g119(.A1(new_n498), .A2(G53), .A3(G543), .A4(new_n500), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n502), .A2(G65), .ZN(new_n547));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT72), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n514), .A2(G91), .B1(new_n550), .B2(G651), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(G299));
  INV_X1    g127(.A(G171), .ZN(G301));
  NAND2_X1  g128(.A1(new_n512), .A2(G49), .ZN(new_n554));
  OAI21_X1  g129(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g132(.A(KEYINPUT73), .B(G651), .C1(new_n502), .C2(G74), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n514), .A2(G87), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(G288));
  NAND4_X1  g136(.A1(new_n498), .A2(G86), .A3(new_n500), .A4(new_n502), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n498), .A2(G48), .A3(G543), .A4(new_n500), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n502), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n505), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT5), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n568), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n574), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n564), .A2(new_n567), .A3(new_n575), .ZN(G305));
  NAND2_X1  g151(.A1(new_n512), .A2(G47), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n514), .A2(G85), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n505), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(G290));
  INV_X1    g156(.A(G92), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n507), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G54), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G651), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n507), .B2(new_n582), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n583), .A2(new_n584), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G171), .B2(new_n590), .ZN(G284));
  OAI21_X1  g167(.A(new_n591), .B1(G171), .B2(new_n590), .ZN(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G299), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(new_n589), .ZN(new_n598));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n537), .A2(new_n590), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n589), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n590), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n482), .A2(G123), .ZN(new_n605));
  INV_X1    g180(.A(new_n478), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G135), .ZN(new_n607));
  OAI21_X1  g182(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n611), .A2(new_n459), .A3(G111), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n459), .B2(G111), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n609), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n610), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n605), .A2(new_n607), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2072), .B(G2078), .Z(new_n638));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n642), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2100), .Z(new_n645));
  AND2_X1   g220(.A1(new_n642), .A2(KEYINPUT17), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  AOI21_X1  g222(.A(KEYINPUT18), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(G227));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT78), .ZN(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n651), .A2(new_n652), .ZN(new_n658));
  AOI22_X1  g233(.A1(new_n656), .A2(new_n657), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n653), .A2(new_n658), .A3(new_n655), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n660), .C1(new_n657), .C2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G1986), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT82), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT79), .B(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(G25), .A2(G29), .ZN(new_n678));
  OR2_X1    g253(.A1(G95), .A2(G2105), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n679), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n680));
  INV_X1    g255(.A(G119), .ZN(new_n681));
  INV_X1    g256(.A(G131), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n680), .B1(new_n481), .B2(new_n681), .C1(new_n682), .C2(new_n478), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n678), .B1(new_n685), .B2(G29), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT35), .B(G1991), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT84), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n686), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  NAND2_X1  g266(.A1(G303), .A2(G16), .ZN(new_n692));
  INV_X1    g267(.A(G22), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G16), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n691), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g271(.A(G1971), .B(new_n694), .C1(G303), .C2(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n554), .A2(new_n559), .A3(new_n560), .A4(G16), .ZN(new_n699));
  OR2_X1    g274(.A1(G16), .A2(G23), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT33), .B(G1976), .Z(new_n701));
  AND3_X1   g276(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n699), .B2(new_n700), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n705), .A2(G6), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G305), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT85), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n707), .A2(new_n709), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n698), .A2(new_n704), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n712), .A2(KEYINPUT86), .A3(KEYINPUT34), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT86), .B1(new_n712), .B2(KEYINPUT34), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n690), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(G16), .A2(G24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G290), .B2(new_n705), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(G1986), .Z(new_n720));
  OAI211_X1 g295(.A(new_n675), .B(new_n677), .C1(new_n717), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n716), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n712), .A2(KEYINPUT86), .A3(KEYINPUT34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n713), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n720), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n724), .A2(new_n725), .A3(new_n690), .A4(new_n676), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n538), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT89), .B(G1341), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n705), .A2(KEYINPUT23), .A3(G20), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n732));
  INV_X1    g307(.A(G20), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n731), .B(new_n734), .C1(new_n595), .C2(new_n705), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1956), .ZN(new_n736));
  NOR2_X1   g311(.A1(G29), .A2(G35), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G162), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT29), .B(G2090), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n721), .A2(new_n726), .A3(new_n730), .A4(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n743));
  INV_X1    g318(.A(G1961), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n705), .B1(new_n529), .B2(new_n531), .ZN(new_n745));
  NOR2_X1   g320(.A1(G5), .A2(G16), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n745), .A2(KEYINPUT93), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(KEYINPUT93), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(G16), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G286), .B2(new_n705), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT92), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n752), .A2(new_n756), .A3(new_n753), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n616), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT91), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(G1966), .B(new_n751), .C1(G286), .C2(new_n705), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT30), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G28), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n759), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n758), .A2(new_n761), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n743), .B1(new_n750), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n770), .ZN(new_n772));
  INV_X1    g347(.A(new_n749), .ZN(new_n773));
  OAI21_X1  g348(.A(G1961), .B1(new_n773), .B2(new_n747), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n772), .A2(KEYINPUT94), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n748), .A2(new_n744), .A3(new_n749), .ZN(new_n777));
  OR2_X1    g352(.A1(G29), .A2(G33), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT25), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  INV_X1    g356(.A(G139), .ZN(new_n782));
  OAI221_X1 g357(.A(new_n780), .B1(new_n459), .B2(new_n781), .C1(new_n478), .C2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n783), .B2(new_n759), .ZN(new_n784));
  INV_X1    g359(.A(G2072), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT90), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT90), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G32), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G129), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n606), .A2(G141), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT26), .Z(new_n796));
  NAND4_X1  g371(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n791), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(G27), .A2(G29), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G164), .B2(G29), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n777), .A2(new_n790), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(KEYINPUT24), .A2(G34), .ZN(new_n807));
  NAND2_X1  g382(.A1(KEYINPUT24), .A2(G34), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n807), .A2(new_n759), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G160), .B2(new_n759), .ZN(new_n810));
  INV_X1    g385(.A(G2084), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n776), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT95), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n776), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n742), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT96), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n759), .A2(G26), .ZN(new_n821));
  OR2_X1    g396(.A1(G104), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n823));
  INV_X1    g398(.A(G128), .ZN(new_n824));
  INV_X1    g399(.A(G140), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n823), .B1(new_n481), .B2(new_n824), .C1(new_n825), .C2(new_n478), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n821), .B1(new_n826), .B2(G29), .ZN(new_n827));
  MUX2_X1   g402(.A(new_n821), .B(new_n827), .S(KEYINPUT28), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2067), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n705), .A2(G4), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n598), .B2(new_n705), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT88), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1348), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n819), .A2(new_n820), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  AND4_X1   g409(.A1(new_n730), .A2(new_n721), .A3(new_n726), .A4(new_n741), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n816), .A2(new_n818), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n829), .A4(new_n833), .ZN(G150));
  NAND2_X1  g412(.A1(G150), .A2(KEYINPUT96), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(G311));
  AOI22_X1  g414(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n505), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n512), .A2(G55), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n845), .B2(new_n507), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n847), .B(new_n537), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n598), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n850), .B1(new_n855), .B2(G860), .ZN(G145));
  XNOR2_X1  g431(.A(new_n616), .B(G160), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(G162), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n797), .B(new_n683), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n783), .B(new_n619), .ZN(new_n861));
  XNOR2_X1  g436(.A(G164), .B(KEYINPUT98), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n606), .A2(G142), .ZN(new_n864));
  OAI21_X1  g439(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n459), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G130), .B2(new_n482), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n826), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n863), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n860), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g449(.A(new_n847), .B(new_n538), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n602), .ZN(new_n876));
  XOR2_X1   g451(.A(G299), .B(new_n589), .Z(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n876), .B(new_n880), .C1(KEYINPUT41), .C2(new_n878), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n877), .B(KEYINPUT99), .Z(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n884), .A2(KEYINPUT101), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(G303), .ZN(new_n887));
  INV_X1    g462(.A(G288), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G305), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(G305), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(KEYINPUT101), .B2(new_n884), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n883), .A2(new_n885), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n886), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n896), .B1(new_n886), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n848), .A2(new_n590), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n901), .ZN(G331));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n895), .B(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G171), .B(G168), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n875), .ZN(new_n908));
  XNOR2_X1  g483(.A(G171), .B(G286), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n851), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n880), .B1(KEYINPUT41), .B2(new_n878), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(KEYINPUT102), .A3(new_n875), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n908), .A2(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n877), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n915), .A2(new_n917), .A3(new_n893), .A4(new_n894), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n872), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n904), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n912), .A2(new_n914), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n923), .A2(new_n882), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n878), .A2(new_n879), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT104), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n916), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n906), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n929), .A2(KEYINPUT43), .A3(new_n872), .A4(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT44), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n919), .B2(new_n921), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(new_n904), .A3(new_n872), .A4(new_n920), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n937), .ZN(G397));
  OAI21_X1  g513(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n939));
  INV_X1    g514(.A(G40), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n463), .A2(new_n466), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n484), .A2(KEYINPUT4), .A3(G138), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n487), .B1(new_n474), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n459), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n492), .A2(new_n493), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G2105), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n489), .A2(new_n490), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n939), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G1956), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n463), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n464), .A2(new_n465), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n459), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n957), .A3(G40), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n948), .A2(new_n950), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT107), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n948), .A2(new_n964), .A3(KEYINPUT45), .A4(new_n950), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT56), .B(G2072), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n961), .A2(new_n963), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n954), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G299), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n546), .A2(new_n551), .A3(new_n969), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT9), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n545), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n550), .A2(G651), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n498), .A2(G91), .A3(new_n500), .A4(new_n502), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n976), .A2(new_n979), .A3(new_n970), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n969), .B1(new_n546), .B2(new_n551), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT117), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n968), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n968), .A2(new_n983), .A3(KEYINPUT118), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1348), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n952), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n941), .A2(new_n950), .A3(new_n948), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n991), .A2(KEYINPUT116), .A3(G2067), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT116), .B1(new_n991), .B2(G2067), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n988), .B1(new_n589), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n971), .A2(new_n972), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n954), .A2(new_n967), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n968), .A2(KEYINPUT118), .A3(new_n983), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT118), .B1(new_n968), .B2(new_n983), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT61), .B(new_n997), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n988), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n997), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n968), .B(new_n996), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(KEYINPUT61), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n589), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n598), .A2(KEYINPUT122), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n994), .A2(KEYINPUT60), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n990), .A2(new_n992), .A3(new_n993), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1007), .B(new_n589), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1010), .B(new_n1013), .C1(KEYINPUT60), .C2(new_n994), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT58), .B(G1341), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n991), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(G1996), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT119), .B(new_n1017), .C1(new_n1018), .C2(G1996), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n538), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1021), .A2(KEYINPUT120), .A3(new_n538), .A4(new_n1022), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(KEYINPUT59), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1023), .A2(new_n1024), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n998), .B1(new_n1015), .B2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n554), .A2(new_n559), .A3(new_n560), .A4(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n991), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1033), .B(new_n1035), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n888), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n991), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G305), .A2(new_n1039), .A3(G1981), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT111), .B(G1981), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(G305), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n567), .A2(new_n575), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(new_n564), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1040), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1038), .B1(new_n1046), .B2(KEYINPUT49), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1040), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1036), .A2(new_n1037), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(KEYINPUT113), .B2(G8), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT109), .B(G2090), .Z(new_n1055));
  INV_X1    g630(.A(new_n952), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT108), .B(G1971), .Z(new_n1057));
  AOI22_X1  g632(.A1(new_n1055), .A2(new_n1056), .B1(new_n1018), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1054), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1051), .B(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1059), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1056), .A2(new_n1055), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1018), .A2(new_n1057), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1050), .A2(new_n1060), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n952), .A2(new_n744), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n961), .A2(KEYINPUT53), .A3(new_n804), .A4(new_n962), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT123), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n961), .A2(new_n963), .A3(new_n804), .A4(new_n965), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT124), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1075), .A2(new_n1079), .A3(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(G171), .B(KEYINPUT54), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n948), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT45), .B1(new_n948), .B2(new_n950), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n958), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT114), .B1(new_n1088), .B2(G1966), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1056), .A2(new_n811), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n961), .A2(new_n962), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n753), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .A4(G168), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT51), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(G286), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1095), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1067), .B(new_n1085), .C1(new_n1097), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1081), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1083), .B1(new_n1076), .B2(new_n1075), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1068), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT125), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1050), .A2(new_n1060), .A3(new_n1066), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n1100), .A2(new_n1095), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(new_n1096), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1106), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1085), .A4(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1031), .A2(new_n1107), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G286), .A2(new_n1059), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1099), .B(new_n1115), .C1(new_n1116), .C2(new_n1053), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1050), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT63), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G305), .A2(new_n1041), .ZN(new_n1120));
  AOI21_X1  g695(.A(G1976), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n888), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1038), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1116), .A2(new_n1053), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1066), .A2(new_n1060), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1099), .A2(new_n1126), .A3(new_n1115), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1128), .B2(new_n1050), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1096), .B(new_n1130), .C1(new_n1095), .C2(new_n1100), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1108), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1133), .A3(G171), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT126), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT62), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1131), .A2(new_n1133), .A3(new_n1137), .A4(G171), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1114), .A2(new_n1129), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1087), .A2(new_n941), .ZN(new_n1141));
  INV_X1    g716(.A(G1996), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n797), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1141), .B(KEYINPUT105), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n826), .B(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n1142), .B2(new_n798), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n683), .B(new_n687), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(G290), .A2(G1986), .ZN(new_n1153));
  NOR2_X1   g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1141), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT106), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1140), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1147), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1145), .B1(new_n797), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1143), .B(KEYINPUT46), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(new_n1162), .B(KEYINPUT47), .Z(new_n1163));
  INV_X1    g738(.A(new_n687), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1149), .A2(new_n1164), .A3(new_n685), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n826), .A2(G2067), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1145), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT127), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1141), .A2(new_n1154), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT48), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1163), .B(new_n1168), .C1(new_n1152), .C2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1158), .A2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g747(.A1(new_n873), .A2(new_n671), .ZN(new_n1174));
  INV_X1    g748(.A(G319), .ZN(new_n1175));
  NOR3_X1   g749(.A1(G401), .A2(new_n1175), .A3(G227), .ZN(new_n1176));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n1174), .A3(new_n1176), .ZN(G225));
  INV_X1    g751(.A(G225), .ZN(G308));
endmodule


