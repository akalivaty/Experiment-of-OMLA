//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(G211gat), .ZN(new_n205));
  INV_X1    g004(.A(G218gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n203), .A3(new_n207), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(KEYINPUT74), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G226gat), .ZN(new_n217));
  INV_X1    g016(.A(G233gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT26), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(KEYINPUT69), .B2(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n222), .A2(new_n223), .A3(new_n220), .A4(new_n221), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT67), .B(G190gat), .Z(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  OR3_X1    g031(.A1(new_n232), .A2(KEYINPUT68), .A3(KEYINPUT27), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT27), .B1(new_n232), .B2(KEYINPUT68), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n230), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(KEYINPUT27), .B(G183gat), .Z(new_n236));
  OR2_X1    g035(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT28), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n228), .A2(new_n229), .A3(new_n235), .A4(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NOR3_X1   g042(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n226), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n232), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n245), .A2(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n226), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n220), .A3(new_n221), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n242), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT25), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n226), .B(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n242), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n247), .B(KEYINPUT66), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n237), .A2(new_n232), .A3(new_n238), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n263), .A2(new_n250), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n241), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n219), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n219), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n229), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n250), .C1(G183gat), .C2(G190gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n255), .B2(KEYINPUT64), .ZN(new_n274));
  AOI211_X1 g073(.A(new_n246), .B(new_n252), .C1(new_n254), .C2(new_n242), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n270), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n262), .A2(new_n250), .A3(new_n263), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n259), .A2(KEYINPUT25), .A3(new_n260), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n269), .B1(new_n280), .B2(new_n241), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n216), .B1(new_n268), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n245), .A2(new_n246), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n256), .A3(new_n273), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n284), .A2(new_n270), .B1(new_n277), .B2(new_n278), .ZN(new_n285));
  INV_X1    g084(.A(new_n241), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n219), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n216), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT29), .B1(new_n280), .B2(new_n241), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(new_n219), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n282), .A2(KEYINPUT75), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n216), .C1(new_n268), .C2(new_n281), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  XOR2_X1   g094(.A(G8gat), .B(G36gat), .Z(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT76), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n297), .B(new_n298), .Z(new_n299));
  NAND4_X1  g098(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT30), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n240), .A2(new_n235), .A3(new_n229), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n276), .A2(new_n279), .B1(new_n302), .B2(new_n228), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n269), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n288), .B1(new_n304), .B2(new_n287), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n293), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT30), .B(new_n299), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n299), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n293), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(KEYINPUT77), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT30), .B1(new_n294), .B2(new_n299), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n300), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT84), .B(KEYINPUT0), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(KEYINPUT85), .ZN(new_n315));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G57gat), .B(G85gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  OR2_X1    g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT79), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT79), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n323), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n322), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT80), .B1(new_n322), .B2(KEYINPUT2), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT81), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G141gat), .B(G148gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n335), .B1(KEYINPUT79), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n322), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n337), .A2(new_n338), .A3(new_n343), .A4(new_n323), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n339), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n336), .A2(KEYINPUT78), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n320), .A2(new_n348), .A3(new_n322), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G120gat), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G113gat), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT1), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G127gat), .B(G134gat), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT70), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G134gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(G127gat), .ZN(new_n360));
  INV_X1    g159(.A(G127gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G134gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(KEYINPUT1), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n354), .A2(KEYINPUT71), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT71), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G120gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(G113gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n354), .B2(G113gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n352), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n363), .A2(KEYINPUT1), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n358), .A2(new_n366), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND4_X1   g175(.A1(KEYINPUT4), .A2(new_n345), .A3(new_n351), .A4(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n350), .B1(new_n334), .B2(new_n344), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT4), .B1(new_n378), .B2(new_n376), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT86), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n345), .A2(new_n351), .A3(new_n376), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n376), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n380), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n345), .A2(new_n351), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n358), .A2(new_n366), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n374), .A2(new_n375), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n392), .B2(new_n394), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n398));
  AND3_X1   g197(.A1(new_n323), .A2(new_n326), .A3(new_n329), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n338), .B1(new_n399), .B2(new_n343), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT81), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n398), .B(new_n351), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n391), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(new_n383), .A3(new_n385), .A4(new_n389), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT1), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n354), .A2(G113gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n352), .A2(G120gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n364), .B1(new_n409), .B2(new_n363), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n356), .A2(KEYINPUT70), .A3(new_n357), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n394), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n376), .A2(new_n393), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n381), .B1(new_n415), .B2(new_n378), .ZN(new_n416));
  INV_X1    g215(.A(new_n389), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n388), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n405), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n405), .B2(new_n418), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n319), .B(new_n404), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n395), .A2(new_n378), .A3(new_n396), .ZN(new_n425));
  INV_X1    g224(.A(new_n381), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n402), .A2(new_n413), .A3(new_n414), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n378), .A2(new_n398), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n389), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n383), .A2(new_n385), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n427), .B(KEYINPUT5), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT83), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n405), .A2(new_n418), .A3(new_n419), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n319), .B1(new_n435), .B2(new_n404), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n424), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n404), .B1(new_n420), .B2(new_n421), .ZN(new_n438));
  INV_X1    g237(.A(new_n319), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n313), .B1(new_n437), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n443));
  INV_X1    g242(.A(G22gat), .ZN(new_n444));
  INV_X1    g243(.A(G228gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n218), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n288), .B1(new_n402), .B2(new_n267), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n211), .A2(new_n213), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n449), .B2(new_n267), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n378), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT88), .B(new_n447), .C1(new_n448), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n398), .B1(new_n216), .B2(KEYINPUT29), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n390), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n446), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n448), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n444), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(G22gat), .B(new_n460), .C1(new_n454), .C2(new_n455), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n443), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(G78gat), .B(G106gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n455), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n378), .B2(new_n398), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n471), .A2(new_n288), .B1(new_n378), .B2(new_n450), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT88), .B1(new_n472), .B2(new_n447), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n461), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(G22gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n444), .A3(new_n461), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(new_n443), .A3(new_n467), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n376), .B1(new_n285), .B2(new_n286), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n280), .A2(new_n412), .A3(new_n241), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G227gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n218), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G43gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(G71gat), .B(G99gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n483), .A3(new_n480), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(KEYINPUT32), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n489), .A2(KEYINPUT73), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT73), .B1(new_n489), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n489), .B(KEYINPUT32), .C1(new_n491), .C2(new_n488), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n485), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n489), .A2(KEYINPUT32), .ZN(new_n500));
  INV_X1    g299(.A(new_n488), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n493), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n489), .A2(KEYINPUT73), .A3(new_n491), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n496), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT34), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n485), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n469), .A2(new_n478), .A3(new_n499), .A4(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n202), .B1(new_n442), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n438), .A2(new_n439), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n423), .A3(new_n422), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n294), .A2(new_n299), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n310), .A2(KEYINPUT77), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n308), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n514), .A2(new_n440), .B1(new_n519), .B2(new_n300), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n467), .B1(new_n477), .B2(new_n443), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT87), .B(new_n468), .C1(new_n475), .C2(new_n476), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n497), .A2(new_n498), .A3(new_n485), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n520), .A2(new_n523), .A3(new_n526), .A4(KEYINPUT35), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n309), .A2(KEYINPUT37), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n310), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n291), .A2(KEYINPUT37), .A3(new_n293), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT38), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n282), .A2(new_n290), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT38), .B1(new_n533), .B2(KEYINPUT37), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n529), .A2(new_n534), .B1(new_n294), .B2(new_n299), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n514), .A2(new_n440), .A3(new_n532), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n523), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n389), .B1(new_n387), .B2(new_n403), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n439), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n416), .A2(new_n417), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n539), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n428), .A2(new_n429), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n380), .B2(new_n386), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n544), .B2(new_n389), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(KEYINPUT40), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(KEYINPUT40), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n540), .B2(new_n545), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n513), .B(new_n546), .C1(new_n548), .C2(KEYINPUT90), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT86), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n403), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n539), .A3(new_n417), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n553), .A3(new_n319), .ZN(new_n554));
  INV_X1    g353(.A(new_n547), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n549), .A2(new_n313), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n537), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n499), .A2(new_n510), .A3(KEYINPUT36), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT36), .B1(new_n499), .B2(new_n510), .ZN(new_n562));
  OAI22_X1  g361(.A1(new_n523), .A2(new_n520), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n512), .B(new_n527), .C1(new_n560), .C2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AND2_X1   g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT93), .ZN(new_n571));
  XOR2_X1   g370(.A(G43gat), .B(G50gat), .Z(new_n572));
  INV_X1    g371(.A(KEYINPUT15), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G29gat), .A2(G36gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT15), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT14), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT91), .A2(KEYINPUT14), .ZN(new_n582));
  OAI22_X1  g381(.A1(new_n581), .A2(new_n582), .B1(G29gat), .B2(G36gat), .ZN(new_n583));
  INV_X1    g382(.A(G29gat), .ZN(new_n584));
  INV_X1    g383(.A(G36gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n584), .B(new_n585), .C1(new_n579), .C2(new_n580), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n583), .A2(new_n589), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n578), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n577), .B1(new_n587), .B2(new_n575), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n571), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n577), .A2(new_n575), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n583), .A2(new_n589), .A3(new_n586), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n589), .B1(new_n583), .B2(new_n586), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n574), .B(new_n594), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT93), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G99gat), .B(G106gat), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n605), .A2(new_n612), .A3(new_n607), .A4(new_n608), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n591), .A2(new_n592), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(KEYINPUT17), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n601), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n593), .A2(new_n599), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n566), .A2(KEYINPUT41), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(G190gat), .B1(new_n618), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n601), .A2(new_n617), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(new_n248), .A3(new_n619), .A4(new_n620), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(G218gat), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT96), .ZN(new_n626));
  AOI21_X1  g425(.A(G218gat), .B1(new_n622), .B2(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n570), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n622), .A2(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n206), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(KEYINPUT96), .A3(new_n625), .A4(new_n569), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G57gat), .B(G64gat), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT9), .ZN(new_n634));
  INV_X1    g433(.A(G71gat), .ZN(new_n635));
  INV_X1    g434(.A(G78gat), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G71gat), .B(G78gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n639), .A3(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT21), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT95), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G183gat), .B(G211gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(G15gat), .B(G22gat), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT16), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(G1gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(G1gat), .B2(new_n651), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(G8gat), .Z(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n644), .B2(new_n643), .ZN(new_n656));
  XNOR2_X1  g455(.A(G127gat), .B(G155gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n656), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n650), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n632), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G113gat), .B(G141gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G197gat), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT11), .B(G169gat), .Z(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT12), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n669), .B(KEYINPUT13), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n591), .A2(new_n571), .A3(new_n592), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT93), .B1(new_n597), .B2(new_n598), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n655), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n654), .B(G8gat), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n593), .A2(new_n599), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n616), .B2(KEYINPUT17), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n601), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n669), .A3(new_n676), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT18), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n679), .A2(KEYINPUT18), .A3(new_n669), .A4(new_n676), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n668), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n668), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n643), .A2(new_n614), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT97), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n610), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n609), .A3(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(new_n641), .A3(new_n642), .A4(new_n613), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n688), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n641), .A4(new_n642), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(G230gat), .A2(G233gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G120gat), .B(G148gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(G176gat), .B(G204gat), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n700), .B(new_n701), .Z(new_n702));
  AND2_X1   g501(.A1(new_n688), .A2(new_n694), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n699), .B(new_n702), .C1(new_n698), .C2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n698), .ZN(new_n706));
  INV_X1    g505(.A(new_n698), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n695), .B2(new_n696), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n704), .A2(KEYINPUT98), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT98), .B1(new_n704), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n663), .A2(new_n687), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n565), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n514), .A2(new_n440), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G1gat), .ZN(G1324gat));
  INV_X1    g518(.A(new_n313), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G8gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(KEYINPUT99), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT100), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  OAI221_X1 g529(.A(new_n722), .B1(new_n721), .B2(new_n724), .C1(new_n729), .C2(new_n730), .ZN(G1325gat));
  AOI21_X1  g530(.A(G15gat), .B1(new_n715), .B2(new_n526), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n561), .A2(new_n562), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G15gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT101), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n732), .B1(new_n715), .B2(new_n735), .ZN(G1326gat));
  NAND2_X1  g535(.A1(new_n469), .A2(new_n478), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n715), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT43), .B(G22gat), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1327gat));
  INV_X1    g539(.A(new_n662), .ZN(new_n741));
  INV_X1    g540(.A(new_n687), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n741), .A2(new_n742), .A3(new_n712), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n564), .A2(new_n632), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n584), .A3(new_n717), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT45), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n628), .A2(new_n631), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n512), .A2(new_n527), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n545), .A2(new_n553), .A3(new_n319), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n750), .A2(KEYINPUT40), .B1(new_n439), .B2(new_n438), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n548), .A2(KEYINPUT90), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n556), .A2(new_n557), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n536), .B(new_n523), .C1(new_n754), .C2(new_n313), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n442), .A2(new_n737), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT36), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n524), .B2(new_n525), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n499), .A2(new_n510), .A3(KEYINPUT36), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  AOI211_X1 g560(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT44), .B1(new_n564), .B2(new_n632), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n743), .B(KEYINPUT102), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n717), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n746), .B1(new_n584), .B2(new_n766), .ZN(G1328gat));
  NAND3_X1  g566(.A1(new_n744), .A2(new_n585), .A3(new_n720), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT103), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT46), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n744), .A2(new_n771), .A3(new_n585), .A4(new_n720), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n769), .B2(new_n772), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n764), .A2(new_n720), .A3(new_n765), .ZN(new_n775));
  OAI22_X1  g574(.A1(new_n773), .A2(new_n774), .B1(new_n585), .B2(new_n775), .ZN(G1329gat));
  AND3_X1   g575(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n512), .A2(new_n527), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n632), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n747), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n564), .A2(KEYINPUT44), .A3(new_n632), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n780), .A2(new_n733), .A3(new_n781), .A4(new_n765), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT104), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n764), .A2(new_n784), .A3(new_n733), .A4(new_n765), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n785), .A3(G43gat), .ZN(new_n786));
  INV_X1    g585(.A(G43gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n744), .A2(new_n787), .A3(new_n526), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n782), .A2(G43gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n788), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n794), .ZN(G1330gat));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n737), .A3(new_n781), .A4(new_n765), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G50gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(G50gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n744), .A2(new_n800), .A3(new_n737), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT48), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n797), .B(new_n801), .C1(new_n798), .C2(KEYINPUT48), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1331gat));
  NAND3_X1  g605(.A1(new_n663), .A2(new_n742), .A3(new_n712), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n565), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n717), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n720), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n565), .A2(new_n807), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT106), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1333gat));
  AOI21_X1  g616(.A(new_n635), .B1(new_n808), .B2(new_n733), .ZN(new_n818));
  INV_X1    g617(.A(new_n526), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(G71gat), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n808), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g621(.A1(new_n808), .A2(new_n737), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g623(.A1(new_n741), .A2(new_n687), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n564), .A2(new_n632), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n564), .A2(KEYINPUT51), .A3(new_n632), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n603), .A3(new_n717), .A4(new_n712), .ZN(new_n831));
  INV_X1    g630(.A(new_n764), .ZN(new_n832));
  INV_X1    g631(.A(new_n825), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n713), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n832), .A2(new_n716), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n831), .B1(new_n836), .B2(new_n603), .ZN(G1336gat));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n720), .A2(new_n712), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(G92gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n830), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n838), .A2(new_n839), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n780), .A2(new_n720), .A3(new_n781), .A4(new_n834), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(G92gat), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n843), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n844), .B1(new_n843), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(G1337gat));
  INV_X1    g648(.A(G99gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n830), .A2(new_n850), .A3(new_n526), .A4(new_n712), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n832), .A2(new_n760), .A3(new_n835), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n850), .ZN(G1338gat));
  NAND4_X1  g652(.A1(new_n780), .A2(new_n737), .A3(new_n781), .A4(new_n834), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G106gat), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n523), .A2(G106gat), .A3(new_n713), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT53), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n855), .B(new_n859), .C1(new_n856), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1339gat));
  NOR4_X1   g663(.A1(new_n632), .A2(new_n662), .A3(new_n687), .A4(new_n712), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n695), .A2(new_n696), .A3(new_n707), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n699), .A2(KEYINPUT54), .A3(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n702), .B1(new_n708), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT55), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT109), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT109), .B(KEYINPUT55), .C1(new_n868), .C2(new_n870), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(KEYINPUT55), .A3(new_n870), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n704), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n866), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n877), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(KEYINPUT110), .C1(new_n873), .C2(new_n874), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n687), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n674), .A2(new_n676), .A3(new_n671), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n679), .A2(new_n676), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n669), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT111), .B1(new_n884), .B2(new_n667), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n669), .B1(new_n679), .B2(new_n676), .ZN(new_n886));
  INV_X1    g685(.A(new_n882), .ZN(new_n887));
  OAI211_X1 g686(.A(KEYINPUT111), .B(new_n667), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n686), .B(new_n712), .C1(new_n885), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n748), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n682), .A2(new_n668), .A3(new_n683), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n884), .A2(new_n667), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n893), .B1(new_n896), .B2(new_n888), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n632), .A2(new_n897), .A3(new_n878), .A4(new_n880), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n865), .B1(new_n899), .B2(new_n662), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n511), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n717), .A2(new_n313), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT112), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n901), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n352), .A3(new_n742), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n904), .A2(new_n742), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(G113gat), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n909), .A2(new_n911), .ZN(G1340gat));
  OAI21_X1  g711(.A(G120gat), .B1(new_n908), .B2(new_n713), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n712), .A2(new_n367), .A3(new_n369), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n904), .B2(new_n914), .ZN(G1341gat));
  NAND2_X1  g714(.A1(new_n741), .A2(G127gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n905), .B2(new_n907), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n361), .B1(new_n904), .B2(new_n662), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n921), .ZN(G1342gat));
  OAI21_X1  g721(.A(G134gat), .B1(new_n908), .B2(new_n748), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n632), .A2(new_n313), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT114), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n901), .A2(new_n359), .A3(new_n717), .A4(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT56), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n927), .ZN(G1343gat));
  NAND3_X1  g727(.A1(new_n760), .A2(new_n903), .A3(KEYINPUT115), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT115), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(new_n733), .B2(new_n902), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n523), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n877), .A2(new_n871), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n893), .B2(new_n684), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n890), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n748), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n741), .B1(new_n938), .B2(new_n898), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n934), .B1(new_n939), .B2(new_n865), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT116), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT116), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n942), .B(new_n934), .C1(new_n939), .C2(new_n865), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n632), .B1(new_n881), .B2(new_n890), .ZN(new_n945));
  AND4_X1   g744(.A1(new_n632), .A2(new_n897), .A3(new_n878), .A4(new_n880), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n662), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n865), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT57), .B1(new_n949), .B2(new_n737), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n687), .B(new_n932), .C1(new_n944), .C2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n523), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n941), .B(new_n943), .C1(new_n954), .C2(KEYINPUT57), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n955), .A2(KEYINPUT120), .A3(new_n687), .A4(new_n932), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(G141gat), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n741), .B1(new_n892), .B2(new_n898), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT117), .B(new_n717), .C1(new_n958), .C2(new_n865), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n733), .A2(new_n523), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT117), .B1(new_n949), .B2(new_n717), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT118), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT117), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n900), .B2(new_n716), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n960), .A4(new_n959), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n742), .A2(G141gat), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n963), .A2(new_n967), .A3(new_n313), .A4(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n957), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n951), .A2(G141gat), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n313), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n961), .A2(new_n962), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g773(.A(KEYINPUT58), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(G1344gat));
  INV_X1    g775(.A(KEYINPUT59), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n932), .B1(new_n944), .B2(new_n950), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n977), .B(G148gat), .C1(new_n978), .C2(new_n713), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n875), .A2(new_n877), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n632), .A2(new_n897), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n741), .B1(new_n938), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n933), .B(new_n737), .C1(new_n982), .C2(new_n865), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n954), .B2(new_n933), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n929), .A2(new_n712), .A3(new_n931), .ZN(new_n985));
  OAI21_X1  g784(.A(G148gat), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT59), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n987), .B1(new_n986), .B2(KEYINPUT59), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n979), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n713), .A2(G148gat), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n963), .A2(new_n967), .A3(new_n313), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1345gat));
  NOR2_X1   g792(.A1(new_n662), .A2(G155gat), .ZN(new_n994));
  NAND4_X1  g793(.A1(new_n963), .A2(new_n967), .A3(new_n313), .A4(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(G155gat), .B1(new_n978), .B2(new_n662), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT122), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT122), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1346gat));
  INV_X1    g800(.A(G162gat), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n963), .A2(new_n967), .A3(new_n1002), .A4(new_n925), .ZN(new_n1003));
  OAI21_X1  g802(.A(G162gat), .B1(new_n978), .B2(new_n748), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1347gat));
  NAND2_X1  g804(.A1(new_n720), .A2(new_n716), .ZN(new_n1006));
  NOR3_X1   g805(.A1(new_n900), .A2(new_n511), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(new_n687), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(G169gat), .ZN(G1348gat));
  AOI21_X1  g808(.A(new_n713), .B1(KEYINPUT123), .B2(new_n221), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n221), .A2(KEYINPUT123), .ZN(new_n1012));
  XNOR2_X1  g811(.A(new_n1011), .B(new_n1012), .ZN(G1349gat));
  INV_X1    g812(.A(new_n511), .ZN(new_n1014));
  INV_X1    g813(.A(new_n1006), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n949), .A2(new_n1014), .A3(new_n741), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(G183gat), .ZN(new_n1017));
  OAI211_X1 g816(.A(new_n1017), .B(KEYINPUT124), .C1(new_n236), .C2(new_n1016), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n1016), .A2(new_n236), .ZN(new_n1019));
  OAI21_X1  g818(.A(new_n1018), .B1(KEYINPUT124), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT60), .ZN(new_n1021));
  XNOR2_X1  g820(.A(new_n1020), .B(new_n1021), .ZN(G1350gat));
  AOI21_X1  g821(.A(new_n248), .B1(new_n1007), .B2(new_n632), .ZN(new_n1023));
  OR2_X1    g822(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(KEYINPUT61), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1007), .A2(new_n230), .A3(new_n632), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(G1351gat));
  AND2_X1   g826(.A1(new_n949), .A2(new_n960), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n1028), .A2(new_n1015), .ZN(new_n1029));
  INV_X1    g828(.A(G197gat), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1029), .A2(new_n1030), .A3(new_n687), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT125), .ZN(new_n1032));
  NOR2_X1   g831(.A1(new_n733), .A2(new_n1006), .ZN(new_n1033));
  OAI211_X1 g832(.A(new_n983), .B(new_n1033), .C1(new_n954), .C2(new_n933), .ZN(new_n1034));
  OAI21_X1  g833(.A(G197gat), .B1(new_n1034), .B2(new_n742), .ZN(new_n1035));
  AND3_X1   g834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g835(.A(new_n1032), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g836(.A1(new_n1036), .A2(new_n1037), .ZN(G1352gat));
  NOR3_X1   g837(.A1(new_n841), .A2(new_n717), .A3(G204gat), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1028), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g839(.A(new_n1040), .B(KEYINPUT62), .Z(new_n1041));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1042), .B1(new_n1034), .B2(new_n713), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1043), .A2(G204gat), .ZN(new_n1044));
  NOR3_X1   g843(.A1(new_n1034), .A2(new_n1042), .A3(new_n713), .ZN(new_n1045));
  OAI21_X1  g844(.A(new_n1041), .B1(new_n1044), .B2(new_n1045), .ZN(G1353gat));
  NAND3_X1  g845(.A1(new_n1029), .A2(new_n205), .A3(new_n741), .ZN(new_n1047));
  OR2_X1    g846(.A1(new_n1034), .A2(new_n662), .ZN(new_n1048));
  AND2_X1   g847(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n1049));
  OAI21_X1  g848(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n1050));
  INV_X1    g849(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g850(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g851(.A(new_n1052), .ZN(new_n1053));
  AOI21_X1  g852(.A(new_n1049), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1054));
  OAI21_X1  g853(.A(new_n1047), .B1(new_n1053), .B2(new_n1054), .ZN(G1354gat));
  NAND3_X1  g854(.A1(new_n1029), .A2(new_n206), .A3(new_n632), .ZN(new_n1056));
  OAI21_X1  g855(.A(G218gat), .B1(new_n1034), .B2(new_n748), .ZN(new_n1057));
  NAND2_X1  g856(.A1(new_n1056), .A2(new_n1057), .ZN(G1355gat));
endmodule


