//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988;
  INV_X1    g000(.A(G204gat), .ZN(new_n202));
  AND2_X1   g001(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT72), .ZN(new_n206));
  INV_X1    g005(.A(G197gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(G204gat), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT22), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  INV_X1    g011(.A(G218gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n205), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G211gat), .B(G218gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n205), .A2(new_n210), .A3(new_n216), .A4(new_n214), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n224), .B(new_n225), .C1(G169gat), .C2(G176gat), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n223), .A2(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NOR4_X1   g026(.A1(new_n225), .A2(KEYINPUT65), .A3(G169gat), .A4(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT65), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n222), .B2(KEYINPUT23), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT64), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n234), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n233), .A2(new_n235), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n227), .A2(new_n231), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT25), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n236), .B1(new_n239), .B2(new_n238), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n232), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n227), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT28), .ZN(new_n251));
  OR2_X1    g050(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n253));
  AOI21_X1  g052(.A(G190gat), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n257));
  NAND2_X1  g056(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n222), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT26), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n222), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263));
  OAI211_X1 g062(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n259), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G190gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n253), .ZN(new_n267));
  NOR2_X1   g066(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(KEYINPUT67), .A3(KEYINPUT28), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n256), .A2(new_n265), .A3(new_n270), .A4(new_n238), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272));
  INV_X1    g071(.A(G226gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n250), .A2(new_n271), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n242), .A2(new_n243), .B1(new_n227), .B2(new_n248), .ZN(new_n278));
  INV_X1    g077(.A(new_n271), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n278), .A2(new_n279), .A3(new_n275), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n221), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT37), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n250), .A2(new_n276), .A3(new_n271), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n276), .A2(new_n272), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n278), .B2(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n285), .A3(new_n220), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT38), .ZN(new_n288));
  XNOR2_X1  g087(.A(G8gat), .B(G36gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(G64gat), .B(G92gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n283), .A2(new_n285), .A3(new_n220), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n282), .B1(new_n293), .B2(KEYINPUT85), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n281), .A2(new_n286), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(KEYINPUT85), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n291), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n286), .A3(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n220), .B1(new_n283), .B2(new_n285), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT73), .A3(new_n297), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n292), .A2(new_n296), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G1gat), .B(G29gat), .ZN(new_n305));
  INV_X1    g104(.A(G85gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT0), .B(G57gat), .ZN(new_n308));
  XOR2_X1   g107(.A(new_n307), .B(new_n308), .Z(new_n309));
  XNOR2_X1  g108(.A(G127gat), .B(G134gat), .ZN(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G113gat), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G120gat), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI211_X1 g116(.A(KEYINPUT70), .B(KEYINPUT1), .C1(new_n312), .C2(new_n314), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G141gat), .B(G148gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n324), .B1(G155gat), .B2(G162gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G148gat), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G155gat), .B(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(G155gat), .ZN(new_n333));
  INV_X1    g132(.A(G162gat), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT2), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(new_n310), .ZN(new_n342));
  XNOR2_X1  g141(.A(G113gat), .B(G120gat), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT70), .B1(new_n343), .B2(KEYINPUT1), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n313), .A2(G120gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n311), .A2(G113gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n316), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n342), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n341), .B1(new_n349), .B2(new_n338), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n344), .A2(new_n348), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n338), .B1(new_n356), .B2(new_n310), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n337), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n357), .A2(KEYINPUT75), .A3(new_n358), .A4(new_n337), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n326), .A2(new_n336), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT74), .B1(new_n368), .B2(new_n357), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n319), .A2(new_n339), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n365), .A4(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n353), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n355), .B1(new_n364), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(new_n359), .ZN(new_n377));
  AND4_X1   g176(.A1(new_n375), .A2(new_n376), .A3(new_n352), .A4(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n309), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n309), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n369), .A2(new_n372), .B1(new_n363), .B2(new_n359), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(new_n375), .A3(new_n352), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n373), .A2(new_n364), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n380), .B(new_n382), .C1(new_n383), .C2(new_n355), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT76), .B(KEYINPUT6), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n309), .B(new_n385), .C1(new_n374), .C2(new_n378), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n302), .A2(new_n282), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n287), .A2(new_n291), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT38), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n304), .A2(new_n387), .A3(new_n388), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G228gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n215), .A2(new_n394), .A3(new_n217), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n272), .B(new_n395), .C1(new_n220), .C2(new_n394), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n337), .B1(new_n396), .B2(new_n366), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n367), .A2(new_n272), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n221), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT29), .B1(new_n218), .B2(new_n219), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n341), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT80), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n406), .B(new_n341), .C1(new_n403), .C2(KEYINPUT3), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n393), .B1(new_n221), .B2(new_n398), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n401), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n402), .B1(new_n401), .B2(new_n409), .ZN(new_n411));
  XNOR2_X1  g210(.A(G78gat), .B(G106gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G22gat), .B(G50gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT31), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n410), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n218), .A2(KEYINPUT79), .A3(new_n219), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n272), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n366), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n341), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n421), .A2(new_n399), .B1(G228gat), .B2(G233gat), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT78), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n402), .A3(new_n409), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n415), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n340), .A2(new_n350), .A3(new_n352), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT39), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT83), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT83), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n431), .A3(KEYINPUT39), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n430), .B(new_n432), .C1(new_n381), .C2(new_n352), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n376), .A2(new_n377), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n353), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n380), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT40), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n433), .A2(new_n436), .A3(KEYINPUT40), .A4(new_n380), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(new_n379), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n437), .A2(KEYINPUT84), .A3(new_n438), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT73), .B1(new_n302), .B2(new_n297), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n298), .A2(new_n299), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n298), .A2(new_n446), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n302), .A2(new_n297), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n392), .B(new_n427), .C1(new_n445), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n452), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n456), .A2(new_n441), .A3(new_n444), .A4(new_n443), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n457), .A2(new_n458), .A3(new_n427), .A4(new_n392), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n250), .A2(new_n370), .A3(new_n271), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n357), .B1(new_n278), .B2(new_n279), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n462), .A2(new_n463), .A3(G227gat), .A4(G233gat), .ZN(new_n464));
  XOR2_X1   g263(.A(G15gat), .B(G43gat), .Z(new_n465));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT33), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(KEYINPUT32), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT71), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n464), .A2(KEYINPUT71), .A3(KEYINPUT32), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n464), .A2(KEYINPUT32), .ZN(new_n474));
  INV_X1    g273(.A(new_n464), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n467), .C1(new_n475), .C2(KEYINPUT33), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n462), .A2(new_n463), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n478));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n482), .B1(new_n473), .B2(new_n476), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n461), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n476), .ZN(new_n486));
  INV_X1    g285(.A(new_n482), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n473), .A2(new_n476), .A3(new_n482), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(KEYINPUT36), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n379), .A2(new_n384), .A3(new_n492), .A4(new_n386), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n493), .A2(new_n388), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n456), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n417), .B2(new_n426), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n416), .B1(new_n410), .B2(new_n411), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n424), .A2(new_n425), .A3(new_n415), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT81), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT82), .B(new_n491), .C1(new_n496), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT82), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n495), .A2(new_n388), .A3(new_n493), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(new_n453), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n485), .A2(new_n490), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n460), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n488), .A2(new_n489), .ZN(new_n510));
  INV_X1    g309(.A(new_n427), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n387), .A2(new_n388), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n509), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT87), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n509), .A2(new_n521), .A3(new_n518), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(KEYINPUT41), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G29gat), .A2(G36gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT89), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n536), .A2(G29gat), .A3(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT90), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n538), .B(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G43gat), .B(G50gat), .Z(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n542), .A3(new_n533), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT91), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n551), .B2(new_n552), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT96), .B(G85gat), .Z(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(G99gat), .ZN(new_n562));
  INV_X1    g361(.A(G106gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT8), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n306), .B2(new_n559), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n560), .A2(new_n561), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n552), .B2(new_n551), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n557), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n569), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(new_n551), .B1(KEYINPUT41), .B2(new_n524), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n530), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n573), .B(new_n529), .C1(new_n557), .C2(new_n570), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n575), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n528), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(new_n527), .A3(new_n579), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G15gat), .B(G22gat), .ZN(new_n587));
  INV_X1    g386(.A(G1gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT16), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(G1gat), .B2(new_n587), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(G8gat), .ZN(new_n592));
  XOR2_X1   g391(.A(G57gat), .B(G64gat), .Z(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G71gat), .B(G78gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT95), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n592), .B1(new_n600), .B2(KEYINPUT21), .ZN(new_n601));
  XOR2_X1   g400(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G127gat), .B(G155gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n603), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G183gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n607), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n606), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n586), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n551), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n592), .B1(new_n617), .B2(KEYINPUT17), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(new_n554), .B2(new_n556), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n592), .A2(new_n551), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n619), .A2(KEYINPUT18), .A3(new_n620), .A4(new_n621), .ZN(new_n625));
  INV_X1    g424(.A(G8gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n591), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n551), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n620), .B(KEYINPUT13), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT11), .B(G169gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT88), .Z(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n631), .B1(new_n624), .B2(KEYINPUT92), .ZN(new_n640));
  INV_X1    g439(.A(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n622), .A2(new_n623), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT92), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT93), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT93), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n647), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n639), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n569), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT99), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n599), .B(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n650), .B(new_n652), .C1(new_n654), .C2(new_n569), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n600), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n652), .B1(new_n654), .B2(new_n569), .ZN(new_n660));
  INV_X1    g459(.A(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n659), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n666), .B1(new_n659), .B2(new_n662), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n616), .A2(new_n649), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n523), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n505), .A2(KEYINPUT100), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n505), .A2(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT101), .B(G1gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n523), .A2(new_n456), .A3(new_n672), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n681), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT102), .B(new_n681), .C1(new_n682), .C2(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n682), .A2(G8gat), .ZN(new_n690));
  INV_X1    g489(.A(new_n673), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n691), .A2(KEYINPUT42), .A3(new_n456), .A4(new_n683), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n689), .B(new_n690), .C1(new_n694), .C2(new_n695), .ZN(G1325gat));
  AND3_X1   g495(.A1(new_n691), .A2(G15gat), .A3(new_n507), .ZN(new_n697));
  INV_X1    g496(.A(new_n510), .ZN(new_n698));
  AOI21_X1  g497(.A(G15gat), .B1(new_n691), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n673), .A2(new_n502), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n649), .ZN(new_n704));
  INV_X1    g503(.A(new_n615), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n670), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n586), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n677), .A2(G29gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n523), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n523), .A2(new_n711), .A3(new_n707), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  INV_X1    g513(.A(new_n518), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n505), .A2(new_n453), .ZN(new_n716));
  INV_X1    g515(.A(new_n502), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n716), .A2(new_n717), .B1(new_n490), .B2(new_n485), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n437), .A2(KEYINPUT84), .A3(new_n438), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT84), .B1(new_n437), .B2(new_n438), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n442), .A2(new_n379), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n511), .B1(new_n722), .B2(new_n456), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n458), .B1(new_n723), .B2(new_n392), .ZN(new_n724));
  AND4_X1   g523(.A1(new_n458), .A2(new_n457), .A3(new_n427), .A4(new_n392), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n718), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n460), .A2(KEYINPUT105), .A3(new_n718), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n715), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n714), .B1(new_n730), .B2(new_n586), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n586), .A2(new_n714), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n520), .A2(new_n522), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n706), .B(KEYINPUT104), .Z(new_n734));
  NAND4_X1  g533(.A1(new_n731), .A2(new_n676), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G29gat), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n713), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1328gat));
  NOR2_X1   g540(.A1(new_n453), .A2(G36gat), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n520), .A2(new_n522), .A3(new_n707), .A4(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n731), .A2(new_n456), .A3(new_n733), .A4(new_n734), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT109), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n752), .B(new_n745), .C1(new_n748), .C2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1329gat));
  AND2_X1   g553(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n510), .A2(G43gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n520), .A2(new_n522), .A3(new_n707), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT110), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n731), .A2(new_n507), .A3(new_n733), .A4(new_n734), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G43gat), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n755), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT111), .A2(KEYINPUT47), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1330gat));
  AND2_X1   g562(.A1(new_n731), .A2(new_n733), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n764), .A2(new_n511), .A3(new_n734), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n523), .A2(new_n707), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n502), .A2(G50gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(KEYINPUT48), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n764), .A2(new_n717), .A3(new_n734), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n769), .B1(new_n772), .B2(G50gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(KEYINPUT48), .B2(new_n773), .ZN(G1331gat));
  NOR2_X1   g573(.A1(new_n704), .A2(new_n670), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n730), .A2(new_n616), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n676), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g578(.A(new_n453), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT112), .ZN(new_n782));
  NOR2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(G1333gat));
  NAND3_X1  g583(.A1(new_n777), .A2(G71gat), .A3(new_n507), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n777), .A2(new_n698), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G71gat), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g587(.A1(new_n777), .A2(new_n717), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT113), .B(G78gat), .Z(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1335gat));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n615), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n764), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(new_n558), .A3(new_n677), .ZN(new_n794));
  INV_X1    g593(.A(new_n729), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT105), .B1(new_n460), .B2(new_n718), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n518), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  AOI211_X1 g598(.A(new_n615), .B(new_n704), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n797), .A2(new_n585), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n802), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n797), .A2(new_n585), .A3(new_n804), .A4(new_n800), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(new_n671), .A3(new_n676), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n794), .B1(new_n558), .B2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n731), .A2(new_n456), .A3(new_n733), .A4(new_n792), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G92gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(KEYINPUT116), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n671), .A2(new_n559), .A3(new_n456), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT115), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n803), .A2(new_n805), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n811), .B(new_n815), .ZN(G1337gat));
  NOR3_X1   g615(.A1(new_n793), .A2(new_n562), .A3(new_n491), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n803), .A2(new_n698), .A3(new_n671), .A4(new_n805), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n562), .B2(new_n818), .ZN(G1338gat));
  OAI21_X1  g618(.A(G106gat), .B1(new_n793), .B2(new_n427), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n427), .A2(G106gat), .ZN(new_n821));
  AND4_X1   g620(.A1(new_n671), .A2(new_n803), .A3(new_n805), .A4(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n731), .A2(new_n717), .A3(new_n733), .A4(new_n792), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n826), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT117), .B1(new_n826), .B2(G106gat), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n827), .A2(new_n822), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n655), .A2(new_n661), .A3(new_n656), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n659), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n661), .B1(new_n655), .B2(new_n656), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n666), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n667), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n833), .A2(new_n836), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n649), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n628), .A2(new_n629), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT119), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n619), .A2(new_n621), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(G229gat), .A3(G233gat), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n636), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n670), .B(new_n850), .C1(new_n646), .C2(new_n648), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n586), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n646), .A2(new_n648), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n838), .B1(new_n841), .B2(new_n840), .ZN(new_n854));
  INV_X1    g653(.A(new_n850), .ZN(new_n855));
  AND4_X1   g654(.A1(new_n853), .A2(new_n854), .A3(new_n585), .A4(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n615), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n616), .A2(new_n704), .A3(new_n671), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n717), .A2(new_n510), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n677), .A2(new_n456), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n704), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G113gat), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n860), .A2(new_n510), .A3(new_n511), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n863), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n649), .A2(G113gat), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT120), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(G1340gat));
  INV_X1    g670(.A(new_n868), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n311), .A3(new_n671), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n864), .A2(new_n671), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n873), .B1(new_n875), .B2(new_n311), .ZN(G1341gat));
  NAND3_X1  g675(.A1(new_n864), .A2(G127gat), .A3(new_n615), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT121), .ZN(new_n878));
  AOI21_X1  g677(.A(G127gat), .B1(new_n872), .B2(new_n615), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  OR2_X1    g679(.A1(new_n586), .A2(G134gat), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n868), .A2(KEYINPUT56), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n585), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(G134gat), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT56), .B1(new_n868), .B2(new_n881), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n863), .A2(new_n491), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n717), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(new_n859), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n853), .A2(new_n671), .A3(new_n855), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n840), .B2(new_n841), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT123), .B(KEYINPUT55), .C1(new_n833), .C2(new_n836), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n839), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n649), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n856), .B1(new_n895), .B2(new_n586), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n615), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n649), .A2(new_n894), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n585), .B1(new_n900), .B2(new_n890), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n705), .B1(new_n901), .B2(new_n856), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n888), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g703(.A(KEYINPUT122), .B(KEYINPUT57), .Z(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n860), .B2(new_n427), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n887), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n327), .B1(new_n908), .B2(new_n704), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n860), .A2(new_n427), .ZN(new_n910));
  INV_X1    g709(.A(new_n887), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n704), .A2(new_n327), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT58), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n914), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n649), .B(new_n887), .C1(new_n904), .C2(new_n907), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n327), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(new_n912), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n921), .A2(new_n329), .A3(new_n671), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT59), .B(new_n329), .C1(new_n908), .C2(new_n671), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n511), .B(new_n905), .C1(new_n858), .C2(new_n859), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n502), .B1(new_n902), .B2(new_n889), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(KEYINPUT57), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n671), .A3(new_n911), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n922), .B1(new_n923), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n921), .B2(new_n615), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n705), .A2(new_n333), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n908), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n921), .B2(new_n585), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n586), .A2(new_n334), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n908), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n676), .A2(new_n453), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n867), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G169gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n704), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n937), .A2(new_n862), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n861), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n704), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n941), .B1(new_n940), .B2(new_n946), .ZN(G1348gat));
  AOI21_X1  g746(.A(G176gat), .B1(new_n939), .B2(new_n671), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n671), .A2(G176gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n944), .B2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n943), .B2(new_n705), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n615), .B1(new_n268), .B2(new_n267), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n938), .B2(new_n952), .ZN(new_n953));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n953), .B(new_n954), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n943), .B2(new_n586), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n266), .A3(new_n585), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  NAND2_X1  g758(.A1(new_n937), .A2(new_n491), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n910), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n207), .A3(new_n704), .ZN(new_n964));
  INV_X1    g763(.A(new_n927), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n965), .A2(new_n649), .A3(new_n960), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n966), .B2(new_n207), .ZN(G1352gat));
  NOR2_X1   g766(.A1(new_n670), .A2(G204gat), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n962), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n962), .B2(new_n969), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n965), .A2(new_n670), .A3(new_n960), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n970), .B(new_n971), .C1(new_n972), .C2(new_n202), .ZN(G1353gat));
  AND4_X1   g772(.A1(new_n212), .A2(new_n910), .A3(new_n615), .A4(new_n961), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT126), .Z(new_n975));
  INV_X1    g774(.A(new_n925), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n889), .B1(new_n896), .B2(new_n615), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT57), .B1(new_n977), .B2(new_n717), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n615), .B(new_n961), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n212), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n927), .A2(KEYINPUT127), .A3(new_n615), .A4(new_n961), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n981), .A2(KEYINPUT63), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n981), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n975), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n963), .B2(new_n585), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n965), .A2(new_n960), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n586), .A2(new_n213), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(G1355gat));
endmodule


