//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(new_n202), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n205), .A2(new_n208), .A3(KEYINPUT70), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n215));
  INV_X1    g014(.A(G169gat), .ZN(new_n216));
  INV_X1    g015(.A(G176gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n217), .ZN(new_n220));
  AND2_X1   g019(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n221));
  NOR2_X1   g020(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(KEYINPUT65), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n225), .B2(new_n220), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n218), .B1(new_n231), .B2(new_n223), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G183gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n236), .A2(new_n238), .A3(KEYINPUT24), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n228), .A2(new_n234), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT25), .ZN(new_n244));
  NOR3_X1   g043(.A1(new_n240), .A2(new_n244), .A3(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n232), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT67), .A3(new_n245), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n243), .A2(new_n244), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT27), .B(G183gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n238), .ZN(new_n252));
  OR2_X1    g051(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n252), .A2(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n214), .A2(KEYINPUT69), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n256), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(KEYINPUT26), .B2(new_n256), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n213), .B1(new_n250), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G227gat), .ZN(new_n262));
  INV_X1    g061(.A(G233gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n213), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n248), .A2(new_n249), .ZN(new_n266));
  INV_X1    g065(.A(new_n242), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(new_n227), .B2(KEYINPUT66), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT25), .B1(new_n268), .B2(new_n234), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n265), .B(new_n259), .C1(new_n266), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n261), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT33), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n277), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT71), .B1(new_n281), .B2(new_n282), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n234), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n242), .B1(new_n232), .B2(new_n233), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n244), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n248), .A2(new_n249), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n260), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(new_n265), .ZN(new_n291));
  AOI211_X1 g090(.A(new_n260), .B(new_n213), .C1(new_n288), .C2(new_n289), .ZN(new_n292));
  OAI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(new_n262), .B2(new_n263), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT34), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  OAI221_X1 g094(.A(new_n295), .B1(new_n262), .B2(new_n263), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n294), .A2(new_n296), .A3(new_n280), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n283), .B2(new_n284), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n298), .B(KEYINPUT73), .C1(new_n283), .C2(new_n284), .ZN(new_n302));
  AOI221_X4 g101(.A(KEYINPUT36), .B1(new_n285), .B2(new_n297), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n297), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(new_n263), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n290), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT74), .B(new_n313), .C1(new_n250), .C2(new_n260), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  XNOR2_X1  g117(.A(G197gat), .B(G204gat), .ZN(new_n319));
  INV_X1    g118(.A(G211gat), .ZN(new_n320));
  INV_X1    g119(.A(G218gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(KEYINPUT22), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G211gat), .B(G218gat), .Z(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n259), .B1(new_n266), .B2(new_n269), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n326), .B1(new_n329), .B2(new_n314), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n317), .A2(new_n318), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n314), .B1(new_n290), .B2(KEYINPUT29), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n332), .A2(new_n315), .A3(new_n316), .A4(new_n325), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT37), .ZN(new_n335));
  INV_X1    g134(.A(new_n332), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n290), .A2(new_n314), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n326), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT76), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  NAND2_X1  g142(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  AND4_X1   g143(.A1(new_n315), .A2(new_n332), .A3(new_n316), .A4(new_n325), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n332), .B1(new_n290), .B2(new_n314), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(new_n318), .B1(new_n326), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n335), .B1(new_n347), .B2(new_n334), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n310), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(G141gat), .ZN(new_n350));
  INV_X1    g149(.A(G148gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G155gat), .ZN(new_n355));
  INV_X1    g154(.A(G162gat), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT2), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358));
  XNOR2_X1  g157(.A(G155gat), .B(G162gat), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n354), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n352), .A3(new_n353), .ZN(new_n361));
  INV_X1    g160(.A(new_n359), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n358), .A3(new_n353), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n211), .B2(new_n212), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT80), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n365), .B2(new_n209), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n365), .A2(new_n209), .A3(new_n369), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n368), .B1(new_n373), .B2(new_n367), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT78), .B1(new_n365), .B2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT78), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n360), .A2(new_n364), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n209), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(KEYINPUT3), .B2(new_n365), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n384), .B(KEYINPUT79), .Z(new_n385));
  NOR2_X1   g184(.A1(new_n385), .A2(KEYINPUT5), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n374), .A2(new_n375), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n365), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n381), .A3(KEYINPUT80), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n367), .B1(new_n389), .B2(new_n370), .ZN(new_n390));
  AOI211_X1 g189(.A(KEYINPUT4), .B(new_n365), .C1(new_n211), .C2(new_n212), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n383), .B(new_n386), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT82), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n385), .B1(new_n366), .B2(KEYINPUT4), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n395), .B(new_n383), .C1(new_n373), .C2(KEYINPUT4), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT5), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n365), .A2(KEYINPUT81), .A3(new_n209), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT81), .B1(new_n365), .B2(new_n209), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n371), .A2(new_n372), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(new_n385), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n387), .A2(new_n393), .B1(new_n396), .B2(new_n401), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n407), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n410), .A2(new_n407), .A3(new_n412), .ZN(new_n414));
  INV_X1    g213(.A(new_n343), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n331), .A2(new_n334), .A3(new_n338), .A4(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n335), .B1(new_n346), .B2(new_n325), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n317), .A2(new_n326), .A3(new_n332), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n310), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n339), .A3(new_n343), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n349), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G78gat), .B(G106gat), .Z(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT31), .B(G50gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT86), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n325), .B1(new_n380), .B2(new_n328), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n325), .A2(new_n328), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n388), .B1(new_n429), .B2(new_n378), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G228gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(new_n263), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n427), .B(G22gat), .C1(new_n428), .C2(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n433), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n426), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n425), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n444), .A3(new_n438), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n416), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n343), .A2(new_n447), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n347), .A2(new_n334), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n338), .B1(new_n333), .B2(KEYINPUT75), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n318), .B1(new_n317), .B2(new_n330), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n343), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n374), .A2(new_n383), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n385), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n400), .A2(new_n385), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n458), .A3(new_n385), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n407), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n460), .A2(KEYINPUT40), .A3(new_n407), .A4(new_n461), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n409), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n446), .B1(new_n454), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n412), .B1(new_n410), .B2(new_n407), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n394), .A2(new_n407), .A3(new_n402), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n409), .A2(KEYINPUT84), .A3(new_n411), .A4(new_n412), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n414), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n473), .A2(new_n448), .A3(new_n450), .A4(new_n453), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n422), .A2(new_n467), .B1(new_n474), .B2(new_n446), .ZN(new_n475));
  INV_X1    g274(.A(new_n454), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n446), .B1(new_n285), .B2(new_n297), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n305), .A2(new_n476), .A3(new_n473), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT35), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n413), .A2(new_n414), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n454), .A2(new_n480), .A3(KEYINPUT35), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n305), .A3(new_n477), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n308), .A2(new_n475), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G36gat), .ZN(new_n484));
  AND2_X1   g283(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(G29gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n492));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n492), .A2(new_n493), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT89), .ZN(new_n499));
  INV_X1    g298(.A(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT17), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(G1gat), .ZN(new_n503));
  AOI21_X1  g302(.A(G8gat), .B1(new_n503), .B2(KEYINPUT90), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(G1gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n504), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n499), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n500), .A2(new_n508), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(KEYINPUT18), .A3(new_n513), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n508), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(new_n513), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n524), .A4(new_n531), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n483), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n471), .A2(new_n472), .A3(new_n414), .ZN(new_n538));
  XOR2_X1   g337(.A(G57gat), .B(G64gat), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT9), .ZN(new_n540));
  INV_X1    g339(.A(G71gat), .ZN(new_n541));
  INV_X1    g340(.A(G78gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n539), .A2(new_n543), .B1(new_n544), .B2(KEYINPUT93), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(KEYINPUT93), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(G127gat), .Z(new_n551));
  INV_X1    g350(.A(new_n547), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT21), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n508), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n551), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G155gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(G183gat), .B(G211gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n555), .B(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G134gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n356), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT7), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT94), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(G99gat), .B(G106gat), .Z(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n571), .B(KEYINPUT94), .ZN(new_n576));
  INV_X1    g375(.A(new_n574), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n579), .A2(new_n496), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n501), .A2(new_n575), .A3(new_n578), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n580), .B1(new_n499), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n564), .B1(new_n584), .B2(KEYINPUT95), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n582), .B(new_n583), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n579), .A2(new_n547), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n552), .B1(new_n575), .B2(new_n578), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G230gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n595), .A2(new_n263), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(new_n591), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n597), .ZN(new_n600));
  XOR2_X1   g399(.A(G120gat), .B(G148gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT96), .ZN(new_n602));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  OR2_X1    g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n560), .A2(new_n589), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n537), .A2(new_n538), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT97), .B(G1gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(G1324gat));
  INV_X1    g410(.A(new_n608), .ZN(new_n612));
  NOR4_X1   g411(.A1(new_n483), .A2(new_n476), .A3(new_n536), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT16), .B(G8gat), .Z(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(G8gat), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT42), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT42), .B2(new_n615), .ZN(G1325gat));
  NAND2_X1  g418(.A1(new_n537), .A2(new_n608), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n308), .B(KEYINPUT98), .ZN(new_n621));
  OAI21_X1  g420(.A(G15gat), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n281), .A2(new_n282), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT71), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n282), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT73), .B1(new_n627), .B2(new_n298), .ZN(new_n628));
  INV_X1    g427(.A(new_n302), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n306), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n612), .A2(G15gat), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n537), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT99), .ZN(G1326gat));
  INV_X1    g433(.A(new_n446), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT43), .B(G22gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(new_n607), .ZN(new_n639));
  AND4_X1   g438(.A1(new_n537), .A2(new_n589), .A3(new_n560), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n488), .A3(new_n538), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT100), .B(KEYINPUT45), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644));
  INV_X1    g443(.A(new_n589), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n483), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n630), .A2(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n454), .A2(new_n466), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n339), .A2(new_n343), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT37), .B1(new_n451), .B2(new_n452), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n309), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n421), .A2(new_n413), .A3(new_n414), .A4(new_n416), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n648), .B(new_n635), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n305), .A2(new_n304), .A3(new_n306), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n474), .A2(new_n446), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n647), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n305), .A2(new_n477), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n657), .A2(new_n481), .B1(new_n478), .B2(KEYINPUT35), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT44), .B(new_n589), .C1(new_n656), .C2(new_n658), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n607), .B(KEYINPUT101), .Z(new_n661));
  INV_X1    g460(.A(new_n560), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n661), .A2(new_n536), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n473), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n643), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT102), .Z(G1328gat));
  NAND3_X1  g466(.A1(new_n640), .A2(new_n484), .A3(new_n454), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT46), .Z(new_n669));
  OAI21_X1  g468(.A(G36gat), .B1(new_n664), .B2(new_n476), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(G1329gat));
  OAI21_X1  g470(.A(G43gat), .B1(new_n664), .B2(new_n308), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n630), .A2(G43gat), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n640), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(KEYINPUT47), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n621), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n676), .A3(new_n663), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n677), .A2(G43gat), .B1(new_n640), .B2(new_n673), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(G1330gat));
  NOR2_X1   g479(.A1(new_n635), .A2(G50gat), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n640), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n646), .A2(new_n446), .A3(new_n659), .A4(new_n663), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(G50gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(KEYINPUT48), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT104), .B(KEYINPUT48), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n684), .A2(KEYINPUT105), .B1(new_n640), .B2(new_n681), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n683), .A2(new_n689), .A3(G50gat), .ZN(new_n690));
  AOI211_X1 g489(.A(KEYINPUT106), .B(new_n687), .C1(new_n688), .C2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n684), .A2(KEYINPUT105), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n690), .A3(new_n682), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(new_n686), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n685), .B1(new_n691), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT107), .B(new_n685), .C1(new_n691), .C2(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1331gat));
  NAND4_X1  g499(.A1(new_n661), .A2(new_n536), .A3(new_n645), .A4(new_n662), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n483), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n483), .B2(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n538), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g507(.A(new_n476), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT109), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1333gat));
  OAI21_X1  g512(.A(G71gat), .B1(new_n705), .B2(new_n621), .ZN(new_n714));
  INV_X1    g513(.A(new_n630), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n541), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n714), .B1(new_n705), .B2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g517(.A1(new_n705), .A2(new_n635), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT110), .B(G78gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1335gat));
  OAI21_X1  g520(.A(new_n589), .B1(new_n656), .B2(new_n658), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n662), .A2(new_n535), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(KEYINPUT51), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n639), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n568), .A3(new_n538), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n724), .A2(new_n639), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n660), .A2(KEYINPUT111), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n646), .A2(new_n659), .A3(new_n730), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n731), .A2(new_n538), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n729), .B1(new_n568), .B2(new_n735), .ZN(G1336gat));
  NAND3_X1  g535(.A1(new_n660), .A2(new_n454), .A3(new_n730), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n569), .B1(new_n737), .B2(KEYINPUT112), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(KEYINPUT112), .B2(new_n737), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n726), .A2(new_n727), .ZN(new_n740));
  INV_X1    g539(.A(new_n661), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(new_n476), .A3(G92gat), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n731), .A2(new_n454), .A3(new_n734), .ZN(new_n746));
  AOI22_X1  g545(.A1(new_n746), .A2(G92gat), .B1(new_n740), .B2(new_n742), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(new_n745), .B2(new_n747), .ZN(G1337gat));
  INV_X1    g547(.A(G99gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n728), .A2(new_n749), .A3(new_n715), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n731), .A2(new_n676), .A3(new_n734), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(G1338gat));
  NOR3_X1   g551(.A1(new_n741), .A2(G106gat), .A3(new_n635), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n740), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  OAI21_X1  g554(.A(G106gat), .B1(new_n732), .B2(new_n635), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n731), .A2(new_n446), .A3(new_n734), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n758), .A2(G106gat), .B1(new_n740), .B2(new_n753), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n759), .B2(new_n755), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n305), .A2(new_n477), .ZN(new_n763));
  INV_X1    g562(.A(new_n604), .ZN(new_n764));
  INV_X1    g563(.A(new_n598), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n592), .A2(new_n593), .A3(new_n596), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n598), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n767), .A2(KEYINPUT55), .A3(new_n769), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n605), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n535), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n512), .A2(new_n513), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n521), .A2(new_n523), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n530), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n534), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n607), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n589), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n776), .A2(new_n589), .A3(new_n783), .A4(new_n778), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n560), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n608), .A2(new_n536), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n763), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n454), .A2(new_n473), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n535), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G113gat), .ZN(G1340gat));
  INV_X1    g593(.A(G120gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n792), .B2(new_n661), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(KEYINPUT115), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n795), .A3(new_n607), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1341gat));
  NAND2_X1  g598(.A1(new_n792), .A2(new_n662), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G127gat), .ZN(G1342gat));
  NOR4_X1   g600(.A1(new_n645), .A2(G134gat), .A3(new_n473), .A4(new_n454), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT56), .Z(new_n804));
  NAND2_X1  g603(.A1(new_n792), .A2(new_n589), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G134gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT116), .ZN(G1343gat));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n308), .A2(new_n791), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n789), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT57), .B1(new_n811), .B2(new_n446), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n635), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n535), .A2(new_n778), .A3(new_n772), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n589), .B1(new_n816), .B2(new_n784), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n786), .B1(new_n817), .B2(KEYINPUT117), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n560), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n820), .B2(new_n789), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n810), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G141gat), .B1(new_n822), .B2(new_n536), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n809), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n811), .A2(new_n446), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n473), .A3(new_n676), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n476), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n535), .A2(new_n350), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n825), .B(new_n830), .ZN(G1344gat));
  NAND4_X1  g630(.A1(new_n827), .A2(new_n351), .A3(new_n476), .A4(new_n607), .ZN(new_n832));
  XOR2_X1   g631(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n833));
  NAND2_X1  g632(.A1(new_n810), .A2(new_n607), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n815), .B1(new_n788), .B2(new_n789), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n778), .A2(new_n589), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n774), .B1(new_n770), .B2(new_n771), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT114), .B(KEYINPUT55), .C1(new_n767), .C2(new_n769), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n836), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n776), .A2(KEYINPUT121), .A3(new_n589), .A4(new_n778), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n783), .ZN(new_n843));
  INV_X1    g642(.A(new_n817), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n662), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n789), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n446), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n813), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n835), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n848), .A2(KEYINPUT122), .A3(new_n813), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n834), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n351), .B1(new_n853), .B2(KEYINPUT123), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n849), .A2(new_n850), .ZN(new_n856));
  INV_X1    g655(.A(new_n835), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n856), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n855), .B1(new_n858), .B2(new_n834), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n833), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n822), .A2(new_n639), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n862), .A2(KEYINPUT59), .A3(new_n351), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n832), .B1(new_n860), .B2(new_n863), .ZN(G1345gat));
  OAI21_X1  g663(.A(G155gat), .B1(new_n822), .B2(new_n560), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n662), .A2(new_n355), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n828), .B2(new_n866), .ZN(G1346gat));
  OAI21_X1  g666(.A(G162gat), .B1(new_n822), .B2(new_n645), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n827), .A2(new_n356), .A3(new_n476), .A4(new_n589), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1347gat));
  NOR2_X1   g669(.A1(new_n476), .A2(new_n538), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n790), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n536), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(new_n216), .ZN(G1348gat));
  OAI21_X1  g673(.A(G176gat), .B1(new_n872), .B2(new_n741), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n607), .A2(new_n217), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n872), .B2(new_n876), .ZN(G1349gat));
  INV_X1    g676(.A(new_n872), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n662), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n236), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n251), .B2(new_n879), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n589), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n238), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n885), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n886), .B(new_n887), .C1(G190gat), .C2(new_n883), .ZN(G1351gat));
  NAND2_X1  g687(.A1(new_n621), .A2(new_n871), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n826), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g689(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(KEYINPUT125), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G197gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n535), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n851), .A2(new_n852), .ZN(new_n897));
  INV_X1    g696(.A(new_n889), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n896), .B1(new_n899), .B2(new_n536), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G197gat), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n899), .A2(new_n896), .A3(new_n536), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n895), .B1(new_n901), .B2(new_n902), .ZN(G1352gat));
  OAI21_X1  g702(.A(G204gat), .B1(new_n899), .B2(new_n741), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n826), .A2(G204gat), .A3(new_n639), .A4(new_n889), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT62), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1353gat));
  NAND3_X1  g706(.A1(new_n893), .A2(new_n320), .A3(new_n662), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n897), .A2(new_n662), .A3(new_n898), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n909), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT63), .B1(new_n909), .B2(G211gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1354gat));
  NOR3_X1   g711(.A1(new_n899), .A2(new_n321), .A3(new_n645), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n891), .A2(new_n589), .A3(new_n892), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n321), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT127), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n917), .A3(new_n321), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n913), .B1(new_n916), .B2(new_n918), .ZN(G1355gat));
endmodule


