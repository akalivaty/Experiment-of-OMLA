//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT3), .B1(new_n187), .B2(G107), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT75), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  OAI211_X1 g004(.A(KEYINPUT75), .B(KEYINPUT3), .C1(new_n187), .C2(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT76), .A4(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  OR3_X1    g013(.A1(new_n194), .A2(KEYINPUT77), .A3(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT77), .B1(new_n194), .B2(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n192), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT78), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n192), .A2(new_n199), .A3(KEYINPUT78), .A4(new_n202), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G101), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G101), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n192), .A2(new_n199), .A3(new_n208), .A4(new_n202), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  XNOR2_X1  g026(.A(G143), .B(G146), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT64), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n212), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n226));
  NAND4_X1  g040(.A1(new_n205), .A2(G101), .A3(new_n206), .A4(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G137), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT11), .A3(G134), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n231), .A2(new_n234), .A3(new_n237), .A4(new_n232), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n217), .A3(new_n219), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n218), .A2(KEYINPUT1), .A3(G146), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n242), .B(new_n243), .C1(G128), .C2(new_n213), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n187), .A2(G107), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n194), .A2(G104), .ZN(new_n246));
  OAI21_X1  g060(.A(G101), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n209), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT80), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(KEYINPUT80), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n248), .B2(new_n250), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n228), .A2(new_n239), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n236), .A2(new_n238), .ZN(new_n255));
  INV_X1    g069(.A(new_n248), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n244), .B1(new_n209), .B2(new_n247), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT12), .B1(new_n255), .B2(KEYINPUT81), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI221_X1 g074(.A(new_n255), .B1(KEYINPUT81), .B2(KEYINPUT12), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n254), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n228), .A2(new_n239), .A3(new_n253), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n239), .B1(new_n228), .B2(new_n253), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n274), .B2(new_n270), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT83), .A2(G469), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT83), .A2(G469), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n275), .A2(new_n276), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n270), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n272), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n270), .B1(new_n254), .B2(new_n262), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT82), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n254), .A2(new_n262), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n228), .A2(new_n253), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n255), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(new_n254), .A3(new_n270), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n280), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n295), .A2(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G221), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT92), .ZN(new_n300));
  AOI21_X1  g114(.A(G237), .B1(new_n264), .B2(new_n266), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G143), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n218), .A2(KEYINPUT89), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n301), .A2(G214), .A3(new_n305), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n301), .A2(G214), .B1(new_n302), .B2(G143), .ZN(new_n307));
  OAI211_X1 g121(.A(KEYINPUT18), .B(G131), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(G125), .B(G140), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n309), .B(new_n216), .ZN(new_n310));
  INV_X1    g124(.A(G237), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n267), .A2(G214), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n303), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n301), .A2(G214), .A3(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n237), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n308), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT19), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n309), .A2(new_n318), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n216), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(new_n309), .B2(KEYINPUT16), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G146), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n313), .A2(new_n314), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(new_n237), .A3(new_n314), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT90), .B1(new_n317), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G113), .B(G122), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(G104), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT90), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n308), .A2(new_n310), .A3(new_n316), .ZN(new_n335));
  INV_X1    g149(.A(new_n329), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n237), .B1(new_n313), .B2(new_n314), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n334), .B(new_n335), .C1(new_n338), .C2(new_n326), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n331), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n328), .A2(new_n341), .A3(new_n329), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n324), .B(new_n216), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n342), .B(new_n343), .C1(new_n341), .C2(new_n328), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n333), .B(KEYINPUT91), .Z(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n335), .A3(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(G475), .B(G902), .C1(new_n340), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n300), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n346), .ZN(new_n350));
  INV_X1    g164(.A(G475), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(new_n351), .A3(new_n276), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT92), .A3(KEYINPUT20), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(new_n348), .A3(new_n351), .A4(new_n276), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n218), .A2(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n240), .A2(G143), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT95), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(KEYINPUT95), .ZN(new_n360));
  AOI21_X1  g174(.A(G134), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G122), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G116), .ZN(new_n364));
  INV_X1    g178(.A(G116), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G122), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(G107), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n240), .A2(G143), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n357), .B1(new_n369), .B2(KEYINPUT13), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT94), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(KEYINPUT13), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n373), .B(new_n357), .C1(new_n369), .C2(KEYINPUT13), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n362), .B(new_n368), .C1(new_n375), .C2(new_n230), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n364), .A2(new_n366), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT96), .B1(new_n377), .B2(new_n194), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT96), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n367), .A2(new_n379), .A3(G107), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n364), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n384));
  OAI21_X1  g198(.A(G107), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n359), .A2(G134), .A3(new_n360), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n381), .B(new_n385), .C1(new_n386), .C2(new_n361), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n376), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n295), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT97), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n376), .A2(new_n387), .A3(new_n390), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n376), .A2(new_n387), .A3(KEYINPUT97), .A4(new_n390), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n276), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT93), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n344), .A2(new_n335), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(new_n333), .ZN(new_n403));
  INV_X1    g217(.A(new_n333), .ZN(new_n404));
  AOI211_X1 g218(.A(KEYINPUT93), .B(new_n404), .C1(new_n344), .C2(new_n335), .ZN(new_n405));
  INV_X1    g219(.A(new_n346), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G475), .B1(new_n407), .B2(G902), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n355), .A2(new_n400), .A3(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n299), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  NAND2_X1  g225(.A1(G234), .A2(G237), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(G952), .A3(new_n263), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n267), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n415), .A2(G902), .A3(new_n412), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT21), .B(G898), .Z(new_n418));
  OAI21_X1  g232(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G116), .B(G119), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT2), .B(G113), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n211), .A2(new_n423), .A3(new_n227), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n425));
  INV_X1    g239(.A(G119), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G116), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(G113), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n420), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n433), .A2(new_n421), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n209), .A2(new_n247), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n439));
  XOR2_X1   g253(.A(G110), .B(G122), .Z(new_n440));
  AND4_X1   g254(.A1(KEYINPUT87), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n440), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n424), .B2(new_n437), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT87), .B1(new_n443), .B2(new_n439), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n424), .A2(new_n437), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n424), .A2(new_n437), .A3(new_n448), .A4(new_n442), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(new_n439), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n244), .A2(G125), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(G125), .B2(new_n224), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n263), .A2(G224), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n455), .B(KEYINPUT88), .Z(new_n456));
  XOR2_X1   g270(.A(new_n454), .B(new_n456), .Z(new_n457));
  NAND3_X1  g271(.A1(new_n445), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G210), .B1(G237), .B2(G902), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n440), .B(KEYINPUT8), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n435), .B1(new_n434), .B2(new_n430), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n447), .B2(new_n449), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n454), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n458), .A2(new_n459), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n459), .B1(new_n458), .B2(new_n467), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n411), .B(new_n419), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n410), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n426), .A2(G128), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n240), .A2(G119), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT24), .B(G110), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n240), .A2(KEYINPUT23), .A3(G119), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n479), .A2(new_n473), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n477), .B1(new_n481), .B2(G110), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n309), .A2(new_n216), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n325), .A3(new_n483), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n484), .B(KEYINPUT70), .Z(new_n485));
  AND2_X1   g299(.A1(new_n481), .A2(G110), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  OR3_X1    g301(.A1(new_n343), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT22), .Z(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n233), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n492), .A3(new_n488), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n276), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(KEYINPUT71), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n389), .B1(G234), .B2(new_n276), .ZN(new_n501));
  INV_X1    g315(.A(new_n499), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(KEYINPUT72), .B2(KEYINPUT25), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n501), .C1(new_n496), .C2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n494), .A2(new_n495), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n501), .A2(G902), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n225), .A2(new_n255), .ZN(new_n510));
  INV_X1    g324(.A(new_n232), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n230), .A2(G137), .ZN(new_n512));
  OAI21_X1  g326(.A(G131), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n244), .A2(new_n238), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(KEYINPUT30), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n244), .A2(new_n238), .A3(new_n513), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n224), .A2(KEYINPUT65), .B1(new_n238), .B2(new_n236), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT65), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n215), .A2(new_n223), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n423), .B(new_n515), .C1(new_n520), .C2(KEYINPUT30), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n301), .A2(new_n522), .A3(G210), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n301), .B2(G210), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT26), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT26), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n526), .A2(new_n529), .A3(G101), .ZN(new_n530));
  AOI21_X1  g344(.A(G101), .B1(new_n526), .B2(new_n529), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n514), .B1(new_n239), .B2(new_n224), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n423), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n521), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT31), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT31), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n521), .A2(new_n532), .A3(new_n538), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n533), .A2(KEYINPUT67), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n510), .A2(new_n541), .A3(new_n514), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n540), .A2(new_n542), .A3(new_n422), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n255), .A3(new_n519), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n422), .B1(new_n547), .B2(new_n514), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT28), .B1(new_n548), .B2(new_n534), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n537), .B(new_n539), .C1(new_n550), .C2(new_n532), .ZN(new_n551));
  NOR2_X1   g365(.A1(G472), .A2(G902), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n551), .A2(KEYINPUT32), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT32), .B1(new_n551), .B2(new_n552), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n521), .A2(new_n535), .ZN(new_n556));
  INV_X1    g370(.A(new_n532), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n545), .A2(new_n549), .A3(new_n532), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT68), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n422), .B1(new_n510), .B2(new_n514), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT28), .B1(new_n534), .B2(new_n563), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n564), .A2(KEYINPUT69), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n545), .A2(KEYINPUT69), .A3(new_n564), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(KEYINPUT29), .A3(new_n532), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT68), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n558), .A2(new_n559), .A3(new_n569), .A4(new_n560), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n562), .A2(new_n568), .A3(new_n276), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G472), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n509), .B1(new_n555), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n472), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(new_n208), .ZN(G3));
  INV_X1    g390(.A(G472), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n551), .B2(new_n276), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT98), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT98), .B1(new_n551), .B2(new_n552), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n509), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n470), .A2(new_n299), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n355), .A2(new_n408), .ZN(new_n586));
  AND4_X1   g400(.A1(new_n398), .A2(new_n395), .A3(new_n276), .A4(new_n396), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n395), .A2(new_n588), .A3(new_n396), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT99), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n388), .B2(new_n391), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT99), .B(new_n390), .C1(new_n376), .C2(new_n387), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT33), .B(new_n394), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n589), .A2(new_n593), .A3(new_n276), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n587), .B1(new_n594), .B2(G478), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n586), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(new_n585), .A3(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT34), .B(G104), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G6));
  NAND2_X1  g415(.A1(new_n408), .A2(KEYINPUT102), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n603), .B(G475), .C1(new_n407), .C2(G902), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n400), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n354), .A2(KEYINPUT101), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n354), .A2(KEYINPUT101), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n349), .B(new_n353), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n584), .A2(new_n585), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NOR2_X1   g427(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(new_n489), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n507), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n504), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n580), .A2(new_n618), .A3(new_n582), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n410), .A2(new_n471), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT37), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G110), .ZN(G12));
  NAND2_X1  g436(.A1(new_n555), .A2(new_n572), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(new_n294), .A3(new_n298), .ZN(new_n624));
  OAI211_X1 g438(.A(new_n411), .B(new_n617), .C1(new_n468), .C2(new_n469), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n413), .B1(new_n416), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n606), .A2(new_n605), .A3(new_n609), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  XNOR2_X1  g446(.A(new_n628), .B(KEYINPUT39), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n299), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n617), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT40), .B1(new_n299), .B2(new_n633), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n556), .A2(new_n532), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n534), .A2(new_n563), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n557), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n639), .B2(new_n642), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(G902), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n555), .B1(new_n577), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n400), .B1(new_n355), .B2(new_n408), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n411), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n468), .A2(new_n469), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n458), .A2(new_n467), .ZN(new_n653));
  INV_X1    g467(.A(new_n459), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n458), .A2(new_n459), .A3(new_n467), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT38), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR3_X1    g471(.A1(new_n650), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT104), .B1(new_n638), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n658), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n660), .A2(new_n636), .A3(new_n661), .A4(new_n637), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n665));
  INV_X1    g479(.A(new_n411), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n655), .B2(new_n656), .ZN(new_n667));
  INV_X1    g481(.A(new_n298), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n282), .A2(KEYINPUT82), .A3(new_n283), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n290), .B1(new_n286), .B2(new_n289), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n276), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G469), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n668), .B1(new_n672), .B2(new_n280), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n667), .A2(new_n673), .A3(new_n623), .A4(new_n617), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n595), .B(KEYINPUT100), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n355), .A2(new_n408), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n676), .A3(new_n629), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n665), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n626), .A2(KEYINPUT105), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  NAND2_X1  g496(.A1(new_n275), .A2(new_n276), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n280), .A3(new_n297), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n471), .A2(new_n573), .A3(new_n598), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT106), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n471), .A2(new_n610), .A3(new_n573), .A4(new_n686), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NAND4_X1  g506(.A1(new_n355), .A2(new_n419), .A3(new_n400), .A4(new_n408), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n555), .B2(new_n572), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n667), .A3(new_n617), .A4(new_n686), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT107), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  AND2_X1   g511(.A1(new_n504), .A2(new_n508), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n537), .B(new_n539), .C1(new_n567), .C2(new_n532), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n552), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n579), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n685), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n471), .A2(new_n702), .A3(new_n649), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NOR2_X1   g518(.A1(new_n625), .A2(new_n685), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n617), .A2(new_n579), .A3(new_n700), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n677), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NAND2_X1  g523(.A1(G469), .A2(G902), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT108), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n286), .B2(new_n289), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT108), .B1(new_n274), .B2(new_n270), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n712), .A2(new_n713), .A3(new_n293), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n710), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT108), .B1(new_n282), .B2(new_n283), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n289), .A2(new_n711), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n715), .A3(G469), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n280), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n655), .A2(new_n411), .A3(new_n656), .ZN(new_n722));
  INV_X1    g536(.A(new_n297), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(KEYINPUT42), .A3(new_n573), .A4(new_n679), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n468), .A2(new_n469), .A3(new_n666), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n717), .A2(G469), .A3(new_n718), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT109), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n280), .A3(new_n719), .A4(new_n710), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n573), .A3(new_n297), .A4(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n726), .B1(new_n731), .B2(new_n677), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT110), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n237), .ZN(G33));
  INV_X1    g549(.A(new_n630), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n731), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n230), .ZN(G36));
  INV_X1    g552(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n586), .A2(new_n675), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n586), .A2(KEYINPUT43), .A3(new_n675), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT112), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT112), .B1(new_n742), .B2(new_n743), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n583), .A2(new_n617), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n739), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n722), .B1(new_n749), .B2(KEYINPUT44), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n669), .B2(new_n670), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n718), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(G469), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n710), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n710), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n280), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n633), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n297), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n748), .A2(new_n750), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  INV_X1    g579(.A(new_n759), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT47), .B1(new_n766), .B2(new_n723), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n722), .A2(new_n698), .A3(new_n623), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n759), .A2(new_n769), .A3(new_n297), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n767), .A2(new_n679), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  AOI21_X1  g586(.A(new_n414), .B1(new_n742), .B2(new_n743), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n722), .A2(new_n685), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n574), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT48), .Z(new_n777));
  NOR2_X1   g591(.A1(new_n648), .A2(new_n414), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n698), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT116), .Z(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n598), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(G952), .A3(new_n263), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n701), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n773), .A2(new_n686), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n652), .A2(new_n657), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n666), .A3(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(KEYINPUT50), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n775), .A2(new_n706), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n773), .A2(new_n783), .A3(new_n727), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT114), .Z(new_n793));
  NAND2_X1  g607(.A1(new_n767), .A2(new_n770), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n684), .A2(new_n280), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n298), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n780), .A2(new_n586), .A3(new_n597), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n790), .A2(new_n791), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AND4_X1   g620(.A1(new_n800), .A2(new_n789), .A3(new_n788), .A4(new_n801), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(KEYINPUT117), .A3(new_n803), .A4(new_n791), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n782), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n784), .A2(new_n667), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n630), .A2(new_n626), .B1(new_n705), .B2(new_n707), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n667), .A2(new_n649), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n297), .A2(new_n648), .A3(new_n618), .A4(new_n629), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n730), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT105), .B1(new_n626), .B2(new_n679), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n624), .A2(new_n625), .A3(new_n677), .A4(new_n665), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n811), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n681), .A2(KEYINPUT52), .A3(new_n811), .A4(new_n814), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n737), .B1(new_n725), .B2(new_n732), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT113), .B(new_n409), .C1(new_n586), .C2(new_n675), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n586), .B2(new_n597), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n584), .A3(new_n585), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n410), .B(new_n471), .C1(new_n573), .C2(new_n619), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n687), .A2(new_n691), .A3(new_n695), .A4(new_n703), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n400), .A2(new_n605), .A3(new_n617), .A4(new_n629), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n609), .A3(new_n727), .ZN(new_n832));
  INV_X1    g646(.A(new_n624), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n832), .A2(new_n833), .B1(new_n707), .B2(new_n724), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n822), .A2(new_n829), .A3(new_n830), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n821), .A2(new_n835), .A3(KEYINPUT53), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n821), .B2(new_n835), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n821), .A2(new_n835), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n821), .A2(new_n835), .A3(KEYINPUT53), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n809), .A2(new_n810), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(G952), .B2(G953), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n848), .A2(new_n849), .A3(new_n509), .A4(new_n666), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n740), .A2(new_n648), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n786), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n847), .B1(new_n668), .B2(new_n852), .ZN(G75));
  AOI21_X1  g667(.A(new_n276), .B1(new_n841), .B2(new_n843), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(G210), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT56), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n445), .A2(new_n452), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(new_n457), .Z(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT55), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n855), .B2(new_n856), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n267), .A2(G952), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G51));
  NAND3_X1  g677(.A1(new_n838), .A2(new_n844), .A3(KEYINPUT118), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n841), .A2(new_n843), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT54), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n710), .B(KEYINPUT57), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n275), .ZN(new_n870));
  INV_X1    g684(.A(new_n754), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n854), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n874));
  INV_X1    g688(.A(new_n862), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n872), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n869), .B2(new_n275), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT119), .B1(new_n878), .B2(new_n862), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(G54));
  NAND3_X1  g694(.A1(KEYINPUT120), .A2(KEYINPUT58), .A3(G475), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n854), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT120), .B1(KEYINPUT58), .B2(G475), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n350), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n862), .ZN(G60));
  NAND2_X1  g702(.A1(new_n589), .A2(new_n593), .ZN(new_n889));
  NAND2_X1  g703(.A1(G478), .A2(G902), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT59), .Z(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n845), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n889), .A2(new_n891), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n864), .A2(new_n867), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n875), .A3(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT122), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT60), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n865), .A2(new_n615), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n865), .A2(new_n898), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n875), .B(new_n899), .C1(new_n900), .C2(new_n505), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT61), .ZN(G66));
  AND2_X1   g717(.A1(new_n829), .A2(new_n830), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n418), .A2(G224), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n904), .A2(new_n415), .B1(new_n263), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(G898), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n857), .B1(new_n907), .B2(new_n415), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n906), .B(new_n908), .Z(G69));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n910));
  INV_X1    g724(.A(new_n663), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n681), .A2(new_n811), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n681), .A2(KEYINPUT123), .A3(new_n811), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n663), .A2(KEYINPUT62), .A3(new_n914), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n515), .B1(new_n520), .B2(KEYINPUT30), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n319), .A2(new_n320), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n920), .B(new_n921), .Z(new_n922));
  AND2_X1   g736(.A1(new_n764), .A2(new_n771), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n826), .A2(new_n573), .A3(new_n634), .A4(new_n727), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n922), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n748), .A2(new_n750), .A3(new_n763), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n764), .A2(KEYINPUT124), .A3(new_n914), .A4(new_n915), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n771), .A2(new_n822), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n763), .A2(new_n573), .A3(new_n812), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n930), .A2(new_n931), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n267), .B(new_n925), .C1(new_n936), .C2(new_n922), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n922), .A2(new_n627), .A3(new_n267), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n937), .A2(new_n939), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n928), .A2(new_n929), .B1(new_n934), .B2(new_n933), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n922), .B1(new_n943), .B2(new_n931), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n925), .A2(new_n267), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n942), .A2(new_n947), .ZN(G72));
  NAND4_X1  g762(.A1(new_n919), .A2(new_n904), .A3(new_n923), .A4(new_n924), .ZN(new_n949));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n640), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n558), .A2(new_n536), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n865), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n875), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n930), .A2(new_n904), .A3(new_n931), .A4(new_n935), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n532), .B(new_n556), .C1(new_n957), .C2(new_n951), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n951), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n535), .A3(new_n557), .A4(new_n521), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n862), .B1(new_n952), .B2(new_n640), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n955), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(G57));
endmodule


