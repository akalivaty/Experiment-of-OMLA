

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n485, n486, n487, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803;

  INV_X1 U368 ( .A(n696), .ZN(n347) );
  INV_X1 U369 ( .A(G902), .ZN(n438) );
  XNOR2_X1 U370 ( .A(G116), .B(KEYINPUT106), .ZN(n562) );
  XNOR2_X1 U371 ( .A(G104), .B(G140), .ZN(n511) );
  NOR2_X1 U372 ( .A1(G953), .A2(G237), .ZN(n574) );
  XOR2_X2 U373 ( .A(n688), .B(KEYINPUT59), .Z(n486) );
  AND2_X2 U374 ( .A1(n407), .A2(n417), .ZN(n406) );
  XNOR2_X1 U375 ( .A(n348), .B(n347), .ZN(G57) );
  NAND2_X1 U376 ( .A1(n695), .A2(n350), .ZN(n348) );
  XOR2_X2 U377 ( .A(n693), .B(n692), .Z(n483) );
  BUF_X1 U378 ( .A(n770), .Z(n349) );
  INV_X1 U379 ( .A(G237), .ZN(n505) );
  XOR2_X1 U380 ( .A(KEYINPUT103), .B(G143), .Z(n580) );
  BUF_X1 U381 ( .A(n794), .Z(n354) );
  XNOR2_X2 U382 ( .A(n362), .B(n395), .ZN(n593) );
  BUF_X2 U383 ( .A(n398), .Z(n774) );
  INV_X1 U384 ( .A(n654), .ZN(n445) );
  XNOR2_X1 U385 ( .A(n573), .B(n572), .ZN(n616) );
  INV_X4 U386 ( .A(G953), .ZN(n794) );
  XNOR2_X1 U387 ( .A(n390), .B(n643), .ZN(n698) );
  NAND2_X1 U388 ( .A1(n705), .A2(n683), .ZN(n393) );
  XNOR2_X1 U389 ( .A(n619), .B(n618), .ZN(n743) );
  XNOR2_X1 U390 ( .A(n627), .B(KEYINPUT117), .ZN(n603) );
  OR2_X1 U391 ( .A1(n614), .A2(n472), .ZN(n750) );
  AND2_X2 U392 ( .A1(n616), .A2(n587), .ZN(n716) );
  INV_X1 U393 ( .A(G125), .ZN(n367) );
  INV_X1 U394 ( .A(KEYINPUT17), .ZN(n368) );
  INV_X1 U395 ( .A(KEYINPUT56), .ZN(n357) );
  INV_X1 U396 ( .A(KEYINPUT60), .ZN(n355) );
  INV_X1 U397 ( .A(n698), .ZN(n353) );
  INV_X1 U398 ( .A(n393), .ZN(n352) );
  XNOR2_X1 U399 ( .A(n411), .B(n648), .ZN(n705) );
  NAND2_X1 U400 ( .A1(n391), .A2(n374), .ZN(n411) );
  XNOR2_X1 U401 ( .A(n656), .B(n655), .ZN(n719) );
  NOR2_X1 U402 ( .A1(n445), .A2(n444), .ZN(n443) );
  AND2_X1 U403 ( .A1(n366), .A2(n590), .ZN(n365) );
  NAND2_X1 U404 ( .A1(n361), .A2(n439), .ZN(n436) );
  XNOR2_X1 U405 ( .A(n412), .B(n585), .ZN(n587) );
  XNOR2_X1 U406 ( .A(n582), .B(n413), .ZN(n688) );
  XNOR2_X1 U407 ( .A(n583), .B(n581), .ZN(n413) );
  XNOR2_X1 U408 ( .A(n792), .B(n490), .ZN(n459) );
  XNOR2_X1 U409 ( .A(n415), .B(n414), .ZN(n577) );
  NAND2_X1 U410 ( .A1(n507), .A2(G214), .ZN(n745) );
  XNOR2_X1 U411 ( .A(n489), .B(G146), .ZN(n792) );
  INV_X1 U412 ( .A(n777), .ZN(n350) );
  XNOR2_X2 U413 ( .A(KEYINPUT79), .B(G110), .ZN(n497) );
  XNOR2_X2 U414 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n534) );
  XNOR2_X2 U415 ( .A(G140), .B(KEYINPUT10), .ZN(n537) );
  XNOR2_X2 U416 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n489) );
  XNOR2_X2 U417 ( .A(G119), .B(G116), .ZN(n500) );
  XOR2_X1 U418 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n563) );
  XNOR2_X2 U419 ( .A(G104), .B(G122), .ZN(n575) );
  XOR2_X1 U420 ( .A(KEYINPUT99), .B(KEYINPUT78), .Z(n516) );
  XNOR2_X1 U421 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n498) );
  XNOR2_X2 U422 ( .A(G122), .B(G107), .ZN(n561) );
  XNOR2_X1 U423 ( .A(KEYINPUT81), .B(KEYINPUT24), .ZN(n530) );
  XNOR2_X1 U424 ( .A(n504), .B(n784), .ZN(n700) );
  NAND2_X1 U425 ( .A1(n351), .A2(KEYINPUT44), .ZN(n466) );
  NAND2_X1 U426 ( .A1(n353), .A2(n352), .ZN(n351) );
  XNOR2_X1 U427 ( .A(n356), .B(n355), .ZN(G60) );
  NAND2_X1 U428 ( .A1(n690), .A2(n350), .ZN(n356) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(G51) );
  NAND2_X1 U430 ( .A1(n359), .A2(n350), .ZN(n358) );
  NAND2_X1 U431 ( .A1(n423), .A2(n612), .ZN(n658) );
  XNOR2_X2 U432 ( .A(n401), .B(n515), .ZN(n612) );
  XNOR2_X1 U433 ( .A(n702), .B(n360), .ZN(n359) );
  INV_X1 U434 ( .A(n701), .ZN(n360) );
  NAND2_X1 U435 ( .A1(n691), .A2(n526), .ZN(n361) );
  XNOR2_X2 U436 ( .A(n525), .B(n524), .ZN(n691) );
  XNOR2_X2 U437 ( .A(n789), .B(n459), .ZN(n525) );
  NOR2_X2 U438 ( .A1(n770), .A2(G902), .ZN(n401) );
  NAND2_X1 U439 ( .A1(n593), .A2(n746), .ZN(n610) );
  NAND2_X1 U440 ( .A1(n365), .A2(n363), .ZN(n362) );
  XNOR2_X1 U441 ( .A(n364), .B(n396), .ZN(n363) );
  NAND2_X1 U442 ( .A1(n381), .A2(n745), .ZN(n364) );
  XNOR2_X1 U443 ( .A(n658), .B(n588), .ZN(n366) );
  NAND2_X1 U444 ( .A1(G125), .A2(n368), .ZN(n369) );
  NAND2_X1 U445 ( .A1(n367), .A2(KEYINPUT17), .ZN(n370) );
  NAND2_X1 U446 ( .A1(n369), .A2(n370), .ZN(n493) );
  BUF_X1 U447 ( .A(n569), .Z(n371) );
  NAND2_X1 U448 ( .A1(n410), .A2(n726), .ZN(n372) );
  NAND2_X1 U449 ( .A1(n410), .A2(n726), .ZN(n676) );
  XNOR2_X1 U450 ( .A(n700), .B(n699), .ZN(n701) );
  XNOR2_X1 U451 ( .A(n394), .B(n459), .ZN(n504) );
  NOR2_X1 U452 ( .A1(n461), .A2(KEYINPUT34), .ZN(n389) );
  NAND2_X1 U453 ( .A1(n420), .A2(n418), .ZN(n417) );
  NAND2_X1 U454 ( .A1(n674), .A2(n419), .ZN(n418) );
  NAND2_X1 U455 ( .A1(n421), .A2(KEYINPUT66), .ZN(n420) );
  NAND2_X1 U456 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n419) );
  XNOR2_X1 U457 ( .A(G137), .B(G131), .ZN(n508) );
  XNOR2_X1 U458 ( .A(G113), .B(KEYINPUT74), .ZN(n501) );
  INV_X1 U459 ( .A(KEYINPUT30), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n599), .B(KEYINPUT111), .ZN(n381) );
  XNOR2_X1 U461 ( .A(KEYINPUT68), .B(G101), .ZN(n490) );
  XNOR2_X1 U462 ( .A(KEYINPUT93), .B(KEYINPUT18), .ZN(n494) );
  XNOR2_X1 U463 ( .A(n635), .B(n634), .ZN(n760) );
  NAND2_X1 U464 ( .A1(n685), .A2(n458), .ZN(n455) );
  INV_X1 U465 ( .A(n760), .ZN(n388) );
  NOR2_X1 U466 ( .A1(n386), .A2(n385), .ZN(n384) );
  AND2_X1 U467 ( .A1(n760), .A2(KEYINPUT34), .ZN(n385) );
  NAND2_X1 U468 ( .A1(n382), .A2(n387), .ZN(n386) );
  INV_X1 U469 ( .A(n642), .ZN(n387) );
  INV_X1 U470 ( .A(KEYINPUT0), .ZN(n462) );
  NAND2_X1 U471 ( .A1(n427), .A2(n426), .ZN(n596) );
  INV_X1 U472 ( .A(n674), .ZN(n421) );
  NAND2_X1 U473 ( .A1(n478), .A2(n477), .ZN(n476) );
  INV_X1 U474 ( .A(KEYINPUT89), .ZN(n477) );
  INV_X1 U475 ( .A(n802), .ZN(n478) );
  AND2_X1 U476 ( .A1(n802), .A2(KEYINPUT89), .ZN(n480) );
  INV_X1 U477 ( .A(KEYINPUT19), .ZN(n468) );
  NAND2_X1 U478 ( .A1(n472), .A2(KEYINPUT19), .ZN(n471) );
  NAND2_X1 U479 ( .A1(n526), .A2(G902), .ZN(n439) );
  NAND2_X1 U480 ( .A1(G472), .A2(n438), .ZN(n437) );
  XNOR2_X1 U481 ( .A(KEYINPUT98), .B(KEYINPUT100), .ZN(n519) );
  XOR2_X1 U482 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n517) );
  INV_X1 U483 ( .A(KEYINPUT92), .ZN(n392) );
  XNOR2_X1 U484 ( .A(G110), .B(G128), .ZN(n527) );
  XNOR2_X1 U485 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U486 ( .A(n425), .ZN(n531) );
  XNOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n425) );
  NAND2_X1 U488 ( .A1(n406), .A2(n404), .ZN(n410) );
  NAND2_X1 U489 ( .A1(n405), .A2(n380), .ZN(n404) );
  NAND2_X1 U490 ( .A1(G234), .A2(G237), .ZN(n547) );
  NAND2_X1 U491 ( .A1(n461), .A2(KEYINPUT34), .ZN(n382) );
  INV_X1 U492 ( .A(KEYINPUT1), .ZN(n424) );
  OR2_X2 U493 ( .A1(n436), .A2(n435), .ZN(n599) );
  XNOR2_X1 U494 ( .A(n416), .B(G113), .ZN(n415) );
  INV_X1 U495 ( .A(KEYINPUT104), .ZN(n416) );
  XNOR2_X1 U496 ( .A(G131), .B(KEYINPUT12), .ZN(n414) );
  XOR2_X1 U497 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n579) );
  AND2_X1 U498 ( .A1(n602), .A2(KEYINPUT36), .ZN(n444) );
  NAND2_X1 U499 ( .A1(n448), .A2(n604), .ZN(n447) );
  INV_X1 U500 ( .A(KEYINPUT80), .ZN(n395) );
  NAND2_X1 U501 ( .A1(n688), .A2(n438), .ZN(n412) );
  XNOR2_X1 U502 ( .A(n496), .B(n403), .ZN(n394) );
  NAND2_X1 U503 ( .A1(n454), .A2(n453), .ZN(n451) );
  AND2_X1 U504 ( .A1(n457), .A2(n373), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n384), .A2(n383), .ZN(n390) );
  NAND2_X1 U506 ( .A1(n388), .A2(n389), .ZN(n383) );
  INV_X1 U507 ( .A(n739), .ZN(n460) );
  XNOR2_X1 U508 ( .A(n776), .B(n429), .ZN(n428) );
  INV_X1 U509 ( .A(n745), .ZN(n472) );
  XOR2_X1 U510 ( .A(n611), .B(KEYINPUT40), .Z(n373) );
  XNOR2_X1 U511 ( .A(n612), .B(n424), .ZN(n729) );
  NOR2_X1 U512 ( .A1(n646), .A2(n645), .ZN(n374) );
  AND2_X1 U513 ( .A1(n687), .A2(n476), .ZN(n375) );
  INV_X1 U514 ( .A(n685), .ZN(n457) );
  NOR2_X1 U515 ( .A1(n747), .A2(n733), .ZN(n376) );
  AND2_X1 U516 ( .A1(n667), .A2(n706), .ZN(n377) );
  AND2_X1 U517 ( .A1(n745), .A2(n468), .ZN(n378) );
  INV_X1 U518 ( .A(n373), .ZN(n458) );
  XNOR2_X1 U519 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n379) );
  INV_X1 U520 ( .A(KEYINPUT111), .ZN(n450) );
  AND2_X1 U521 ( .A1(n674), .A2(KEYINPUT66), .ZN(n380) );
  INV_X1 U522 ( .A(n391), .ZN(n652) );
  XNOR2_X2 U523 ( .A(n644), .B(n379), .ZN(n391) );
  NAND2_X1 U524 ( .A1(n391), .A2(n666), .ZN(n706) );
  XNOR2_X1 U525 ( .A(n393), .B(n392), .ZN(n669) );
  INV_X1 U526 ( .A(n427), .ZN(n684) );
  XNOR2_X2 U527 ( .A(n397), .B(KEYINPUT83), .ZN(n427) );
  NAND2_X2 U528 ( .A1(n613), .A2(n560), .ZN(n397) );
  XNOR2_X2 U529 ( .A(n559), .B(n558), .ZN(n613) );
  XNOR2_X1 U530 ( .A(n372), .B(KEYINPUT65), .ZN(n398) );
  XNOR2_X1 U531 ( .A(n676), .B(KEYINPUT65), .ZN(n767) );
  INV_X1 U532 ( .A(n469), .ZN(n399) );
  XNOR2_X1 U533 ( .A(n431), .B(KEYINPUT71), .ZN(n430) );
  OR2_X2 U534 ( .A1(n436), .A2(n435), .ZN(n400) );
  INV_X1 U535 ( .A(n728), .ZN(n423) );
  XNOR2_X1 U536 ( .A(n536), .B(n485), .ZN(n538) );
  XNOR2_X1 U537 ( .A(n533), .B(n532), .ZN(n536) );
  XNOR2_X1 U538 ( .A(n599), .B(n450), .ZN(n649) );
  BUF_X1 U539 ( .A(n775), .Z(n402) );
  XNOR2_X1 U540 ( .A(n538), .B(n583), .ZN(n775) );
  INV_X1 U541 ( .A(n402), .ZN(n429) );
  BUF_X1 U542 ( .A(n449), .Z(n403) );
  NAND2_X1 U543 ( .A1(n672), .A2(n422), .ZN(n407) );
  XNOR2_X1 U544 ( .A(n409), .B(KEYINPUT87), .ZN(n408) );
  INV_X1 U545 ( .A(n672), .ZN(n405) );
  NAND2_X1 U546 ( .A1(n408), .A2(n778), .ZN(n726) );
  NAND2_X1 U547 ( .A1(n722), .A2(KEYINPUT2), .ZN(n409) );
  AND2_X1 U548 ( .A1(n671), .A2(n675), .ZN(n422) );
  XNOR2_X1 U549 ( .A(n595), .B(KEYINPUT85), .ZN(n432) );
  NAND2_X1 U550 ( .A1(n432), .A2(n607), .ZN(n431) );
  NAND2_X1 U551 ( .A1(n703), .A2(n623), .ZN(n434) );
  XNOR2_X1 U552 ( .A(n434), .B(n624), .ZN(n433) );
  XNOR2_X1 U553 ( .A(n440), .B(n625), .ZN(n482) );
  NAND2_X1 U554 ( .A1(n722), .A2(n778), .ZN(n672) );
  NOR2_X2 U555 ( .A1(n475), .A2(n481), .ZN(n722) );
  INV_X1 U556 ( .A(n487), .ZN(n426) );
  NAND2_X1 U557 ( .A1(n466), .A2(n377), .ZN(n465) );
  NAND2_X1 U558 ( .A1(n482), .A2(n480), .ZN(n479) );
  XNOR2_X1 U559 ( .A(n465), .B(KEYINPUT91), .ZN(n464) );
  NOR2_X1 U560 ( .A1(n428), .A2(n777), .ZN(G66) );
  NAND2_X1 U561 ( .A1(n433), .A2(n430), .ZN(n440) );
  NAND2_X1 U562 ( .A1(n452), .A2(n451), .ZN(n703) );
  NOR2_X1 U563 ( .A1(n691), .A2(n437), .ZN(n435) );
  NOR2_X1 U564 ( .A1(n400), .A2(n728), .ZN(n653) );
  XNOR2_X2 U565 ( .A(n400), .B(KEYINPUT6), .ZN(n664) );
  NAND2_X2 U566 ( .A1(n442), .A2(n441), .ZN(n682) );
  NAND2_X1 U567 ( .A1(n603), .A2(KEYINPUT36), .ZN(n441) );
  AND2_X2 U568 ( .A1(n446), .A2(n443), .ZN(n442) );
  OR2_X2 U569 ( .A1(n603), .A2(n447), .ZN(n446) );
  INV_X1 U570 ( .A(n602), .ZN(n448) );
  XNOR2_X1 U571 ( .A(n682), .B(KEYINPUT90), .ZN(n605) );
  XNOR2_X2 U572 ( .A(n449), .B(G134), .ZN(n569) );
  XNOR2_X2 U573 ( .A(n491), .B(G128), .ZN(n449) );
  INV_X1 U574 ( .A(n400), .ZN(n657) );
  NAND2_X1 U575 ( .A1(n632), .A2(n458), .ZN(n456) );
  XNOR2_X2 U576 ( .A(n610), .B(n609), .ZN(n632) );
  INV_X1 U577 ( .A(n632), .ZN(n454) );
  AND2_X1 U578 ( .A1(n456), .A2(n455), .ZN(n452) );
  AND2_X1 U579 ( .A1(n660), .A2(n460), .ZN(n656) );
  INV_X1 U580 ( .A(n660), .ZN(n461) );
  XNOR2_X2 U581 ( .A(n641), .B(n462), .ZN(n660) );
  XNOR2_X2 U582 ( .A(n463), .B(KEYINPUT45), .ZN(n778) );
  NAND2_X1 U583 ( .A1(n464), .A2(n670), .ZN(n463) );
  NAND2_X1 U584 ( .A1(n469), .A2(n745), .ZN(n602) );
  NAND2_X1 U585 ( .A1(n470), .A2(n467), .ZN(n640) );
  NAND2_X1 U586 ( .A1(n469), .A2(n378), .ZN(n467) );
  INV_X1 U587 ( .A(n591), .ZN(n469) );
  AND2_X1 U588 ( .A1(n473), .A2(n471), .ZN(n470) );
  NAND2_X1 U589 ( .A1(n591), .A2(KEYINPUT19), .ZN(n473) );
  XNOR2_X2 U590 ( .A(n474), .B(n506), .ZN(n591) );
  NAND2_X1 U591 ( .A1(n700), .A2(n673), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n479), .A2(n375), .ZN(n475) );
  NOR2_X1 U593 ( .A1(n482), .A2(KEYINPUT89), .ZN(n481) );
  XNOR2_X2 U594 ( .A(n569), .B(n509), .ZN(n789) );
  XNOR2_X1 U595 ( .A(n678), .B(n677), .ZN(n680) );
  XNOR2_X2 U596 ( .A(n543), .B(n542), .ZN(n732) );
  AND2_X1 U597 ( .A1(n680), .A2(n350), .ZN(G63) );
  AND2_X1 U598 ( .A1(G221), .A2(n566), .ZN(n485) );
  NOR2_X1 U599 ( .A1(n718), .A2(n716), .ZN(n487) );
  AND2_X1 U600 ( .A1(n679), .A2(G953), .ZN(n777) );
  INV_X1 U601 ( .A(KEYINPUT46), .ZN(n624) );
  NOR2_X1 U602 ( .A1(n729), .A2(n728), .ZN(n633) );
  BUF_X1 U603 ( .A(n703), .Z(n704) );
  XNOR2_X2 U604 ( .A(G143), .B(KEYINPUT84), .ZN(n491) );
  NAND2_X1 U605 ( .A1(G224), .A2(n794), .ZN(n492) );
  XNOR2_X1 U606 ( .A(n493), .B(n492), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n497), .B(G107), .ZN(n513) );
  XNOR2_X1 U609 ( .A(n575), .B(n498), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n513), .B(n499), .ZN(n503) );
  XNOR2_X1 U611 ( .A(n500), .B(KEYINPUT3), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n502), .B(n501), .ZN(n522) );
  XNOR2_X1 U613 ( .A(n503), .B(n522), .ZN(n784) );
  XNOR2_X1 U614 ( .A(G902), .B(KEYINPUT15), .ZN(n673) );
  NAND2_X1 U615 ( .A1(n438), .A2(n505), .ZN(n507) );
  NAND2_X1 U616 ( .A1(n507), .A2(G210), .ZN(n506) );
  XNOR2_X1 U617 ( .A(n508), .B(KEYINPUT70), .ZN(n509) );
  NAND2_X1 U618 ( .A1(n354), .A2(G227), .ZN(n510) );
  XNOR2_X1 U619 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U620 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U621 ( .A(n525), .B(n514), .ZN(n770) );
  XNOR2_X1 U622 ( .A(KEYINPUT73), .B(G469), .ZN(n515) );
  AND2_X1 U623 ( .A1(n612), .A2(n640), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n517), .B(n516), .ZN(n521) );
  NAND2_X1 U625 ( .A1(n574), .A2(G210), .ZN(n518) );
  XNOR2_X1 U626 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n521), .B(n520), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n523), .B(n522), .ZN(n524) );
  INV_X1 U629 ( .A(G472), .ZN(n526) );
  INV_X1 U630 ( .A(n527), .ZN(n529) );
  XNOR2_X1 U631 ( .A(G119), .B(G137), .ZN(n528) );
  XNOR2_X1 U632 ( .A(n529), .B(n528), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n794), .A2(G234), .ZN(n535) );
  XNOR2_X1 U634 ( .A(n535), .B(n534), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n537), .B(G125), .ZN(n791) );
  XNOR2_X1 U636 ( .A(n791), .B(G146), .ZN(n583) );
  NAND2_X1 U637 ( .A1(n775), .A2(n438), .ZN(n543) );
  NAND2_X1 U638 ( .A1(G234), .A2(n673), .ZN(n539) );
  XNOR2_X1 U639 ( .A(KEYINPUT20), .B(n539), .ZN(n544) );
  NAND2_X1 U640 ( .A1(G217), .A2(n544), .ZN(n540) );
  XNOR2_X1 U641 ( .A(KEYINPUT96), .B(n540), .ZN(n541) );
  XNOR2_X1 U642 ( .A(n541), .B(KEYINPUT25), .ZN(n542) );
  AND2_X1 U643 ( .A1(n544), .A2(G221), .ZN(n546) );
  INV_X1 U644 ( .A(KEYINPUT21), .ZN(n545) );
  XNOR2_X1 U645 ( .A(n546), .B(n545), .ZN(n733) );
  XNOR2_X1 U646 ( .A(n547), .B(KEYINPUT14), .ZN(n552) );
  NAND2_X1 U647 ( .A1(G902), .A2(n552), .ZN(n548) );
  XOR2_X1 U648 ( .A(KEYINPUT94), .B(n548), .Z(n549) );
  NAND2_X1 U649 ( .A1(G953), .A2(n549), .ZN(n636) );
  NOR2_X1 U650 ( .A1(G900), .A2(n636), .ZN(n551) );
  INV_X1 U651 ( .A(KEYINPUT112), .ZN(n550) );
  XNOR2_X1 U652 ( .A(n551), .B(n550), .ZN(n553) );
  NAND2_X1 U653 ( .A1(G952), .A2(n552), .ZN(n758) );
  OR2_X1 U654 ( .A1(n758), .A2(G953), .ZN(n637) );
  AND2_X1 U655 ( .A1(n553), .A2(n637), .ZN(n589) );
  NOR2_X1 U656 ( .A1(n733), .A2(n589), .ZN(n554) );
  NAND2_X1 U657 ( .A1(n732), .A2(n554), .ZN(n556) );
  INV_X1 U658 ( .A(KEYINPUT72), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n600) );
  INV_X1 U660 ( .A(n600), .ZN(n557) );
  OR2_X2 U661 ( .A1(n649), .A2(n557), .ZN(n559) );
  INV_X1 U662 ( .A(KEYINPUT28), .ZN(n558) );
  XNOR2_X1 U663 ( .A(n561), .B(KEYINPUT9), .ZN(n565) );
  XNOR2_X1 U664 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U665 ( .A(n565), .B(n564), .Z(n568) );
  NAND2_X1 U666 ( .A1(G217), .A2(n566), .ZN(n567) );
  XNOR2_X1 U667 ( .A(n568), .B(n567), .ZN(n570) );
  XNOR2_X1 U668 ( .A(n371), .B(n570), .ZN(n677) );
  NAND2_X1 U669 ( .A1(n677), .A2(n438), .ZN(n573) );
  INV_X1 U670 ( .A(KEYINPUT108), .ZN(n571) );
  XNOR2_X1 U671 ( .A(n571), .B(G478), .ZN(n572) );
  INV_X1 U672 ( .A(n616), .ZN(n586) );
  NAND2_X1 U673 ( .A1(G214), .A2(n574), .ZN(n576) );
  XNOR2_X1 U674 ( .A(n576), .B(n575), .ZN(n578) );
  XNOR2_X1 U675 ( .A(n578), .B(n577), .ZN(n582) );
  XNOR2_X1 U676 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U677 ( .A(KEYINPUT13), .B(G475), .ZN(n584) );
  XNOR2_X1 U678 ( .A(n584), .B(KEYINPUT105), .ZN(n585) );
  INV_X1 U679 ( .A(n587), .ZN(n615) );
  AND2_X1 U680 ( .A1(n586), .A2(n615), .ZN(n718) );
  NAND2_X1 U681 ( .A1(n596), .A2(KEYINPUT47), .ZN(n594) );
  OR2_X2 U682 ( .A1(n732), .A2(n733), .ZN(n728) );
  INV_X1 U683 ( .A(KEYINPUT114), .ZN(n588) );
  INV_X1 U684 ( .A(n589), .ZN(n590) );
  OR2_X1 U685 ( .A1(n615), .A2(n616), .ZN(n642) );
  NOR2_X1 U686 ( .A1(n399), .A2(n642), .ZN(n592) );
  NAND2_X1 U687 ( .A1(n593), .A2(n592), .ZN(n697) );
  NAND2_X1 U688 ( .A1(n594), .A2(n697), .ZN(n595) );
  INV_X1 U689 ( .A(n596), .ZN(n598) );
  INV_X1 U690 ( .A(KEYINPUT47), .ZN(n597) );
  NAND2_X1 U691 ( .A1(n598), .A2(n597), .ZN(n606) );
  AND2_X1 U692 ( .A1(n600), .A2(n716), .ZN(n601) );
  AND2_X2 U693 ( .A1(n664), .A2(n601), .ZN(n627) );
  INV_X1 U694 ( .A(KEYINPUT36), .ZN(n604) );
  AND2_X1 U695 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U696 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n608) );
  XNOR2_X1 U697 ( .A(n591), .B(n608), .ZN(n614) );
  INV_X1 U698 ( .A(n614), .ZN(n746) );
  INV_X1 U699 ( .A(KEYINPUT39), .ZN(n609) );
  INV_X1 U700 ( .A(n716), .ZN(n685) );
  INV_X1 U701 ( .A(KEYINPUT115), .ZN(n611) );
  AND2_X1 U702 ( .A1(n612), .A2(n613), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U704 ( .A(n617), .B(KEYINPUT110), .ZN(n747) );
  OR2_X1 U705 ( .A1(n750), .A2(n747), .ZN(n619) );
  XNOR2_X1 U706 ( .A(KEYINPUT116), .B(KEYINPUT41), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n620), .A2(n743), .ZN(n622) );
  INV_X1 U708 ( .A(KEYINPUT42), .ZN(n621) );
  XNOR2_X1 U709 ( .A(n622), .B(n621), .ZN(n803) );
  INV_X1 U710 ( .A(n803), .ZN(n623) );
  INV_X1 U711 ( .A(KEYINPUT48), .ZN(n625) );
  AND2_X1 U712 ( .A1(n729), .A2(n745), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U714 ( .A(n628), .B(KEYINPUT43), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n629), .A2(n399), .ZN(n631) );
  INV_X1 U716 ( .A(KEYINPUT113), .ZN(n630) );
  XNOR2_X1 U717 ( .A(n631), .B(n630), .ZN(n802) );
  INV_X1 U718 ( .A(n718), .ZN(n712) );
  OR2_X1 U719 ( .A1(n632), .A2(n712), .ZN(n687) );
  NAND2_X1 U720 ( .A1(n633), .A2(n664), .ZN(n635) );
  INV_X1 U721 ( .A(KEYINPUT33), .ZN(n634) );
  OR2_X1 U722 ( .A1(n636), .A2(G898), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U725 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n660), .A2(n376), .ZN(n644) );
  XNOR2_X1 U727 ( .A(n664), .B(KEYINPUT82), .ZN(n646) );
  INV_X1 U728 ( .A(n732), .ZN(n663) );
  OR2_X1 U729 ( .A1(n729), .A2(n663), .ZN(n645) );
  INV_X1 U730 ( .A(KEYINPUT67), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n647), .B(KEYINPUT32), .ZN(n648) );
  AND2_X1 U732 ( .A1(n649), .A2(n732), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n650), .A2(n445), .ZN(n651) );
  OR2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n683) );
  INV_X1 U735 ( .A(n729), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n654), .A2(n653), .ZN(n739) );
  XNOR2_X1 U737 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n655) );
  NOR2_X1 U738 ( .A1(n657), .A2(n658), .ZN(n659) );
  AND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n708) );
  NOR2_X1 U740 ( .A1(n719), .A2(n708), .ZN(n661) );
  NOR2_X1 U741 ( .A1(n661), .A2(n487), .ZN(n662) );
  XNOR2_X1 U742 ( .A(n662), .B(KEYINPUT109), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n445), .A2(n663), .ZN(n665) );
  NOR2_X1 U744 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U745 ( .A1(n698), .A2(KEYINPUT44), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n670) );
  INV_X1 U747 ( .A(KEYINPUT2), .ZN(n671) );
  INV_X1 U748 ( .A(n673), .ZN(n674) );
  INV_X1 U749 ( .A(KEYINPUT66), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n774), .A2(G478), .ZN(n678) );
  INV_X1 U751 ( .A(G952), .ZN(n679) );
  XOR2_X1 U752 ( .A(G125), .B(KEYINPUT37), .Z(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(G27) );
  XNOR2_X1 U754 ( .A(n683), .B(G110), .ZN(G12) );
  NOR2_X1 U755 ( .A1(n684), .A2(n685), .ZN(n686) );
  XOR2_X1 U756 ( .A(G146), .B(n686), .Z(G48) );
  XNOR2_X1 U757 ( .A(n687), .B(G134), .ZN(G36) );
  NAND2_X1 U758 ( .A1(n398), .A2(G475), .ZN(n689) );
  XNOR2_X1 U759 ( .A(n689), .B(n486), .ZN(n690) );
  NAND2_X1 U760 ( .A1(n767), .A2(G472), .ZN(n694) );
  BUF_X1 U761 ( .A(n691), .Z(n693) );
  XNOR2_X1 U762 ( .A(KEYINPUT118), .B(KEYINPUT62), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n694), .B(n483), .ZN(n695) );
  XNOR2_X1 U764 ( .A(KEYINPUT119), .B(KEYINPUT63), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n697), .B(G143), .ZN(G45) );
  XOR2_X1 U766 ( .A(G122), .B(n698), .Z(G24) );
  NAND2_X1 U767 ( .A1(n767), .A2(G210), .ZN(n702) );
  XNOR2_X1 U768 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n704), .B(G131), .ZN(G33) );
  XNOR2_X1 U770 ( .A(n705), .B(G119), .ZN(G21) );
  XNOR2_X1 U771 ( .A(G101), .B(n706), .ZN(G3) );
  NAND2_X1 U772 ( .A1(n708), .A2(n716), .ZN(n707) );
  XNOR2_X1 U773 ( .A(n707), .B(G104), .ZN(G6) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n710) );
  NAND2_X1 U775 ( .A1(n708), .A2(n718), .ZN(n709) );
  XNOR2_X1 U776 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(G107), .B(n711), .ZN(G9) );
  XOR2_X1 U778 ( .A(KEYINPUT29), .B(KEYINPUT120), .Z(n714) );
  NOR2_X1 U779 ( .A1(n684), .A2(n712), .ZN(n713) );
  XOR2_X1 U780 ( .A(n714), .B(n713), .Z(n715) );
  XNOR2_X1 U781 ( .A(G128), .B(n715), .ZN(G30) );
  NAND2_X1 U782 ( .A1(n719), .A2(n716), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(G113), .ZN(G15) );
  NAND2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U785 ( .A(n720), .B(G116), .ZN(G18) );
  NOR2_X1 U786 ( .A1(n778), .A2(KEYINPUT2), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT86), .ZN(n725) );
  BUF_X1 U788 ( .A(n722), .Z(n723) );
  NOR2_X1 U789 ( .A1(n723), .A2(KEYINPUT2), .ZN(n724) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U791 ( .A1(n726), .A2(n727), .ZN(n764) );
  XOR2_X1 U792 ( .A(KEYINPUT122), .B(KEYINPUT50), .Z(n731) );
  NAND2_X1 U793 ( .A1(n445), .A2(n728), .ZN(n730) );
  XOR2_X1 U794 ( .A(n731), .B(n730), .Z(n738) );
  XOR2_X1 U795 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n735) );
  NAND2_X1 U796 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U797 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U798 ( .A1(n736), .A2(n657), .ZN(n737) );
  NAND2_X1 U799 ( .A1(n738), .A2(n737), .ZN(n740) );
  NAND2_X1 U800 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U801 ( .A(n741), .B(KEYINPUT123), .ZN(n742) );
  XOR2_X1 U802 ( .A(KEYINPUT51), .B(n742), .Z(n744) );
  INV_X1 U803 ( .A(n743), .ZN(n759) );
  NOR2_X1 U804 ( .A1(n744), .A2(n759), .ZN(n755) );
  NOR2_X1 U805 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U807 ( .A(n749), .B(KEYINPUT124), .ZN(n752) );
  NOR2_X1 U808 ( .A1(n750), .A2(n487), .ZN(n751) );
  NOR2_X1 U809 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U810 ( .A1(n760), .A2(n753), .ZN(n754) );
  NOR2_X1 U811 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U812 ( .A(n756), .B(KEYINPUT52), .ZN(n757) );
  NOR2_X1 U813 ( .A1(n758), .A2(n757), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n760), .A2(n759), .ZN(n761) );
  OR2_X1 U815 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U816 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U817 ( .A1(n765), .A2(G953), .ZN(n766) );
  XNOR2_X1 U818 ( .A(n766), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U819 ( .A1(n774), .A2(G469), .ZN(n772) );
  XOR2_X1 U820 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n768) );
  XOR2_X1 U821 ( .A(n768), .B(KEYINPUT125), .Z(n769) );
  XNOR2_X1 U822 ( .A(n349), .B(n769), .ZN(n771) );
  XNOR2_X1 U823 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U824 ( .A1(n777), .A2(n773), .ZN(G54) );
  NAND2_X1 U825 ( .A1(n774), .A2(G217), .ZN(n776) );
  NAND2_X1 U826 ( .A1(n778), .A2(n354), .ZN(n783) );
  NAND2_X1 U827 ( .A1(G224), .A2(G953), .ZN(n779) );
  XNOR2_X1 U828 ( .A(n779), .B(KEYINPUT126), .ZN(n780) );
  XNOR2_X1 U829 ( .A(KEYINPUT61), .B(n780), .ZN(n781) );
  NAND2_X1 U830 ( .A1(n781), .A2(G898), .ZN(n782) );
  NAND2_X1 U831 ( .A1(n783), .A2(n782), .ZN(n788) );
  XOR2_X1 U832 ( .A(G101), .B(n784), .Z(n786) );
  NOR2_X1 U833 ( .A1(n354), .A2(G898), .ZN(n785) );
  NOR2_X1 U834 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U835 ( .A(n788), .B(n787), .ZN(G69) );
  BUF_X1 U836 ( .A(n789), .Z(n790) );
  XNOR2_X1 U837 ( .A(n792), .B(n791), .ZN(n793) );
  XNOR2_X1 U838 ( .A(n790), .B(n793), .ZN(n796) );
  XNOR2_X1 U839 ( .A(n723), .B(n796), .ZN(n795) );
  NAND2_X1 U840 ( .A1(n795), .A2(n354), .ZN(n801) );
  XOR2_X1 U841 ( .A(G227), .B(n796), .Z(n797) );
  NAND2_X1 U842 ( .A1(n797), .A2(G900), .ZN(n798) );
  XOR2_X1 U843 ( .A(KEYINPUT127), .B(n798), .Z(n799) );
  NAND2_X1 U844 ( .A1(G953), .A2(n799), .ZN(n800) );
  NAND2_X1 U845 ( .A1(n801), .A2(n800), .ZN(G72) );
  XNOR2_X1 U846 ( .A(G140), .B(n802), .ZN(G42) );
  XOR2_X1 U847 ( .A(n803), .B(G137), .Z(G39) );
endmodule

