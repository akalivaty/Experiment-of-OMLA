//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OR2_X1    g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n188), .A2(G146), .A3(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(G146), .B1(new_n188), .B2(new_n191), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n196), .A2(KEYINPUT72), .A3(G119), .ZN(new_n197));
  INV_X1    g011(.A(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT72), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G119), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT73), .B1(new_n198), .B2(G128), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .B1(new_n198), .B2(G128), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n202), .A2(KEYINPUT73), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n203), .A2(new_n205), .B1(G110), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n195), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT74), .B(G110), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n201), .A2(new_n202), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n204), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n207), .A2(KEYINPUT75), .A3(new_n209), .A4(new_n213), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n192), .B1(new_n221), .B2(new_n187), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT76), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n226), .A2(new_n228), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n212), .A2(new_n223), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(KEYINPUT77), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n229), .B2(new_n230), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n195), .A2(new_n211), .B1(new_n220), .B2(new_n222), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n232), .B(new_n233), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n212), .A2(new_n223), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(KEYINPUT25), .A3(new_n233), .A4(new_n232), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G217), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(G234), .B2(new_n233), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n233), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(KEYINPUT78), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n252), .A3(new_n232), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G134), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  INV_X1    g071(.A(G134), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n257), .B1(new_n258), .B2(G137), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n259), .B2(KEYINPUT11), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n257), .B(new_n261), .C1(new_n258), .C2(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(G137), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n265), .A2(new_n266), .A3(new_n262), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(KEYINPUT0), .B2(G128), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT0), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n196), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n270), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  INV_X1    g089(.A(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(KEYINPUT65), .A2(G143), .ZN(new_n278));
  AOI21_X1  g092(.A(G146), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n221), .A2(G143), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n273), .B(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(G146), .A3(new_n278), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n276), .A2(G146), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n282), .A2(KEYINPUT0), .A3(G128), .A4(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n258), .A2(G137), .ZN(new_n287));
  OAI21_X1  g101(.A(G131), .B1(new_n287), .B2(new_n256), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n268), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n291));
  OAI21_X1  g105(.A(G128), .B1(new_n291), .B2(new_n283), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT65), .A2(G143), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT65), .A2(G143), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n221), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n280), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n282), .A2(G128), .A3(new_n291), .A4(new_n284), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n269), .A2(new_n286), .B1(new_n290), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G116), .B(G119), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT2), .B(G113), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n307), .A2(new_n224), .A3(G210), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n306), .B(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n307), .A2(new_n224), .A3(G210), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n306), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n310), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n290), .A2(new_n300), .ZN(new_n318));
  INV_X1    g132(.A(new_n268), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n266), .B1(new_n260), .B2(new_n262), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n285), .B(new_n281), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT67), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n289), .A2(new_n323), .B1(new_n298), .B2(new_n299), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n268), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n324), .A2(new_n325), .B1(new_n269), .B2(new_n286), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n322), .B1(new_n317), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n305), .B(new_n316), .C1(new_n327), .C2(new_n304), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n281), .A2(new_n285), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(new_n268), .B2(new_n264), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n293), .A2(new_n294), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n283), .B1(new_n333), .B2(G146), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT1), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT68), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT68), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT1), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n336), .A2(new_n338), .A3(G128), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n334), .A2(new_n339), .B1(new_n292), .B2(new_n297), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n289), .ZN(new_n341));
  XOR2_X1   g155(.A(G116), .B(G119), .Z(new_n342));
  XNOR2_X1  g156(.A(new_n342), .B(new_n303), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n332), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(KEYINPUT30), .B1(new_n332), .B2(new_n341), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n289), .A2(new_n323), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n325), .A3(new_n300), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n317), .A3(new_n321), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n349), .B2(new_n343), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT31), .A3(new_n316), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n347), .A2(new_n321), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n343), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n301), .B2(new_n304), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n354), .A2(new_n318), .A3(new_n321), .A4(new_n304), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT70), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n316), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n312), .A2(new_n315), .A3(KEYINPUT70), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n330), .A2(new_n351), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(G472), .A2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT32), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n362), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT31), .B1(new_n350), .B2(new_n316), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n304), .B1(new_n345), .B2(new_n348), .ZN(new_n369));
  INV_X1    g183(.A(new_n316), .ZN(new_n370));
  NOR4_X1   g184(.A1(new_n369), .A2(new_n344), .A3(new_n329), .A4(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT32), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(new_n364), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n350), .A2(new_n316), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n361), .B(new_n353), .C1(new_n355), .C2(new_n356), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT71), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n370), .B1(new_n369), .B2(new_n344), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT71), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n378), .A4(new_n377), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n301), .A2(new_n304), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n305), .A2(KEYINPUT28), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n301), .A2(new_n354), .A3(new_n304), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n370), .A2(new_n378), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n380), .A2(new_n383), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G472), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n254), .B1(new_n375), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT9), .B(G234), .ZN(new_n393));
  OAI21_X1  g207(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n269), .ZN(new_n396));
  INV_X1    g210(.A(G104), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT3), .B1(new_n397), .B2(G107), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n399), .A3(G104), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g219(.A1(KEYINPUT80), .A2(G101), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(G107), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT80), .A2(G101), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n401), .B(KEYINPUT10), .C1(new_n405), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n410), .B1(new_n299), .B2(new_n298), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(new_n404), .A3(new_n407), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT4), .B1(new_n405), .B2(new_n409), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n406), .A2(new_n408), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n402), .A3(new_n404), .A4(new_n407), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(G101), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT81), .A4(KEYINPUT4), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n413), .A2(new_n422), .A3(G101), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n281), .A2(new_n423), .A3(new_n285), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n411), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n282), .A2(new_n284), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT65), .B(G143), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n335), .B1(new_n428), .B2(new_n221), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n429), .B2(new_n196), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n299), .A2(KEYINPUT82), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n339), .A2(new_n432), .A3(new_n284), .A4(new_n282), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n418), .A2(new_n401), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n396), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT10), .B1(new_n434), .B2(new_n435), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n424), .B1(new_n416), .B2(new_n420), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n441), .A2(new_n442), .A3(new_n411), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT83), .B1(new_n443), .B2(new_n396), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n426), .A2(new_n438), .A3(KEYINPUT83), .A4(new_n396), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n224), .A2(G227), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n426), .A2(new_n438), .A3(new_n396), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n439), .B1(new_n455), .B2(new_n445), .ZN(new_n456));
  INV_X1    g270(.A(new_n450), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n450), .B1(new_n455), .B2(new_n445), .ZN(new_n459));
  OR3_X1    g273(.A1(new_n435), .A2(new_n300), .A3(KEYINPUT84), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT84), .B1(new_n435), .B2(new_n300), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n436), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT12), .A3(new_n269), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT12), .B1(new_n462), .B2(new_n269), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G469), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n233), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n233), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n455), .A2(new_n445), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n464), .B2(new_n465), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n450), .B(KEYINPUT79), .Z(new_n473));
  AOI22_X1  g287(.A1(new_n472), .A2(new_n473), .B1(new_n459), .B2(new_n440), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n474), .B2(G469), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n395), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G110), .B(G122), .Z(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT8), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n342), .A2(new_n303), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n198), .A3(G116), .ZN(new_n481));
  OAI211_X1 g295(.A(G113), .B(new_n481), .C1(new_n342), .C2(new_n480), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n435), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n418), .A2(new_n401), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n478), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G125), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n298), .A2(new_n488), .A3(new_n299), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT90), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n298), .A2(new_n491), .A3(new_n488), .A4(new_n299), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n331), .A2(G125), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n224), .A2(G224), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT7), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n487), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT89), .B1(new_n331), .B2(G125), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n501), .B(new_n488), .C1(new_n281), .C2(new_n285), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT7), .B1(new_n496), .B2(KEYINPUT91), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(KEYINPUT91), .B2(new_n496), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n493), .A2(new_n500), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT92), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n499), .A2(new_n502), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n493), .A4(new_n505), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n498), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n343), .A2(new_n423), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n421), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n477), .ZN(new_n515));
  AND4_X1   g329(.A1(KEYINPUT87), .A2(new_n514), .A3(new_n515), .A4(new_n483), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n484), .A2(new_n485), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n517), .B1(new_n421), .B2(new_n513), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT87), .B1(new_n518), .B2(new_n515), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G902), .B1(new_n511), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n512), .B1(new_n416), .B2(new_n420), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n477), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT88), .B1(new_n523), .B2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n483), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT88), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n477), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n508), .A2(new_n493), .ZN(new_n530));
  INV_X1    g344(.A(new_n496), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n516), .A2(new_n519), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n534), .A3(new_n477), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT86), .B1(new_n518), .B2(new_n515), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(KEYINPUT6), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n529), .B(new_n532), .C1(new_n533), .C2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(G210), .B1(G237), .B2(G902), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT93), .Z(new_n540));
  AND3_X1   g354(.A1(new_n521), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n521), .B2(new_n538), .ZN(new_n542));
  OAI21_X1  g356(.A(G214), .B1(G237), .B2(G902), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT100), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(KEYINPUT20), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT99), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n307), .A2(new_n224), .A3(G214), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n550), .A2(new_n277), .A3(KEYINPUT94), .A4(new_n278), .ZN(new_n551));
  INV_X1    g365(.A(G214), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n552), .A2(G237), .A3(G953), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G143), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(KEYINPUT94), .B1(new_n333), .B2(new_n550), .ZN(new_n556));
  OAI21_X1  g370(.A(G131), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n428), .B2(new_n553), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n266), .A3(new_n554), .A4(new_n551), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n549), .B1(new_n561), .B2(KEYINPUT17), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT17), .B(G131), .C1(new_n555), .C2(new_n556), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n194), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n557), .A2(KEYINPUT99), .A3(new_n565), .A4(new_n560), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G113), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n397), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT18), .B(G131), .C1(new_n555), .C2(new_n556), .ZN(new_n570));
  NAND2_X1  g384(.A1(KEYINPUT18), .A2(G131), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n559), .A2(new_n571), .A3(new_n554), .A4(new_n551), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n187), .B(new_n221), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT95), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n570), .A2(new_n576), .A3(new_n572), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n567), .A2(new_n569), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n187), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n488), .A2(G140), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n190), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT97), .B1(new_n585), .B2(new_n580), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(KEYINPUT19), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n192), .B1(new_n588), .B2(new_n221), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n575), .A2(new_n577), .B1(new_n589), .B2(new_n561), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT98), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n569), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n579), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(G475), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n547), .B(new_n548), .C1(new_n594), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n589), .A2(new_n561), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n578), .A2(new_n591), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n569), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n590), .A2(new_n591), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n567), .A2(new_n578), .ZN(new_n603));
  OAI22_X1  g417(.A1(new_n601), .A2(new_n602), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(new_n546), .A3(KEYINPUT20), .A4(new_n595), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n569), .B1(new_n567), .B2(new_n578), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n579), .A2(new_n606), .A3(KEYINPUT101), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(KEYINPUT101), .A3(new_n600), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n233), .ZN(new_n609));
  OAI21_X1  g423(.A(G475), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n333), .A2(G128), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n196), .A2(G143), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n258), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n611), .A2(new_n258), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g430(.A1(KEYINPUT102), .A2(G122), .ZN(new_n617));
  NAND2_X1  g431(.A1(KEYINPUT102), .A2(G122), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G116), .ZN(new_n620));
  INV_X1    g434(.A(G116), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G122), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n399), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(KEYINPUT14), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n621), .B1(new_n617), .B2(new_n618), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT103), .B(G107), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n625), .A3(new_n624), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n630), .B2(G107), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n616), .B(new_n623), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n620), .A2(new_n622), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(G107), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n611), .A2(KEYINPUT13), .A3(new_n612), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n636), .B(G134), .C1(KEYINPUT13), .C2(new_n611), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n637), .A3(new_n615), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n393), .A2(new_n247), .A3(G953), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n632), .A2(new_n638), .A3(new_n640), .ZN(new_n643));
  AOI21_X1  g457(.A(G902), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G478), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(KEYINPUT15), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n597), .A2(new_n605), .A3(new_n610), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(G234), .A2(G237), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(G952), .A3(new_n224), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(G902), .A3(G953), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT104), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT21), .B(G898), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n392), .A2(new_n476), .A3(new_n545), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(new_n417), .Z(G3));
  OAI21_X1  g471(.A(G472), .B1(new_n363), .B2(G902), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n365), .B2(new_n363), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n254), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n521), .A2(new_n538), .ZN(new_n661));
  INV_X1    g475(.A(new_n540), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n521), .A2(new_n538), .A3(new_n540), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n543), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n654), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n660), .A2(new_n476), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n597), .A2(new_n610), .A3(new_n605), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n641), .B2(KEYINPUT105), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n643), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n640), .B1(new_n632), .B2(new_n638), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n642), .A2(new_n643), .A3(new_n670), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n645), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n645), .B(new_n233), .C1(new_n672), .C2(new_n673), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n645), .A2(new_n233), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(KEYINPUT106), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n672), .A2(new_n673), .A3(new_n671), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n670), .B1(new_n642), .B2(new_n643), .ZN(new_n683));
  OAI21_X1  g497(.A(G478), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n678), .B1(new_n644), .B2(new_n645), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n668), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n667), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT34), .B(G104), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G6));
  NAND2_X1  g506(.A1(new_n597), .A2(new_n605), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n647), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n610), .A2(new_n696), .ZN(new_n697));
  OAI211_X1 g511(.A(KEYINPUT107), .B(G475), .C1(new_n607), .C2(new_n609), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n694), .A2(new_n695), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n667), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G107), .ZN(new_n702));
  XNOR2_X1  g516(.A(KEYINPUT108), .B(KEYINPUT35), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n238), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n242), .B1(new_n243), .B2(KEYINPUT36), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n707), .A2(new_n252), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n249), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n250), .B1(new_n241), .B2(new_n245), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT109), .B1(new_n712), .B2(new_n709), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n659), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n476), .A3(new_n655), .A4(new_n545), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT37), .B(G110), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G12));
  AOI21_X1  g532(.A(new_n714), .B1(new_n375), .B2(new_n391), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n697), .A2(new_n698), .ZN(new_n720));
  INV_X1    g534(.A(G900), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n650), .B1(new_n652), .B2(new_n721), .ZN(new_n722));
  NOR4_X1   g536(.A1(new_n720), .A2(new_n693), .A3(new_n647), .A4(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n719), .A2(new_n723), .A3(new_n476), .A4(new_n545), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  NAND2_X1  g539(.A1(new_n663), .A2(new_n664), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT38), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n362), .B1(new_n384), .B2(new_n344), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n328), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(G472), .B1(new_n730), .B2(G902), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n375), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n668), .A2(new_n695), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n711), .A2(new_n713), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n733), .A2(new_n544), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n728), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n722), .B(KEYINPUT39), .Z(new_n737));
  NAND2_X1  g551(.A1(new_n476), .A2(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT40), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n333), .B(KEYINPUT110), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G45));
  INV_X1    g557(.A(new_n722), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n668), .A2(new_n688), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n719), .A2(new_n476), .A3(new_n545), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G146), .ZN(G48));
  INV_X1    g561(.A(new_n469), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n468), .B1(new_n467), .B2(new_n233), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n748), .A2(new_n749), .A3(new_n395), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n392), .A3(new_n689), .A4(new_n666), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  NAND4_X1  g567(.A1(new_n750), .A2(new_n700), .A3(new_n392), .A4(new_n666), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G116), .ZN(G18));
  INV_X1    g569(.A(new_n648), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n750), .A2(new_n719), .A3(new_n756), .A4(new_n666), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G119), .ZN(G21));
  INV_X1    g572(.A(new_n254), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n387), .A2(new_n361), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n330), .B2(new_n351), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n760), .B1(new_n762), .B2(new_n365), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n368), .A2(new_n371), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT111), .B(new_n364), .C1(new_n764), .C2(new_n761), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n759), .A2(new_n658), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n733), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n750), .A2(new_n766), .A3(new_n666), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND4_X1  g583(.A1(new_n734), .A2(new_n658), .A3(new_n763), .A4(new_n765), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n668), .A2(new_n688), .A3(new_n744), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n750), .A3(new_n545), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n469), .A2(new_n475), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n544), .B1(new_n663), .B2(new_n664), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n394), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n775), .B1(new_n476), .B2(new_n777), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n392), .B(new_n745), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT113), .B(KEYINPUT42), .Z(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n776), .A2(new_n777), .A3(new_n394), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT112), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n476), .A2(new_n775), .A3(new_n777), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(KEYINPUT113), .A2(KEYINPUT42), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n787), .A2(new_n392), .A3(new_n745), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G131), .ZN(G33));
  OAI211_X1 g606(.A(new_n392), .B(new_n723), .C1(new_n778), .C2(new_n779), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  AND2_X1   g608(.A1(new_n681), .A2(new_n687), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n668), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT43), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n659), .A2(new_n734), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT44), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n777), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n474), .A2(KEYINPUT45), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n468), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n474), .A2(KEYINPUT45), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n470), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(KEYINPUT46), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n469), .B1(new_n806), .B2(KEYINPUT46), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n394), .B(new_n737), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n810), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n802), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(new_n255), .ZN(G39));
  NAND4_X1  g629(.A1(new_n777), .A2(new_n375), .A3(new_n391), .A4(new_n254), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n394), .B1(new_n807), .B2(new_n808), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n771), .B(new_n816), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(new_n189), .ZN(G42));
  NAND3_X1  g636(.A1(new_n759), .A2(new_n394), .A3(new_n543), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n728), .A2(new_n668), .A3(new_n795), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n467), .A2(new_n233), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(G469), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n469), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n732), .B1(new_n827), .B2(KEYINPUT49), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n824), .B(new_n828), .C1(KEYINPUT49), .C2(new_n827), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT115), .Z(new_n830));
  INV_X1    g644(.A(new_n766), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n797), .A2(new_n650), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT117), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n777), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n819), .B(new_n820), .C1(new_n394), .C2(new_n827), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT118), .ZN(new_n839));
  INV_X1    g653(.A(new_n750), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n728), .A3(new_n543), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT50), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n777), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n732), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n759), .A3(new_n650), .A4(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n668), .A3(new_n688), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n833), .A2(new_n834), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n850), .A2(new_n846), .ZN(new_n851));
  INV_X1    g665(.A(new_n770), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n844), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n839), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n689), .ZN(new_n856));
  OAI211_X1 g670(.A(G952), .B(new_n224), .C1(new_n848), .C2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n545), .A2(new_n826), .A3(new_n394), .A4(new_n469), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n835), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n851), .B2(new_n392), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n861), .A2(new_n850), .A3(new_n392), .A4(new_n846), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n844), .A2(new_n838), .A3(KEYINPUT51), .A4(new_n853), .ZN(new_n867));
  OAI211_X1 g681(.A(KEYINPUT119), .B(new_n860), .C1(new_n862), .C2(new_n863), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n751), .A2(new_n754), .A3(new_n656), .A4(new_n716), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n756), .B1(new_n668), .B2(new_n795), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n660), .A3(new_n476), .A4(new_n666), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n757), .A2(new_n768), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n720), .A2(new_n693), .A3(new_n695), .A4(new_n722), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n719), .A2(new_n876), .A3(new_n476), .A4(new_n777), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n793), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n791), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n665), .A2(new_n733), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n712), .A2(new_n709), .A3(new_n722), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n476), .A3(new_n732), .A4(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n773), .A2(new_n724), .A3(new_n746), .A4(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT52), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT53), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n879), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n776), .A2(new_n545), .A3(new_n394), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n372), .A2(new_n373), .A3(new_n364), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n373), .B1(new_n372), .B2(new_n364), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n391), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n734), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n697), .A2(new_n698), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(new_n694), .A3(new_n695), .A4(new_n744), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n889), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n658), .A2(new_n763), .A3(new_n765), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n745), .A3(new_n734), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n858), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT116), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n773), .A2(new_n724), .A3(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n900), .A2(new_n746), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n879), .B1(new_n888), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n886), .B1(KEYINPUT53), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n885), .B1(new_n879), .B2(new_n884), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n888), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n793), .A2(new_n875), .A3(new_n877), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n910), .A2(new_n873), .A3(new_n870), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(new_n911), .A3(KEYINPUT53), .A4(new_n791), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n855), .A2(new_n869), .A3(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(G952), .A2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n830), .B1(new_n916), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n224), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n233), .B1(new_n908), .B2(new_n912), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(new_n540), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n529), .B1(new_n537), .B2(new_n533), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(new_n532), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n920), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n922), .B2(new_n925), .ZN(G51));
  XNOR2_X1  g741(.A(new_n913), .B(KEYINPUT54), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n470), .B(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n467), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n921), .A2(new_n805), .A3(new_n804), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n919), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND3_X1  g747(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n919), .B1(new_n934), .B2(new_n594), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n594), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(KEYINPUT120), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(KEYINPUT120), .B2(new_n936), .ZN(G60));
  NAND2_X1  g752(.A1(new_n674), .A2(new_n675), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT121), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n678), .B(KEYINPUT59), .Z(new_n941));
  AOI21_X1  g755(.A(new_n940), .B1(new_n915), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n928), .A2(new_n940), .A3(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n919), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n913), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(KEYINPUT122), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n244), .A2(new_n232), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n913), .A2(new_n951), .A3(new_n947), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n707), .A2(new_n708), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT123), .Z(new_n955));
  AOI21_X1  g769(.A(new_n951), .B1(new_n913), .B2(new_n947), .ZN(new_n956));
  AOI211_X1 g770(.A(KEYINPUT122), .B(new_n946), .C1(new_n908), .C2(new_n912), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n958), .A3(new_n920), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n956), .A2(new_n957), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n919), .B1(new_n964), .B2(new_n950), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n960), .A4(new_n958), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n963), .A2(new_n966), .ZN(G66));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n653), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n874), .B2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n923), .B1(G898), .B2(new_n224), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G69));
  XNOR2_X1  g786(.A(new_n327), .B(new_n588), .ZN(new_n973));
  NAND3_X1  g787(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n871), .A2(new_n392), .A3(new_n777), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(new_n738), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT125), .Z(new_n977));
  NOR3_X1   g791(.A1(new_n814), .A2(new_n821), .A3(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n900), .A2(new_n746), .A3(new_n902), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n741), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n973), .B(new_n974), .C1(new_n983), .C2(G953), .ZN(new_n984));
  INV_X1    g798(.A(new_n793), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n814), .A2(new_n821), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n813), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n392), .B(new_n880), .C1(new_n987), .C2(new_n811), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n979), .A2(new_n791), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n986), .A2(new_n993), .A3(new_n988), .A4(new_n990), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n721), .A2(new_n224), .A3(G227), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n973), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n984), .B1(new_n995), .B2(new_n997), .ZN(G72));
  XNOR2_X1  g812(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n874), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1001), .B1(new_n983), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n350), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1003), .A2(new_n316), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n328), .A2(new_n381), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n906), .A2(new_n1001), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1005), .A2(new_n1007), .A3(new_n920), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n350), .A2(new_n370), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n992), .A2(new_n994), .A3(new_n874), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1009), .B1(new_n1010), .B2(new_n1001), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1008), .A2(new_n1011), .ZN(G57));
endmodule


