

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767;

  NOR2_X1 U374 ( .A1(n753), .A2(n418), .ZN(n686) );
  NAND2_X1 U375 ( .A1(n363), .A2(n625), .ZN(n753) );
  XNOR2_X1 U376 ( .A(n622), .B(n621), .ZN(n363) );
  OR2_X1 U377 ( .A1(n642), .A2(n626), .ZN(n485) );
  XNOR2_X1 U378 ( .A(n750), .B(n446), .ZN(n465) );
  INV_X2 U379 ( .A(G128), .ZN(n392) );
  INV_X2 U380 ( .A(G953), .ZN(n754) );
  NOR2_X2 U381 ( .A1(n557), .A2(n527), .ZN(n705) );
  XNOR2_X1 U382 ( .A(n446), .B(G125), .ZN(n473) );
  NAND2_X1 U383 ( .A1(n619), .A2(n708), .ZN(n611) );
  BUF_X1 U384 ( .A(n655), .Z(n731) );
  NAND2_X1 U385 ( .A1(n705), .A2(n703), .ZN(n711) );
  NAND2_X1 U386 ( .A1(n424), .A2(n421), .ZN(n367) );
  NAND2_X1 U387 ( .A1(n423), .A2(n422), .ZN(n421) );
  XNOR2_X1 U388 ( .A(n365), .B(n361), .ZN(n535) );
  NAND2_X2 U389 ( .A1(n689), .A2(n690), .ZN(n369) );
  XNOR2_X1 U390 ( .A(n397), .B(n470), .ZN(n742) );
  XNOR2_X1 U391 ( .A(n472), .B(n471), .ZN(n397) );
  XNOR2_X1 U392 ( .A(n447), .B(n473), .ZN(n748) );
  NAND2_X1 U393 ( .A1(n754), .A2(G234), .ZN(n405) );
  XNOR2_X2 U394 ( .A(n584), .B(KEYINPUT81), .ZN(n669) );
  XNOR2_X2 U395 ( .A(n400), .B(KEYINPUT0), .ZN(n551) );
  XNOR2_X1 U396 ( .A(n369), .B(n458), .ZN(n545) );
  INV_X1 U397 ( .A(KEYINPUT76), .ZN(n458) );
  AND2_X1 U398 ( .A1(n637), .A2(KEYINPUT66), .ZN(n394) );
  NOR2_X1 U399 ( .A1(n766), .A2(n767), .ZN(n407) );
  INV_X1 U400 ( .A(n639), .ZN(n389) );
  AND2_X1 U401 ( .A1(n408), .A2(n389), .ZN(n382) );
  XNOR2_X1 U402 ( .A(KEYINPUT15), .B(G902), .ZN(n569) );
  XOR2_X1 U403 ( .A(G116), .B(KEYINPUT97), .Z(n460) );
  XNOR2_X1 U404 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n402) );
  INV_X1 U405 ( .A(KEYINPUT8), .ZN(n440) );
  XOR2_X1 U406 ( .A(G140), .B(G104), .Z(n503) );
  XNOR2_X1 U407 ( .A(G143), .B(G113), .ZN(n502) );
  XNOR2_X1 U408 ( .A(n501), .B(n430), .ZN(n429) );
  XNOR2_X1 U409 ( .A(n431), .B(KEYINPUT4), .ZN(n430) );
  INV_X1 U410 ( .A(G137), .ZN(n431) );
  INV_X1 U411 ( .A(KEYINPUT39), .ZN(n379) );
  NAND2_X1 U412 ( .A1(n376), .A2(n380), .ZN(n375) );
  NOR2_X1 U413 ( .A1(n591), .A2(n377), .ZN(n376) );
  NAND2_X1 U414 ( .A1(n360), .A2(KEYINPUT39), .ZN(n377) );
  INV_X1 U415 ( .A(KEYINPUT92), .ZN(n366) );
  XOR2_X1 U416 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n434) );
  INV_X1 U417 ( .A(G101), .ZN(n436) );
  XNOR2_X1 U418 ( .A(n396), .B(G107), .ZN(n470) );
  XNOR2_X1 U419 ( .A(G110), .B(G104), .ZN(n396) );
  XNOR2_X1 U420 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n476) );
  INV_X1 U421 ( .A(n686), .ZN(n417) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n413) );
  NAND2_X1 U423 ( .A1(n628), .A2(n506), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n454), .B(KEYINPUT25), .ZN(n411) );
  OR2_X2 U425 ( .A1(n732), .A2(G902), .ZN(n412) );
  BUF_X1 U426 ( .A(G953), .Z(n759) );
  NAND2_X1 U427 ( .A1(n353), .A2(n371), .ZN(n601) );
  NOR2_X1 U428 ( .A1(n694), .A2(n693), .ZN(n690) );
  XNOR2_X1 U429 ( .A(n570), .B(KEYINPUT84), .ZN(n368) );
  NOR2_X1 U430 ( .A1(n736), .A2(n569), .ZN(n570) );
  AND2_X1 U431 ( .A1(n638), .A2(n394), .ZN(n393) );
  NAND2_X1 U432 ( .A1(n383), .A2(n381), .ZN(n622) );
  NAND2_X1 U433 ( .A1(n355), .A2(n382), .ZN(n381) );
  NAND2_X1 U434 ( .A1(n384), .A2(n389), .ZN(n383) );
  INV_X1 U435 ( .A(G902), .ZN(n506) );
  XNOR2_X1 U436 ( .A(n465), .B(n464), .ZN(n628) );
  XNOR2_X1 U437 ( .A(n404), .B(n401), .ZN(n445) );
  XNOR2_X1 U438 ( .A(n403), .B(n402), .ZN(n401) );
  XNOR2_X1 U439 ( .A(G119), .B(KEYINPUT78), .ZN(n403) );
  XNOR2_X1 U440 ( .A(G137), .B(G128), .ZN(n443) );
  INV_X1 U441 ( .A(G134), .ZN(n391) );
  XNOR2_X1 U442 ( .A(n505), .B(n504), .ZN(n647) );
  NAND2_X1 U443 ( .A1(n545), .A2(n608), .ZN(n469) );
  NAND2_X1 U444 ( .A1(n373), .A2(n379), .ZN(n372) );
  AND2_X1 U445 ( .A1(n378), .A2(n375), .ZN(n374) );
  NAND2_X1 U446 ( .A1(n371), .A2(n360), .ZN(n373) );
  NOR2_X1 U447 ( .A1(n427), .A2(n426), .ZN(n425) );
  NOR2_X1 U448 ( .A1(n493), .A2(n494), .ZN(n427) );
  INV_X1 U449 ( .A(n594), .ZN(n426) );
  XNOR2_X1 U450 ( .A(n611), .B(KEYINPUT19), .ZN(n583) );
  AND2_X1 U451 ( .A1(n535), .A2(n531), .ZN(n560) );
  XNOR2_X1 U452 ( .A(n438), .B(n465), .ZN(n657) );
  XNOR2_X1 U453 ( .A(n742), .B(n480), .ZN(n642) );
  AND2_X1 U454 ( .A1(n631), .A2(n759), .ZN(n735) );
  NAND2_X1 U455 ( .A1(n419), .A2(KEYINPUT2), .ZN(n418) );
  INV_X1 U456 ( .A(n736), .ZN(n419) );
  XNOR2_X1 U457 ( .A(n537), .B(KEYINPUT32), .ZN(n637) );
  INV_X1 U458 ( .A(G143), .ZN(n636) );
  AND2_X1 U459 ( .A1(n380), .A2(n593), .ZN(n353) );
  AND2_X1 U460 ( .A1(n681), .A2(KEYINPUT48), .ZN(n354) );
  AND2_X1 U461 ( .A1(n406), .A2(n354), .ZN(n355) );
  XOR2_X1 U462 ( .A(n501), .B(KEYINPUT11), .Z(n356) );
  XOR2_X1 U463 ( .A(n435), .B(n749), .Z(n357) );
  AND2_X1 U464 ( .A1(n493), .A2(n494), .ZN(n358) );
  OR2_X1 U465 ( .A1(n575), .A2(n492), .ZN(n359) );
  NOR2_X1 U466 ( .A1(n603), .A2(n592), .ZN(n360) );
  XOR2_X1 U467 ( .A(n530), .B(KEYINPUT22), .Z(n361) );
  XNOR2_X1 U468 ( .A(n450), .B(n449), .ZN(n732) );
  XNOR2_X1 U469 ( .A(KEYINPUT64), .B(n627), .ZN(n362) );
  INV_X1 U470 ( .A(KEYINPUT48), .ZN(n390) );
  NAND2_X1 U471 ( .A1(n657), .A2(n506), .ZN(n414) );
  NAND2_X1 U472 ( .A1(n364), .A2(KEYINPUT44), .ZN(n541) );
  NAND2_X1 U473 ( .A1(n393), .A2(n540), .ZN(n364) );
  NOR2_X2 U474 ( .A1(n551), .A2(n529), .ZN(n365) );
  XNOR2_X2 U475 ( .A(n441), .B(n366), .ZN(n749) );
  XNOR2_X2 U476 ( .A(n367), .B(KEYINPUT35), .ZN(n654) );
  NAND2_X1 U477 ( .A1(n368), .A2(n420), .ZN(n416) );
  NAND2_X1 U478 ( .A1(n655), .A2(G475), .ZN(n649) );
  AND2_X2 U479 ( .A1(n415), .A2(n417), .ZN(n655) );
  NAND2_X1 U480 ( .A1(n583), .A2(n359), .ZN(n400) );
  XNOR2_X2 U481 ( .A(n549), .B(n413), .ZN(n689) );
  NAND2_X1 U482 ( .A1(n587), .A2(n708), .ZN(n589) );
  XNOR2_X2 U483 ( .A(n370), .B(G472), .ZN(n587) );
  INV_X1 U484 ( .A(n591), .ZN(n371) );
  INV_X1 U485 ( .A(n590), .ZN(n380) );
  NAND2_X1 U486 ( .A1(n590), .A2(n379), .ZN(n378) );
  NAND2_X1 U487 ( .A1(n374), .A2(n372), .ZN(n624) );
  NAND2_X1 U488 ( .A1(n387), .A2(n385), .ZN(n384) );
  NAND2_X1 U489 ( .A1(n386), .A2(n390), .ZN(n385) );
  NAND2_X1 U490 ( .A1(n406), .A2(n681), .ZN(n386) );
  NAND2_X1 U491 ( .A1(n388), .A2(n390), .ZN(n387) );
  INV_X1 U492 ( .A(n408), .ZN(n388) );
  XNOR2_X2 U493 ( .A(n474), .B(n391), .ZN(n511) );
  XNOR2_X2 U494 ( .A(n392), .B(G143), .ZN(n474) );
  NAND2_X1 U495 ( .A1(n416), .A2(n362), .ZN(n415) );
  XOR2_X2 U496 ( .A(KEYINPUT68), .B(G140), .Z(n441) );
  XNOR2_X2 U497 ( .A(n395), .B(KEYINPUT104), .ZN(n638) );
  NAND2_X1 U498 ( .A1(n560), .A2(n532), .ZN(n395) );
  XNOR2_X2 U499 ( .A(n399), .B(n398), .ZN(n471) );
  XNOR2_X2 U500 ( .A(KEYINPUT3), .B(G119), .ZN(n398) );
  XNOR2_X2 U501 ( .A(G113), .B(G101), .ZN(n399) );
  NAND2_X1 U502 ( .A1(n512), .A2(G221), .ZN(n404) );
  XNOR2_X2 U503 ( .A(n405), .B(n440), .ZN(n512) );
  XNOR2_X1 U504 ( .A(n407), .B(KEYINPUT46), .ZN(n406) );
  XNOR2_X1 U505 ( .A(n409), .B(KEYINPUT73), .ZN(n408) );
  NAND2_X1 U506 ( .A1(n410), .A2(n598), .ZN(n409) );
  XNOR2_X1 U507 ( .A(n586), .B(n585), .ZN(n410) );
  XNOR2_X2 U508 ( .A(n412), .B(n411), .ZN(n694) );
  INV_X1 U509 ( .A(n689), .ZN(n531) );
  XNOR2_X2 U510 ( .A(n414), .B(n439), .ZN(n549) );
  NOR2_X1 U511 ( .A1(n753), .A2(n736), .ZN(n684) );
  INV_X1 U512 ( .A(n753), .ZN(n420) );
  INV_X1 U513 ( .A(n494), .ZN(n422) );
  INV_X1 U514 ( .A(n721), .ZN(n423) );
  AND2_X2 U515 ( .A1(n428), .A2(n425), .ZN(n424) );
  NAND2_X1 U516 ( .A1(n721), .A2(n358), .ZN(n428) );
  XNOR2_X2 U517 ( .A(n469), .B(n468), .ZN(n721) );
  XNOR2_X2 U518 ( .A(n511), .B(n429), .ZN(n750) );
  NOR2_X2 U519 ( .A1(n650), .A2(n735), .ZN(n653) );
  NOR2_X2 U520 ( .A1(n645), .A2(n735), .ZN(n646) );
  NOR2_X2 U521 ( .A1(n632), .A2(n735), .ZN(n634) );
  BUF_X1 U522 ( .A(n549), .Z(n580) );
  XOR2_X1 U523 ( .A(n503), .B(n502), .Z(n432) );
  INV_X1 U524 ( .A(KEYINPUT85), .ZN(n621) );
  INV_X1 U525 ( .A(n683), .ZN(n625) );
  XNOR2_X1 U526 ( .A(n356), .B(n432), .ZN(n504) );
  XNOR2_X1 U527 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n588) );
  XNOR2_X1 U528 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X2 U529 ( .A(KEYINPUT67), .B(G131), .Z(n501) );
  INV_X2 U530 ( .A(G146), .ZN(n446) );
  NAND2_X1 U531 ( .A1(G227), .A2(n754), .ZN(n433) );
  XNOR2_X1 U532 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U533 ( .A(n470), .B(n436), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n357), .B(n437), .ZN(n438) );
  INV_X1 U535 ( .A(G469), .ZN(n439) );
  INV_X1 U536 ( .A(n441), .ZN(n442) );
  XOR2_X1 U537 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n450) );
  XNOR2_X1 U539 ( .A(G110), .B(KEYINPUT83), .ZN(n448) );
  INV_X1 U540 ( .A(KEYINPUT10), .ZN(n447) );
  XNOR2_X1 U541 ( .A(n448), .B(n748), .ZN(n449) );
  XOR2_X1 U542 ( .A(KEYINPUT94), .B(KEYINPUT20), .Z(n452) );
  NAND2_X1 U543 ( .A1(G234), .A2(n569), .ZN(n451) );
  XNOR2_X1 U544 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U545 ( .A(KEYINPUT93), .B(n453), .ZN(n455) );
  NAND2_X1 U546 ( .A1(n455), .A2(G217), .ZN(n454) );
  AND2_X1 U547 ( .A1(n455), .A2(G221), .ZN(n457) );
  XNOR2_X1 U548 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n456) );
  XNOR2_X1 U549 ( .A(n457), .B(n456), .ZN(n693) );
  XNOR2_X1 U550 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n459) );
  XNOR2_X1 U551 ( .A(n460), .B(n459), .ZN(n462) );
  NOR2_X1 U552 ( .A1(n759), .A2(G237), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n498), .A2(G210), .ZN(n461) );
  XNOR2_X1 U554 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U555 ( .A(n471), .B(n463), .ZN(n464) );
  INV_X1 U556 ( .A(KEYINPUT6), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n587), .B(n466), .ZN(n608) );
  XOR2_X1 U558 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n467) );
  XNOR2_X1 U559 ( .A(n467), .B(KEYINPUT105), .ZN(n468) );
  XNOR2_X2 U560 ( .A(G122), .B(G116), .ZN(n509) );
  XNOR2_X1 U561 ( .A(n509), .B(KEYINPUT16), .ZN(n472) );
  XNOR2_X1 U562 ( .A(n474), .B(n473), .ZN(n479) );
  NAND2_X1 U563 ( .A1(n754), .A2(G224), .ZN(n475) );
  XNOR2_X1 U564 ( .A(n475), .B(KEYINPUT4), .ZN(n477) );
  XNOR2_X1 U565 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U566 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U567 ( .A(n569), .ZN(n626) );
  INV_X1 U568 ( .A(G237), .ZN(n481) );
  NAND2_X1 U569 ( .A1(n506), .A2(n481), .ZN(n486) );
  NAND2_X1 U570 ( .A1(n486), .A2(G210), .ZN(n483) );
  INV_X1 U571 ( .A(KEYINPUT88), .ZN(n482) );
  XNOR2_X1 U572 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X2 U573 ( .A(n485), .B(n484), .ZN(n619) );
  NAND2_X1 U574 ( .A1(n486), .A2(G214), .ZN(n488) );
  INV_X1 U575 ( .A(KEYINPUT89), .ZN(n487) );
  XNOR2_X1 U576 ( .A(n488), .B(n487), .ZN(n708) );
  NAND2_X1 U577 ( .A1(G234), .A2(G237), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n489), .B(KEYINPUT14), .ZN(n491) );
  NAND2_X1 U579 ( .A1(G952), .A2(n491), .ZN(n719) );
  NOR2_X1 U580 ( .A1(n759), .A2(n719), .ZN(n490) );
  XNOR2_X1 U581 ( .A(n490), .B(KEYINPUT90), .ZN(n575) );
  NAND2_X1 U582 ( .A1(G902), .A2(n491), .ZN(n571) );
  XNOR2_X1 U583 ( .A(G898), .B(KEYINPUT91), .ZN(n739) );
  NAND2_X1 U584 ( .A1(n759), .A2(n739), .ZN(n743) );
  NOR2_X1 U585 ( .A1(n571), .A2(n743), .ZN(n492) );
  INV_X1 U586 ( .A(n551), .ZN(n493) );
  XNOR2_X1 U587 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n494) );
  XOR2_X1 U588 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n496) );
  XNOR2_X1 U589 ( .A(G122), .B(KEYINPUT12), .ZN(n495) );
  XNOR2_X1 U590 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U591 ( .A(n748), .B(n497), .Z(n500) );
  NAND2_X1 U592 ( .A1(G214), .A2(n498), .ZN(n499) );
  XNOR2_X1 U593 ( .A(n500), .B(n499), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n647), .A2(n506), .ZN(n508) );
  XOR2_X1 U595 ( .A(KEYINPUT13), .B(G475), .Z(n507) );
  XNOR2_X1 U596 ( .A(n508), .B(n507), .ZN(n557) );
  XOR2_X1 U597 ( .A(KEYINPUT101), .B(G478), .Z(n519) );
  XNOR2_X1 U598 ( .A(n509), .B(G107), .ZN(n510) );
  XNOR2_X1 U599 ( .A(n511), .B(n510), .ZN(n517) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(KEYINPUT100), .Z(n514) );
  NAND2_X1 U601 ( .A1(G217), .A2(n512), .ZN(n513) );
  XNOR2_X1 U602 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U603 ( .A(n515), .B(KEYINPUT7), .Z(n516) );
  XNOR2_X1 U604 ( .A(n517), .B(n516), .ZN(n728) );
  NOR2_X1 U605 ( .A1(G902), .A2(n728), .ZN(n518) );
  XNOR2_X1 U606 ( .A(n519), .B(n518), .ZN(n556) );
  INV_X1 U607 ( .A(n556), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n557), .A2(n527), .ZN(n521) );
  INV_X1 U609 ( .A(KEYINPUT106), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n521), .B(n520), .ZN(n594) );
  INV_X1 U611 ( .A(KEYINPUT44), .ZN(n522) );
  NAND2_X1 U612 ( .A1(n522), .A2(KEYINPUT66), .ZN(n523) );
  OR2_X2 U613 ( .A1(n654), .A2(n523), .ZN(n526) );
  INV_X1 U614 ( .A(KEYINPUT66), .ZN(n524) );
  NAND2_X1 U615 ( .A1(n654), .A2(n524), .ZN(n525) );
  NAND2_X1 U616 ( .A1(n526), .A2(n525), .ZN(n539) );
  INV_X1 U617 ( .A(n693), .ZN(n528) );
  NAND2_X1 U618 ( .A1(n705), .A2(n528), .ZN(n529) );
  INV_X1 U619 ( .A(KEYINPUT72), .ZN(n530) );
  INV_X1 U620 ( .A(n587), .ZN(n554) );
  INV_X1 U621 ( .A(n694), .ZN(n533) );
  NOR2_X1 U622 ( .A1(n587), .A2(n533), .ZN(n532) );
  OR2_X1 U623 ( .A1(n531), .A2(n533), .ZN(n534) );
  NOR2_X1 U624 ( .A1(n534), .A2(n608), .ZN(n536) );
  NAND2_X1 U625 ( .A1(n536), .A2(n535), .ZN(n537) );
  AND2_X1 U626 ( .A1(n638), .A2(n637), .ZN(n538) );
  NAND2_X1 U627 ( .A1(n539), .A2(n538), .ZN(n542) );
  NAND2_X1 U628 ( .A1(n654), .A2(KEYINPUT86), .ZN(n540) );
  NAND2_X1 U629 ( .A1(n542), .A2(n541), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n654), .A2(KEYINPUT44), .ZN(n544) );
  INV_X1 U631 ( .A(KEYINPUT86), .ZN(n543) );
  NAND2_X1 U632 ( .A1(n544), .A2(n543), .ZN(n565) );
  BUF_X1 U633 ( .A(n545), .Z(n546) );
  NAND2_X1 U634 ( .A1(n546), .A2(n587), .ZN(n688) );
  NOR2_X1 U635 ( .A1(n688), .A2(n551), .ZN(n548) );
  INV_X1 U636 ( .A(KEYINPUT31), .ZN(n547) );
  XNOR2_X1 U637 ( .A(n548), .B(n547), .ZN(n676) );
  INV_X1 U638 ( .A(n690), .ZN(n550) );
  OR2_X1 U639 ( .A1(n580), .A2(n550), .ZN(n591) );
  OR2_X1 U640 ( .A1(n591), .A2(n551), .ZN(n553) );
  INV_X1 U641 ( .A(KEYINPUT96), .ZN(n552) );
  XNOR2_X1 U642 ( .A(n553), .B(n552), .ZN(n555) );
  AND2_X1 U643 ( .A1(n555), .A2(n554), .ZN(n664) );
  OR2_X1 U644 ( .A1(n676), .A2(n664), .ZN(n558) );
  NOR2_X1 U645 ( .A1(n557), .A2(n556), .ZN(n675) );
  XOR2_X1 U646 ( .A(KEYINPUT102), .B(n675), .Z(n623) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n661) );
  NAND2_X1 U648 ( .A1(n623), .A2(n661), .ZN(n704) );
  NAND2_X1 U649 ( .A1(n558), .A2(n704), .ZN(n563) );
  NOR2_X1 U650 ( .A1(n608), .A2(n694), .ZN(n559) );
  NAND2_X1 U651 ( .A1(n560), .A2(n559), .ZN(n562) );
  INV_X1 U652 ( .A(KEYINPUT103), .ZN(n561) );
  XNOR2_X1 U653 ( .A(n562), .B(n561), .ZN(n765) );
  AND2_X1 U654 ( .A1(n563), .A2(n765), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X2 U656 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X2 U657 ( .A(n568), .B(KEYINPUT45), .ZN(n736) );
  NOR2_X1 U658 ( .A1(G900), .A2(n571), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n759), .A2(n572), .ZN(n573) );
  XNOR2_X1 U660 ( .A(KEYINPUT107), .B(n573), .ZN(n574) );
  NOR2_X1 U661 ( .A1(n575), .A2(n574), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n592), .A2(n693), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n694), .A2(n576), .ZN(n577) );
  XNOR2_X2 U664 ( .A(n577), .B(KEYINPUT69), .ZN(n609) );
  NAND2_X1 U665 ( .A1(n609), .A2(n587), .ZN(n579) );
  XOR2_X1 U666 ( .A(KEYINPUT109), .B(KEYINPUT28), .Z(n578) );
  XNOR2_X1 U667 ( .A(n579), .B(n578), .ZN(n581) );
  NOR2_X2 U668 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U669 ( .A(n582), .B(KEYINPUT110), .ZN(n606) );
  NAND2_X1 U670 ( .A1(n606), .A2(n583), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n669), .A2(n704), .ZN(n586) );
  INV_X1 U672 ( .A(KEYINPUT74), .ZN(n596) );
  NOR2_X1 U673 ( .A1(n596), .A2(KEYINPUT47), .ZN(n585) );
  INV_X1 U674 ( .A(n592), .ZN(n593) );
  NAND2_X1 U675 ( .A1(n594), .A2(n619), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n601), .A2(n595), .ZN(n635) );
  AND2_X1 U677 ( .A1(n596), .A2(KEYINPUT47), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n635), .A2(n597), .ZN(n598) );
  INV_X1 U679 ( .A(KEYINPUT75), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT38), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n619), .B(n600), .ZN(n603) );
  NOR2_X1 U682 ( .A1(n661), .A2(n624), .ZN(n602) );
  XNOR2_X1 U683 ( .A(n602), .B(KEYINPUT40), .ZN(n766) );
  INV_X1 U684 ( .A(n708), .ZN(n617) );
  INV_X1 U685 ( .A(n603), .ZN(n703) );
  NOR2_X1 U686 ( .A1(n617), .A2(n711), .ZN(n605) );
  XOR2_X1 U687 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n604) );
  XOR2_X1 U688 ( .A(n605), .B(n604), .Z(n720) );
  AND2_X1 U689 ( .A1(n606), .A2(n720), .ZN(n607) );
  XNOR2_X1 U690 ( .A(n607), .B(KEYINPUT42), .ZN(n767) );
  NAND2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U692 ( .A1(n661), .A2(n610), .ZN(n615) );
  XOR2_X1 U693 ( .A(KEYINPUT112), .B(n615), .Z(n612) );
  NOR2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U695 ( .A(n613), .B(KEYINPUT36), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n614), .A2(n689), .ZN(n681) );
  NAND2_X1 U697 ( .A1(n531), .A2(n615), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT43), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n639) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n683) );
  NAND2_X1 U702 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n655), .A2(G472), .ZN(n630) );
  XOR2_X1 U704 ( .A(KEYINPUT62), .B(n628), .Z(n629) );
  XNOR2_X1 U705 ( .A(n630), .B(n629), .ZN(n632) );
  INV_X1 U706 ( .A(G952), .ZN(n631) );
  INV_X1 U707 ( .A(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n634), .B(n633), .ZN(G57) );
  XNOR2_X1 U709 ( .A(n636), .B(n635), .ZN(G45) );
  XNOR2_X1 U710 ( .A(n637), .B(G119), .ZN(G21) );
  XNOR2_X1 U711 ( .A(n638), .B(G110), .ZN(G12) );
  XOR2_X1 U712 ( .A(G140), .B(n639), .Z(G42) );
  NAND2_X1 U713 ( .A1(n655), .A2(G210), .ZN(n644) );
  XNOR2_X1 U714 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n640) );
  XNOR2_X1 U715 ( .A(n640), .B(KEYINPUT55), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U717 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U719 ( .A(n647), .B(KEYINPUT59), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n651) );
  XOR2_X1 U722 ( .A(n651), .B(KEYINPUT65), .Z(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(G60) );
  XOR2_X1 U724 ( .A(G122), .B(n654), .Z(G24) );
  NAND2_X1 U725 ( .A1(n731), .A2(G469), .ZN(n659) );
  XNOR2_X1 U726 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n660), .A2(n735), .ZN(G54) );
  INV_X1 U730 ( .A(n661), .ZN(n673) );
  NAND2_X1 U731 ( .A1(n664), .A2(n673), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT114), .ZN(n663) );
  XNOR2_X1 U733 ( .A(G104), .B(n663), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n666) );
  NAND2_X1 U735 ( .A1(n664), .A2(n675), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U737 ( .A(G107), .B(KEYINPUT27), .Z(n667) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(G9) );
  XOR2_X1 U739 ( .A(G128), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U740 ( .A1(n669), .A2(n675), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G30) );
  NAND2_X1 U742 ( .A1(n673), .A2(n669), .ZN(n672) );
  XNOR2_X1 U743 ( .A(G146), .B(n672), .ZN(G48) );
  NAND2_X1 U744 ( .A1(n676), .A2(n673), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(G113), .ZN(G15) );
  XOR2_X1 U746 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n678) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U749 ( .A(G116), .B(n679), .ZN(G18) );
  XOR2_X1 U750 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(G125), .B(n682), .ZN(G27) );
  XOR2_X1 U753 ( .A(G134), .B(n683), .Z(G36) );
  NOR2_X1 U754 ( .A1(n684), .A2(KEYINPUT2), .ZN(n685) );
  XNOR2_X1 U755 ( .A(n685), .B(KEYINPUT82), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n726) );
  XOR2_X1 U757 ( .A(KEYINPUT121), .B(KEYINPUT52), .Z(n717) );
  INV_X1 U758 ( .A(n688), .ZN(n700) );
  NOR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n692) );
  XNOR2_X1 U760 ( .A(KEYINPUT119), .B(KEYINPUT50), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n692), .B(n691), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT49), .B(n695), .Z(n696) );
  NAND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U765 ( .A1(n587), .A2(n698), .ZN(n699) );
  NOR2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT51), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n702), .A2(n720), .ZN(n715) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n707) );
  INV_X1 U770 ( .A(n705), .ZN(n706) );
  NAND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U774 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  NAND2_X1 U775 ( .A1(n713), .A2(n721), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U777 ( .A(n717), .B(n716), .Z(n718) );
  NOR2_X1 U778 ( .A1(n719), .A2(n718), .ZN(n723) );
  AND2_X1 U779 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U781 ( .A1(n724), .A2(n754), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n727), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U784 ( .A1(n731), .A2(G478), .ZN(n729) );
  XNOR2_X1 U785 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U786 ( .A1(n735), .A2(n730), .ZN(G63) );
  NAND2_X1 U787 ( .A1(n731), .A2(G217), .ZN(n733) );
  XNOR2_X1 U788 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U789 ( .A1(n735), .A2(n734), .ZN(G66) );
  NOR2_X1 U790 ( .A1(n736), .A2(n759), .ZN(n741) );
  NAND2_X1 U791 ( .A1(n759), .A2(G224), .ZN(n737) );
  XOR2_X1 U792 ( .A(KEYINPUT61), .B(n737), .Z(n738) );
  NOR2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U794 ( .A1(n741), .A2(n740), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n742), .B(KEYINPUT123), .ZN(n744) );
  NAND2_X1 U796 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U797 ( .A(n745), .B(KEYINPUT124), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(G69) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(n748), .Z(n752) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n757) );
  XNOR2_X1 U802 ( .A(n753), .B(n757), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U804 ( .A(n756), .B(KEYINPUT126), .ZN(n762) );
  XNOR2_X1 U805 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U809 ( .A(KEYINPUT127), .B(n763), .Z(G72) );
  XOR2_X1 U810 ( .A(G101), .B(KEYINPUT113), .Z(n764) );
  XNOR2_X1 U811 ( .A(n765), .B(n764), .ZN(G3) );
  XOR2_X1 U812 ( .A(G131), .B(n766), .Z(G33) );
  XOR2_X1 U813 ( .A(G137), .B(n767), .Z(G39) );
endmodule

