//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n568, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n469), .A2(G2105), .B1(G101), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n465), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n463), .A3(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(new_n476), .A3(new_n466), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n477), .A2(new_n470), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n478), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n484), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  AND3_X1   g066(.A1(new_n474), .A2(new_n476), .A3(new_n466), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(G138), .A3(new_n470), .ZN(new_n493));
  INV_X1    g068(.A(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n493), .A2(KEYINPUT4), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n492), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n470), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT5), .B1(KEYINPUT70), .B2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT5), .A4(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(KEYINPUT73), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n510), .B2(KEYINPUT73), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI221_X4 g091(.A(KEYINPUT72), .B1(new_n515), .B2(new_n516), .C1(new_n507), .C2(new_n508), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n509), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n515), .B2(new_n516), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n522), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AND3_X1   g102(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(new_n524), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(new_n519), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT72), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n509), .A2(new_n518), .A3(new_n519), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n507), .A2(new_n508), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(G52), .B2(new_n524), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n536), .A2(G90), .A3(new_n537), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n543), .C2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n552), .B1(new_n507), .B2(new_n508), .ZN(new_n554));
  INV_X1    g129(.A(new_n551), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT74), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(G651), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n536), .A2(G81), .A3(new_n537), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT75), .B(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n524), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n557), .A2(KEYINPUT76), .A3(new_n558), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  AND3_X1   g147(.A1(new_n536), .A2(G91), .A3(new_n537), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G651), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n524), .A2(new_n576), .A3(G53), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n576), .B1(new_n524), .B2(G53), .ZN(new_n578));
  OAI22_X1  g153(.A1(new_n574), .A2(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n573), .A2(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n521), .A2(G87), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n509), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G49), .B2(new_n524), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n543), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n521), .A2(new_n589), .A3(G86), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n589), .B1(new_n521), .B2(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(G305));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(G47), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n538), .A2(new_n593), .B1(new_n594), .B2(new_n531), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI221_X1 g172(.A(KEYINPUT79), .B1(new_n594), .B2(new_n531), .C1(new_n538), .C2(new_n593), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n575), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n543), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(G54), .B2(new_n524), .ZN(new_n608));
  AOI21_X1  g183(.A(KEYINPUT10), .B1(new_n521), .B2(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  NOR4_X1   g186(.A1(new_n517), .A2(new_n520), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n608), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT80), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n604), .B1(new_n614), .B2(new_n603), .ZN(G321));
  XOR2_X1   g190(.A(G321), .B(KEYINPUT81), .Z(G284));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n573), .A2(new_n579), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(G868), .B2(new_n618), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n565), .A2(new_n603), .ZN(new_n623));
  INV_X1    g198(.A(new_n614), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n494), .A2(new_n472), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G123), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT82), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n486), .A2(G135), .ZN(new_n634));
  OR2_X1    g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n635), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n631), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT84), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(KEYINPUT14), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT86), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  INV_X1    g233(.A(G14), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT87), .ZN(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(KEYINPUT17), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n663), .B(new_n664), .C1(new_n442), .C2(new_n666), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n665), .A3(new_n663), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n680), .A3(KEYINPUT88), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n679), .A2(new_n680), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(new_n682), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n678), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT29), .Z(new_n701));
  INV_X1    g276(.A(G2090), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT91), .B(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G20), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT23), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n618), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1956), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n698), .A2(G26), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT28), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n482), .A2(G128), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n470), .A2(G116), .ZN(new_n714));
  OAI21_X1  g289(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n478), .B(KEYINPUT68), .ZN(new_n716));
  INV_X1    g291(.A(G140), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n713), .B1(new_n714), .B2(new_n715), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G2067), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n703), .A2(new_n704), .A3(new_n710), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G4), .A2(G16), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n614), .B2(G16), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT97), .B(G1348), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n705), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n566), .B2(new_n727), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(G1341), .Z(new_n730));
  AND3_X1   g305(.A1(new_n722), .A2(new_n726), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  NAND2_X1  g308(.A1(G115), .A2(G2104), .ZN(new_n734));
  INV_X1    g309(.A(G127), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n467), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n733), .B1(G2105), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G139), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n737), .B1(new_n716), .B2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT98), .Z(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  OR2_X1    g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G2072), .ZN(new_n743));
  NOR2_X1   g318(.A1(G168), .A2(new_n708), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n708), .B2(G21), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G171), .A2(new_n708), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G5), .B2(new_n708), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n698), .A2(G32), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT26), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n754), .A2(new_n755), .B1(G105), .B2(new_n472), .ZN(new_n756));
  INV_X1    g331(.A(G129), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n498), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n486), .B2(G141), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n751), .B1(new_n759), .B2(new_n698), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n749), .A2(new_n750), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n742), .A2(new_n743), .A3(new_n747), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n765), .B2(KEYINPUT24), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(KEYINPUT24), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n480), .B2(new_n698), .ZN(new_n768));
  INV_X1    g343(.A(G2084), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G28), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(KEYINPUT30), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n772), .B2(KEYINPUT30), .ZN(new_n775));
  NOR2_X1   g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n774), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n771), .A2(new_n779), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n770), .B(new_n780), .C1(new_n746), .C2(new_n745), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n698), .A2(G27), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n698), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT100), .B(G2078), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n786), .B(new_n787), .C1(new_n698), .C2(new_n637), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n749), .A2(new_n750), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n760), .A2(new_n762), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n781), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n764), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT101), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(G166), .A2(new_n727), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G22), .B2(new_n727), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT93), .B(G1971), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n708), .A2(G6), .ZN(new_n803));
  INV_X1    g378(.A(G305), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n708), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n801), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(G288), .A2(G16), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n708), .A2(G23), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(KEYINPUT92), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT33), .B(G1976), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n805), .A2(new_n806), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n808), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT34), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G1991), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n486), .A2(G131), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(new_n470), .B2(G107), .ZN(new_n824));
  OR3_X1    g399(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n482), .B2(G119), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G29), .ZN(new_n830));
  OR2_X1    g405(.A1(G25), .A2(G29), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(KEYINPUT90), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT90), .B1(new_n830), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n822), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  INV_X1    g411(.A(new_n822), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n837), .A3(new_n832), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  MUX2_X1   g414(.A(G24), .B(G290), .S(new_n727), .Z(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(G1986), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(G1986), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n808), .A2(new_n844), .A3(new_n817), .A4(new_n818), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n843), .A2(new_n845), .A3(KEYINPUT94), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT94), .B1(new_n843), .B2(new_n845), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n820), .B(new_n821), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n731), .B(new_n796), .C1(new_n848), .C2(KEYINPUT96), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n820), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n849), .B1(new_n851), .B2(new_n853), .ZN(G311));
  OR2_X1    g429(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n796), .A2(new_n731), .ZN(new_n856));
  INV_X1    g431(.A(new_n851), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n852), .ZN(G150));
  NAND2_X1  g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(G67), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n543), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G651), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n524), .A2(G55), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n862), .B(new_n863), .C1(new_n538), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n563), .B2(new_n564), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n561), .A2(new_n865), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n614), .A2(G559), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(new_n874), .A3(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n865), .A2(G860), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n877), .ZN(G145));
  OAI21_X1  g453(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n879));
  INV_X1    g454(.A(G118), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(G2105), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n482), .B2(G130), .ZN(new_n882));
  INV_X1    g457(.A(G142), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n716), .B2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT102), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n629), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n829), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n718), .B(G164), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(new_n740), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n740), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n759), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n759), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n637), .B(new_n480), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n490), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT103), .B1(new_n892), .B2(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n889), .A2(new_n890), .ZN(new_n899));
  INV_X1    g474(.A(new_n759), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n891), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n887), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT104), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n907), .B(new_n887), .C1(new_n898), .C2(new_n903), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n894), .B(new_n897), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n894), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n887), .A2(new_n892), .A3(new_n893), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n896), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT40), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT40), .B1(new_n909), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(G395));
  INV_X1    g492(.A(G288), .ZN(new_n918));
  XNOR2_X1  g493(.A(G303), .B(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n599), .A2(G305), .A3(new_n601), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G305), .B1(new_n599), .B2(new_n601), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G303), .B(G288), .ZN(new_n924));
  NAND2_X1  g499(.A1(G290), .A2(new_n804), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n927), .B(KEYINPUT42), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n625), .B(new_n869), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n613), .A2(G299), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n610), .B1(new_n538), .B2(new_n611), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n618), .B1(new_n933), .B2(new_n608), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n613), .A2(G299), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n618), .B(new_n608), .C1(new_n609), .C2(new_n612), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n937), .A2(KEYINPUT41), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT41), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n936), .B1(new_n942), .B2(new_n929), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n928), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n943), .A2(new_n944), .A3(new_n928), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g525(.A(new_n949), .B1(G868), .B2(new_n866), .ZN(G331));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n521), .A2(G81), .B1(new_n524), .B2(new_n559), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT76), .B1(new_n953), .B2(new_n557), .ZN(new_n954));
  INV_X1    g529(.A(new_n564), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n865), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n868), .ZN(new_n957));
  INV_X1    g532(.A(G90), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n517), .A2(new_n520), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n524), .A2(G52), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n961), .B2(new_n575), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT106), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n546), .A2(new_n964), .A3(new_n547), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G168), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n963), .A2(new_n965), .A3(G286), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n956), .A2(new_n957), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n963), .A2(new_n965), .A3(G286), .ZN(new_n970));
  AOI21_X1  g545(.A(G286), .B1(new_n963), .B2(new_n965), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n867), .A2(new_n868), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT41), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n930), .B2(new_n934), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT41), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n969), .A2(new_n972), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n941), .A2(KEYINPUT107), .A3(new_n969), .A4(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n969), .A2(new_n972), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n935), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n978), .A2(new_n979), .A3(new_n927), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n976), .A2(new_n977), .B1(new_n980), .B2(new_n935), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n985), .A2(KEYINPUT108), .A3(new_n927), .A4(new_n979), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n979), .ZN(new_n988));
  INV_X1    g563(.A(new_n927), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n981), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n980), .A2(KEYINPUT110), .A3(new_n935), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n941), .A2(new_n998), .A3(new_n969), .A4(new_n972), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(G37), .B1(new_n1000), .B2(new_n989), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n987), .A2(new_n1001), .A3(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n952), .B1(new_n993), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n987), .A2(new_n1001), .A3(new_n992), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT44), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT111), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1002), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT43), .B1(new_n987), .B2(new_n990), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1005), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n992), .B1(new_n987), .B2(new_n990), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n952), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1007), .A2(new_n1015), .ZN(G397));
  XNOR2_X1  g591(.A(new_n718), .B(new_n720), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n829), .A2(new_n822), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n759), .B(G1996), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n829), .A2(new_n822), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(G1986), .B2(G290), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n497), .B2(new_n502), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n1027), .B2(KEYINPUT112), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(KEYINPUT112), .B2(new_n1027), .ZN(new_n1029));
  INV_X1    g604(.A(G40), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n480), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G168), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1027), .A2(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1026), .C1(new_n497), .C2(new_n502), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1027), .A2(KEYINPUT50), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1042), .A2(new_n769), .A3(new_n1031), .A4(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT45), .B(new_n1026), .C1(new_n497), .C2(new_n502), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1031), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1044), .B1(new_n1049), .B2(G1966), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT122), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1044), .B(new_n1052), .C1(new_n1049), .C2(G1966), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1037), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(G168), .A3(new_n1053), .ZN(new_n1055));
  AND2_X1   g630(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1050), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n1037), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT62), .B(new_n1054), .C1(new_n1057), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2078), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1049), .A2(KEYINPUT53), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1042), .A2(new_n1031), .A3(new_n1043), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n750), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1027), .A2(new_n1048), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1031), .A3(new_n1045), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1068), .B2(G2078), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1063), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1073), .A3(G171), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G303), .A2(G8), .ZN(new_n1076));
  XNOR2_X1  g651(.A(new_n1076), .B(KEYINPUT55), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1971), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1068), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1064), .B2(G2090), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1081), .A3(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  INV_X1    g658(.A(G1981), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n521), .A2(G86), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n588), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT115), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1038), .A2(new_n1031), .A3(new_n1041), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n918), .A2(G1976), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT52), .ZN(new_n1097));
  INV_X1    g672(.A(G1976), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT52), .B1(G288), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1082), .A2(new_n1094), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1039), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1031), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1104), .A2(G2090), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1080), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1077), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1077), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT116), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1075), .A2(new_n1103), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT126), .B1(new_n1061), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1101), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n1115), .A3(new_n1082), .A4(new_n1110), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1070), .A2(new_n1073), .A3(G171), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1073), .B1(new_n1070), .B2(G171), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1054), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1120), .B(new_n1121), .C1(new_n1124), .C2(KEYINPUT62), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(KEYINPUT62), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1114), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1081), .A2(G8), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1115), .A2(new_n1078), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1083), .B1(new_n1094), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1092), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1050), .A2(G8), .A3(G168), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1116), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1133), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1103), .B(new_n1136), .C1(new_n1078), .C2(new_n1128), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1091), .A2(G2067), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT117), .ZN(new_n1140));
  INV_X1    g715(.A(G1348), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1064), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1956), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n618), .B(KEYINPUT57), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT56), .B(G2072), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1067), .A2(new_n1031), .A3(new_n1045), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1143), .A2(new_n614), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1146), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT58), .B(G1341), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1091), .A2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT118), .B(G1996), .Z(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1068), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n565), .A2(KEYINPUT119), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT59), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1153), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT60), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n614), .B2(KEYINPUT121), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1140), .A2(new_n1165), .A3(new_n1142), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n614), .A2(KEYINPUT121), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1166), .A2(new_n1167), .B1(new_n1143), .B2(new_n1164), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT61), .B1(new_n1153), .B2(new_n1149), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  AOI21_X1  g747(.A(new_n1154), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT53), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1046), .A2(new_n1174), .A3(G2078), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1029), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT125), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1178));
  AOI21_X1  g753(.A(G301), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT54), .B1(new_n1070), .B2(G171), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1116), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT54), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1177), .A2(G301), .A3(new_n1178), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1075), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1185), .A3(new_n1124), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1138), .B1(new_n1173), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1034), .B1(new_n1127), .B2(new_n1187), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n1029), .A2(G1996), .A3(new_n1032), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT46), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1033), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1017), .A2(new_n759), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(KEYINPUT127), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT47), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OR2_X1    g771(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1024), .A2(new_n1191), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1198), .A2(KEYINPUT48), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1021), .A2(new_n1033), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1198), .A2(KEYINPUT48), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1203), .A2(new_n1020), .B1(G2067), .B2(new_n718), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1033), .ZN(new_n1205));
  AND4_X1   g780(.A1(new_n1196), .A2(new_n1197), .A3(new_n1202), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1188), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g782(.A1(G227), .A2(new_n460), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n696), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n657), .B2(new_n660), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n894), .A2(new_n897), .ZN(new_n1212));
  NOR3_X1   g786(.A1(new_n892), .A2(KEYINPUT103), .A3(new_n893), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n902), .B1(new_n901), .B2(new_n891), .ZN(new_n1214));
  OAI21_X1  g788(.A(new_n905), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1215), .A2(new_n907), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n904), .A2(KEYINPUT104), .A3(new_n905), .ZN(new_n1217));
  AOI21_X1  g791(.A(new_n1212), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n912), .A2(new_n913), .ZN(new_n1219));
  OAI221_X1 g793(.A(new_n1211), .B1(new_n1011), .B2(new_n1012), .C1(new_n1218), .C2(new_n1219), .ZN(G225));
  INV_X1    g794(.A(G225), .ZN(G308));
endmodule


