//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n189), .B(new_n191), .C1(new_n192), .C2(KEYINPUT23), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(KEYINPUT16), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G140), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n196), .A2(new_n201), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n200), .B(new_n205), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n193), .A2(G110), .ZN(new_n209));
  AND3_X1   g023(.A1(new_n194), .A2(KEYINPUT74), .A3(new_n195), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT74), .B1(new_n194), .B2(new_n195), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G137), .ZN(new_n214));
  INV_X1    g028(.A(G953), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(G221), .A3(G234), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n214), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n207), .B(new_n217), .C1(new_n208), .C2(new_n212), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n187), .B1(new_n221), .B2(G902), .ZN(new_n222));
  INV_X1    g036(.A(G902), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n219), .A2(KEYINPUT25), .A3(new_n223), .A4(new_n220), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G234), .B2(new_n223), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n225), .B2(new_n228), .ZN(new_n231));
  NOR3_X1   g045(.A1(new_n221), .A2(G902), .A3(new_n228), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G472), .ZN(new_n234));
  NOR2_X1   g048(.A1(G237), .A2(G953), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G210), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n236), .B(KEYINPUT27), .Z(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT26), .B(G101), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT28), .ZN(new_n241));
  XOR2_X1   g055(.A(KEYINPUT2), .B(G113), .Z(new_n242));
  OR2_X1    g056(.A1(KEYINPUT70), .A2(G116), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT70), .A2(G116), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(G119), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n190), .A2(G116), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n242), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n242), .B1(new_n246), .B2(new_n245), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT64), .B1(new_n205), .B2(G143), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n254), .A2(new_n251), .A3(G146), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT0), .A3(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n205), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  OR2_X1    g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n260), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(KEYINPUT67), .A3(G137), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n267), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(G134), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n265), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT68), .B(G131), .C1(new_n272), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(G137), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n268), .A2(new_n277), .B1(new_n273), .B2(new_n265), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n266), .A2(G137), .ZN(new_n279));
  AND2_X1   g093(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n280));
  NOR2_X1   g094(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(KEYINPUT66), .B(G131), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n271), .A4(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G131), .B1(new_n272), .B2(new_n275), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n264), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n273), .A2(new_n277), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G131), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n256), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n260), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n292), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n250), .B1(new_n289), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n293), .ZN(new_n304));
  AOI21_X1  g118(.A(KEYINPUT69), .B1(new_n256), .B2(new_n293), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n292), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n257), .A2(new_n263), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n276), .A2(new_n284), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n282), .A2(new_n271), .A3(new_n267), .A4(new_n270), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT68), .B1(new_n311), .B2(G131), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n313), .A3(new_n249), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n241), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n288), .A2(new_n276), .A3(new_n284), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n316), .A2(new_n309), .B1(new_n306), .B2(new_n307), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT28), .B1(new_n317), .B2(new_n249), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n240), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT30), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n308), .A2(new_n313), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n308), .B2(new_n313), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n250), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n314), .A3(new_n239), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT29), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n314), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n249), .B1(new_n308), .B2(new_n313), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT28), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n239), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n303), .A2(new_n314), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n318), .B1(new_n333), .B2(KEYINPUT28), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n330), .B(new_n332), .C1(new_n334), .C2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n223), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n325), .B1(new_n336), .B2(KEYINPUT73), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n338), .A3(new_n223), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n234), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n318), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n240), .B1(new_n328), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n323), .A2(new_n314), .A3(new_n240), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT31), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n323), .A2(KEYINPUT31), .A3(new_n314), .A4(new_n240), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(G472), .A2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT30), .B1(new_n289), .B2(new_n302), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n308), .A2(new_n313), .A3(new_n320), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n326), .B1(new_n356), .B2(new_n250), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT31), .B1(new_n357), .B2(new_n240), .ZN(new_n358));
  INV_X1    g172(.A(new_n348), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n350), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n352), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n233), .B1(new_n340), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT9), .B(G234), .ZN(new_n365));
  OAI21_X1  g179(.A(G221), .B1(new_n365), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n368));
  INV_X1    g182(.A(new_n256), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n299), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n258), .A2(KEYINPUT78), .A3(KEYINPUT1), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(G128), .A3(new_n372), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n296), .A2(new_n297), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n375), .B2(G107), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G104), .ZN(new_n379));
  INV_X1    g193(.A(G101), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(G107), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n376), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT77), .B1(new_n375), .B2(G107), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n375), .B2(G107), .ZN(new_n386));
  OAI21_X1  g200(.A(G101), .B1(new_n381), .B2(KEYINPUT77), .ZN(new_n387));
  OAI22_X1  g201(.A1(new_n383), .A2(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n374), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n368), .B1(new_n389), .B2(KEYINPUT10), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n298), .B2(new_n301), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n386), .A2(new_n387), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n376), .A2(new_n379), .A3(new_n381), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT4), .B(new_n398), .C1(new_n383), .C2(new_n384), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n400), .A3(G101), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n257), .A2(new_n263), .A3(new_n401), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n392), .A2(new_n396), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n316), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n372), .A2(G128), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT78), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n369), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n304), .B2(new_n305), .ZN(new_n408));
  AOI21_X1  g222(.A(KEYINPUT10), .B1(new_n408), .B2(new_n396), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT79), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n390), .A2(new_n403), .A3(new_n404), .A4(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n316), .A2(KEYINPUT80), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n306), .A2(new_n396), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n389), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT12), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT12), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n412), .B(new_n416), .C1(new_n389), .C2(new_n413), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G140), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n215), .A2(G227), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n306), .A2(new_n396), .A3(KEYINPUT10), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n399), .A2(new_n402), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(new_n424), .C1(new_n409), .C2(KEYINPUT79), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n368), .B(KEYINPUT10), .C1(new_n408), .C2(new_n396), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n316), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n411), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n422), .A2(G469), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G469), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(new_n223), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AND4_X1   g248(.A1(new_n411), .A2(new_n415), .A3(new_n428), .A4(new_n417), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n428), .B1(new_n427), .B2(new_n411), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n431), .B(new_n223), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n367), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n283), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n235), .A2(G143), .A3(G214), .ZN(new_n440));
  AOI21_X1  g254(.A(G143), .B1(new_n235), .B2(G214), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n235), .A2(G214), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n251), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n235), .A2(G143), .A3(G214), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n283), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n442), .A2(new_n446), .B1(new_n200), .B2(G146), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT19), .B1(new_n199), .B2(KEYINPUT84), .ZN(new_n448));
  AND4_X1   g262(.A1(KEYINPUT84), .A2(new_n203), .A3(new_n204), .A4(KEYINPUT19), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n205), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n206), .A2(KEYINPUT83), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n203), .A2(new_n204), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G146), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(KEYINPUT83), .A3(G146), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n444), .A2(KEYINPUT18), .A3(G131), .A4(new_n445), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT18), .A2(G131), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n440), .B2(new_n441), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n447), .A2(new_n450), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n375), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT85), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n442), .A2(new_n446), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n450), .A3(new_n201), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n456), .A2(new_n460), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n469));
  INV_X1    g283(.A(new_n463), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n200), .A2(G146), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n439), .B(KEYINPUT17), .C1(new_n440), .C2(new_n441), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n201), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n465), .A2(KEYINPUT17), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n463), .B(new_n467), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n464), .A2(new_n471), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(G475), .A2(G902), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(KEYINPUT86), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT20), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT86), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n478), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n208), .B(new_n473), .C1(KEYINPUT17), .C2(new_n465), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n463), .B1(new_n487), .B2(new_n467), .ZN(new_n488));
  INV_X1    g302(.A(new_n476), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n223), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G475), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G952), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(KEYINPUT87), .ZN(new_n496));
  AOI21_X1  g310(.A(G953), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(G234), .A2(G237), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT88), .Z(new_n500));
  AND3_X1   g314(.A1(new_n498), .A2(G902), .A3(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT21), .B(G898), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G128), .B(G143), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(new_n266), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n243), .A2(G122), .A3(new_n244), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n378), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n508), .A2(new_n512), .A3(new_n510), .ZN(new_n513));
  OAI21_X1  g327(.A(G107), .B1(new_n508), .B2(new_n512), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n507), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n506), .A2(KEYINPUT13), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n188), .A2(KEYINPUT13), .A3(G143), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n266), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n516), .A2(new_n518), .B1(new_n266), .B2(new_n506), .ZN(new_n519));
  INV_X1    g333(.A(new_n511), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n378), .B1(new_n508), .B2(new_n510), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n365), .A2(new_n227), .A3(G953), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n522), .A3(new_n524), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G478), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n528), .B(new_n223), .C1(KEYINPUT15), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI211_X1 g345(.A(KEYINPUT15), .B(new_n529), .C1(new_n528), .C2(new_n223), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n493), .A2(KEYINPUT89), .A3(new_n505), .A4(new_n533), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT86), .B(KEYINPUT20), .C1(new_n477), .C2(new_n478), .ZN(new_n535));
  INV_X1    g349(.A(G475), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n487), .A2(new_n467), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n470), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n476), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n223), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n483), .A2(new_n484), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT20), .A3(new_n479), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n541), .A2(new_n505), .A3(new_n543), .A4(new_n533), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT89), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n534), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G214), .B1(G237), .B2(G902), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT81), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n401), .B1(new_n247), .B2(new_n248), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n394), .A2(new_n395), .ZN(new_n553));
  INV_X1    g367(.A(new_n398), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(new_n400), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n247), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n245), .A2(KEYINPUT5), .A3(new_n246), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n559));
  INV_X1    g373(.A(G113), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n388), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n551), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n552), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n399), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n247), .B1(new_n558), .B2(new_n561), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n396), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n550), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT6), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT6), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n572), .B(new_n551), .C1(new_n556), .C2(new_n564), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n197), .B1(new_n257), .B2(new_n263), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n296), .A2(new_n297), .B1(new_n260), .B2(new_n300), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n197), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n215), .A2(G224), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n574), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n306), .B2(G125), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(G224), .A3(new_n215), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n573), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n388), .A2(new_n563), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n569), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n550), .B(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n577), .A2(KEYINPUT7), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n585), .A2(new_n586), .B1(new_n576), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n566), .A2(new_n399), .B1(new_n396), .B2(new_n568), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n590), .A2(new_n550), .B1(new_n580), .B2(new_n587), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n583), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n583), .B2(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n548), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT82), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n548), .C1(new_n594), .C2(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n438), .A2(new_n547), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n364), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT90), .B(G101), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  NAND3_X1  g418(.A1(new_n437), .A2(new_n433), .A3(new_n430), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n366), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n349), .B2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n361), .ZN(new_n608));
  INV_X1    g422(.A(new_n233), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n592), .ZN(new_n611));
  INV_X1    g425(.A(new_n593), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT91), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n583), .A2(new_n592), .A3(new_n593), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n548), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n595), .B2(KEYINPUT91), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT92), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n620), .A2(KEYINPUT92), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n528), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n620), .A4(new_n527), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n223), .A2(G478), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n526), .B2(new_n527), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT93), .B(G478), .ZN(new_n629));
  OAI22_X1  g443(.A1(new_n626), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n630), .B(new_n505), .C1(new_n482), .C2(new_n492), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n619), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n610), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT94), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT34), .B(G104), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G6));
  INV_X1    g450(.A(new_n533), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n637), .A2(new_n541), .A3(new_n505), .A4(new_n543), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n610), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NAND2_X1  g456(.A1(new_n225), .A2(new_n228), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT75), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n218), .A2(KEYINPUT36), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n213), .B(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n646), .B(new_n223), .C1(new_n227), .C2(G234), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n229), .A3(new_n647), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n607), .A2(new_n361), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n547), .A3(new_n438), .A4(new_n600), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  INV_X1    g466(.A(new_n619), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n653), .B(new_n648), .C1(new_n340), .C2(new_n363), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n541), .A2(new_n543), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n533), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n501), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n500), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT95), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n656), .A2(KEYINPUT95), .A3(new_n660), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n438), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n654), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n188), .ZN(G30));
  XOR2_X1   g481(.A(new_n659), .B(KEYINPUT39), .Z(new_n668));
  AND2_X1   g482(.A1(new_n438), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT40), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n349), .A2(new_n362), .A3(new_n351), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n361), .B2(new_n342), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n357), .A2(new_n239), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n223), .B1(new_n333), .B2(new_n240), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n594), .A2(new_n595), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n655), .A2(new_n637), .ZN(new_n679));
  NOR4_X1   g493(.A1(new_n678), .A2(new_n617), .A3(new_n648), .A4(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n670), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  NAND2_X1  g496(.A1(new_n655), .A2(new_n630), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n438), .A2(new_n684), .A3(new_n660), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n654), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(new_n205), .ZN(G48));
  NAND2_X1  g501(.A1(new_n337), .A2(new_n339), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G472), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n609), .B1(new_n689), .B2(new_n672), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n223), .B1(new_n435), .B2(new_n436), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(G469), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n366), .A3(new_n437), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT96), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n692), .A2(KEYINPUT96), .A3(new_n366), .A4(new_n437), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n690), .A2(new_n697), .A3(new_n632), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND3_X1  g514(.A1(new_n690), .A2(new_n697), .A3(new_n639), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  OAI21_X1  g516(.A(new_n648), .B1(new_n340), .B2(new_n363), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n693), .A2(new_n619), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n547), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n190), .ZN(G21));
  OAI21_X1  g521(.A(new_n330), .B1(new_n334), .B2(new_n329), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n239), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n347), .A2(new_n348), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n351), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT97), .B(G472), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n349), .B2(G902), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT98), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(KEYINPUT98), .B(new_n712), .C1(new_n349), .C2(G902), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n711), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n233), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n619), .A2(new_n679), .A3(new_n504), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n695), .A3(new_n696), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n509), .ZN(G24));
  NAND3_X1  g536(.A1(new_n704), .A2(new_n684), .A3(new_n660), .ZN(new_n723));
  INV_X1    g537(.A(new_n711), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n360), .A2(new_n223), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT98), .B1(new_n725), .B2(new_n712), .ZN(new_n726));
  INV_X1    g540(.A(new_n716), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n648), .B(new_n724), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT99), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n717), .A2(KEYINPUT99), .A3(new_n648), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n197), .ZN(G27));
  XNOR2_X1  g547(.A(new_n361), .B(new_n362), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n233), .B1(new_n734), .B2(new_n340), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n655), .A2(new_n630), .A3(new_n660), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n677), .A2(new_n548), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n606), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n690), .A2(KEYINPUT100), .A3(new_n739), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT100), .ZN(new_n744));
  INV_X1    g558(.A(new_n738), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n438), .A2(new_n684), .A3(new_n660), .A4(new_n745), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n364), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n740), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G131), .ZN(G33));
  OAI211_X1 g564(.A(new_n233), .B(new_n745), .C1(new_n340), .C2(new_n363), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n665), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n266), .ZN(G36));
  NAND2_X1  g567(.A1(new_n493), .A2(new_n630), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n608), .A3(new_n648), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT103), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  XOR2_X1   g575(.A(new_n761), .B(KEYINPUT104), .Z(new_n762));
  NOR3_X1   g576(.A1(new_n760), .A2(new_n762), .A3(new_n738), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n422), .A2(KEYINPUT45), .A3(new_n429), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT45), .B1(new_n422), .B2(new_n429), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n431), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n432), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n767), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT101), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n768), .A2(new_n437), .A3(new_n769), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n366), .A3(new_n668), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT102), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(KEYINPUT102), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n763), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NAND2_X1  g590(.A1(new_n771), .A2(new_n366), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n771), .A2(new_n366), .A3(new_n778), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n745), .A2(new_n609), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n783), .A2(new_n340), .A3(new_n363), .A4(new_n737), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT106), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  OAI22_X1  g601(.A1(new_n718), .A2(new_n720), .B1(new_n703), .B2(new_n705), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n605), .A2(new_n233), .A3(new_n366), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n597), .A2(new_n599), .B1(new_n631), .B2(new_n638), .ZN(new_n790));
  INV_X1    g604(.A(new_n608), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n650), .B(new_n792), .C1(new_n364), .C2(new_n601), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n690), .B(new_n697), .C1(new_n632), .C2(new_n639), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n730), .A2(new_n731), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n739), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n655), .A2(new_n637), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n438), .A2(new_n798), .A3(new_n660), .A4(new_n745), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n703), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n752), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n795), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n735), .A2(new_n742), .A3(new_n746), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n364), .A2(new_n746), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT42), .B1(new_n804), .B2(KEYINPUT100), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n805), .B2(new_n747), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT109), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n795), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n808), .A2(new_n793), .A3(new_n788), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n746), .B1(new_n730), .B2(new_n731), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n810), .A2(new_n752), .A3(new_n800), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(new_n749), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n654), .B1(new_n665), .B2(new_n685), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n732), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  OR3_X1    g631(.A1(new_n648), .A2(new_n817), .A3(new_n659), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n648), .B2(new_n659), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n619), .A2(new_n679), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n676), .A2(new_n820), .A3(new_n438), .A4(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT112), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(KEYINPUT112), .A3(new_n822), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(new_n822), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n732), .A2(new_n828), .A3(new_n815), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n814), .A2(new_n826), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n802), .A2(new_n806), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n816), .A2(new_n822), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n831), .A2(KEYINPUT53), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n807), .A2(KEYINPUT110), .A3(new_n813), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT110), .B1(new_n807), .B2(new_n813), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n837), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI22_X1  g658(.A1(new_n844), .A2(KEYINPUT53), .B1(new_n832), .B2(new_n833), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(KEYINPUT54), .B2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n500), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n756), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n693), .A2(new_n738), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n736), .ZN(new_n851));
  XOR2_X1   g665(.A(new_n851), .B(KEYINPUT48), .Z(new_n852));
  XOR2_X1   g666(.A(new_n497), .B(KEYINPUT119), .Z(new_n853));
  INV_X1    g667(.A(new_n676), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n233), .A3(new_n847), .A4(new_n849), .ZN(new_n855));
  INV_X1    g669(.A(new_n704), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n848), .A2(new_n233), .A3(new_n717), .ZN(new_n857));
  OAI221_X1 g671(.A(new_n853), .B1(new_n855), .B2(new_n683), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n855), .A2(new_n655), .A3(new_n630), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n692), .A2(new_n437), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT114), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n367), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n780), .A2(new_n781), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n857), .A2(new_n738), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n859), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n678), .A2(new_n617), .ZN(new_n868));
  OR3_X1    g682(.A1(new_n857), .A2(new_n693), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT50), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n869), .B2(KEYINPUT115), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n850), .A2(new_n796), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT117), .Z(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n867), .A2(new_n874), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT118), .B1(new_n865), .B2(new_n866), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(KEYINPUT51), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n852), .B(new_n858), .C1(new_n879), .C2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n846), .B(new_n882), .C1(new_n881), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n494), .A2(new_n215), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n609), .A2(new_n754), .A3(new_n367), .A4(new_n617), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT49), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n861), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT107), .Z(new_n889));
  OAI21_X1  g703(.A(new_n678), .B1(KEYINPUT49), .B2(new_n860), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n676), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n885), .A2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n215), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n838), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n832), .B2(new_n833), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n223), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n571), .A2(new_n573), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n582), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n895), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n899), .B2(new_n902), .ZN(G51));
  XNOR2_X1  g718(.A(new_n432), .B(KEYINPUT57), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n834), .B2(new_n838), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n840), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n435), .A2(new_n436), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT120), .B(new_n905), .C1(new_n840), .C2(new_n907), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n898), .A2(new_n766), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n894), .B1(new_n913), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n898), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  INV_X1    g730(.A(new_n477), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n918), .A2(new_n919), .A3(new_n894), .ZN(G60));
  NAND2_X1  g734(.A1(G478), .A2(G902), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT59), .Z(new_n922));
  OR2_X1    g736(.A1(new_n626), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n897), .A2(new_n906), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n894), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT121), .B1(new_n926), .B2(new_n894), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n626), .B1(new_n846), .B2(new_n922), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n221), .B1(new_n897), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n932), .ZN(new_n934));
  INV_X1    g748(.A(new_n833), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n823), .A2(new_n830), .ZN(new_n936));
  AOI22_X1  g750(.A1(KEYINPUT52), .A2(new_n936), .B1(new_n807), .B2(new_n813), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n831), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n646), .B(new_n934), .C1(new_n938), .C2(new_n896), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n895), .A4(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n895), .A4(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n839), .A2(new_n947), .A3(new_n646), .A4(new_n934), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n946), .A2(new_n895), .A3(new_n933), .A4(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n949), .A2(KEYINPUT123), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT123), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n502), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n809), .B2(G953), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n900), .B1(G898), .B2(new_n215), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n681), .A2(new_n816), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT62), .Z(new_n960));
  INV_X1    g774(.A(new_n751), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n669), .C1(new_n684), .C2(new_n656), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n786), .A2(new_n775), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n215), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n448), .A2(new_n449), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n356), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n773), .A2(new_n821), .A3(new_n736), .A4(new_n774), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n775), .A2(new_n816), .A3(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n806), .A2(new_n752), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n786), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n968), .B1(new_n973), .B2(G953), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n215), .B1(G227), .B2(G900), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n976), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n975), .B(new_n978), .ZN(G72));
  XOR2_X1   g793(.A(new_n324), .B(KEYINPUT127), .Z(new_n980));
  INV_X1    g794(.A(new_n673), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n973), .A2(new_n980), .B1(new_n963), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n809), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n981), .ZN(new_n984));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT63), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n894), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n324), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n673), .A2(new_n989), .A3(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n988), .B1(new_n845), .B2(new_n990), .ZN(G57));
endmodule


