

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  BUF_X2 U321 ( .A(n560), .Z(n289) );
  BUF_X1 U322 ( .A(n555), .Z(n290) );
  XOR2_X1 U323 ( .A(n346), .B(n345), .Z(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n358) );
  XNOR2_X1 U325 ( .A(n359), .B(n358), .ZN(n376) );
  XNOR2_X1 U326 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U327 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n387) );
  XNOR2_X1 U328 ( .A(n357), .B(n356), .ZN(n380) );
  XNOR2_X1 U329 ( .A(n388), .B(n387), .ZN(n540) );
  XOR2_X1 U330 ( .A(n405), .B(n404), .Z(n511) );
  XNOR2_X1 U331 ( .A(n449), .B(KEYINPUT124), .ZN(n450) );
  XNOR2_X1 U332 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT64), .B(KEYINPUT73), .Z(n293) );
  XNOR2_X1 U334 ( .A(G92GAT), .B(KEYINPUT78), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U336 ( .A(KEYINPUT76), .B(KEYINPUT10), .Z(n295) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(G162GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U339 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U340 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n299) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U343 ( .A(KEYINPUT11), .B(n300), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT70), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n351) );
  XNOR2_X1 U349 ( .A(G218GAT), .B(n351), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U351 ( .A(n308), .B(n307), .Z(n314) );
  XNOR2_X1 U352 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n309), .B(G29GAT), .ZN(n310) );
  XOR2_X1 U354 ( .A(n310), .B(KEYINPUT7), .Z(n312) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G50GAT), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n312), .B(n311), .ZN(n342) );
  XNOR2_X1 U357 ( .A(n342), .B(G134GAT), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n536) );
  INV_X1 U359 ( .A(n536), .ZN(n548) );
  XOR2_X1 U360 ( .A(G120GAT), .B(G71GAT), .Z(n344) );
  XOR2_X1 U361 ( .A(G99GAT), .B(G15GAT), .Z(n316) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G43GAT), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U364 ( .A(n344), .B(n317), .Z(n319) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U367 ( .A(KEYINPUT80), .B(KEYINPUT82), .Z(n321) );
  XNOR2_X1 U368 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U370 ( .A(n323), .B(n322), .Z(n332) );
  XNOR2_X1 U371 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n324), .B(KEYINPUT81), .ZN(n325) );
  XOR2_X1 U373 ( .A(n325), .B(KEYINPUT18), .Z(n327) );
  XNOR2_X1 U374 ( .A(G183GAT), .B(G190GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n400) );
  XOR2_X1 U376 ( .A(KEYINPUT79), .B(G134GAT), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U379 ( .A(G113GAT), .B(n330), .Z(n422) );
  XNOR2_X1 U380 ( .A(n400), .B(n422), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n522) );
  XOR2_X1 U382 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n334) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U385 ( .A(n335), .B(KEYINPUT66), .Z(n337) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n431) );
  XOR2_X1 U387 ( .A(G169GAT), .B(G8GAT), .Z(n392) );
  XNOR2_X1 U388 ( .A(n431), .B(n392), .ZN(n336) );
  XNOR2_X1 U389 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U390 ( .A(G15GAT), .B(G1GAT), .Z(n371) );
  XOR2_X1 U391 ( .A(n338), .B(n371), .Z(n340) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G113GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n565) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n343), .B(G64GAT), .ZN(n396) );
  XOR2_X1 U397 ( .A(n396), .B(n344), .Z(n346) );
  NAND2_X1 U398 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XOR2_X1 U399 ( .A(G57GAT), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U400 ( .A(n291), .B(n360), .ZN(n348) );
  XNOR2_X1 U401 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n357) );
  XOR2_X1 U403 ( .A(G78GAT), .B(G148GAT), .Z(n350) );
  XNOR2_X1 U404 ( .A(KEYINPUT69), .B(G204GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n436) );
  XOR2_X1 U406 ( .A(n436), .B(n351), .Z(n355) );
  XOR2_X1 U407 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n353) );
  XNOR2_X1 U408 ( .A(KEYINPUT68), .B(KEYINPUT31), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n380), .B(KEYINPUT41), .Z(n555) );
  NAND2_X1 U411 ( .A1(n565), .A2(n290), .ZN(n359) );
  XNOR2_X1 U412 ( .A(G22GAT), .B(G211GAT), .ZN(n361) );
  XOR2_X1 U413 ( .A(n361), .B(n360), .Z(n375) );
  XOR2_X1 U414 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n363) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U417 ( .A(KEYINPUT14), .B(G64GAT), .Z(n365) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(G127GAT), .ZN(n364) );
  XNOR2_X1 U419 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U420 ( .A(n367), .B(n366), .Z(n373) );
  XOR2_X1 U421 ( .A(G78GAT), .B(G155GAT), .Z(n369) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n573) );
  NOR2_X1 U427 ( .A1(n376), .A2(n573), .ZN(n377) );
  AND2_X1 U428 ( .A1(n536), .A2(n377), .ZN(n379) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n379), .B(n378), .ZN(n386) );
  BUF_X1 U431 ( .A(n380), .Z(n570) );
  XOR2_X1 U432 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT36), .B(n536), .Z(n575) );
  NAND2_X1 U434 ( .A1(n573), .A2(n575), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U436 ( .A(KEYINPUT67), .B(n565), .ZN(n552) );
  NAND2_X1 U437 ( .A1(n383), .A2(n552), .ZN(n384) );
  NOR2_X1 U438 ( .A1(n570), .A2(n384), .ZN(n385) );
  NOR2_X1 U439 ( .A1(n386), .A2(n385), .ZN(n388) );
  XOR2_X1 U440 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n390) );
  XNOR2_X1 U441 ( .A(G36GAT), .B(G204GAT), .ZN(n389) );
  XNOR2_X1 U442 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U443 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U446 ( .A(n395), .B(KEYINPUT90), .Z(n398) );
  XNOR2_X1 U447 ( .A(n396), .B(KEYINPUT91), .ZN(n397) );
  XNOR2_X1 U448 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U449 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U450 ( .A(KEYINPUT21), .B(G218GAT), .Z(n402) );
  XNOR2_X1 U451 ( .A(KEYINPUT85), .B(G211GAT), .ZN(n401) );
  XNOR2_X1 U452 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U453 ( .A(G197GAT), .B(n403), .Z(n439) );
  INV_X1 U454 ( .A(n439), .ZN(n404) );
  INV_X1 U455 ( .A(n511), .ZN(n406) );
  NAND2_X1 U456 ( .A1(n540), .A2(n406), .ZN(n408) );
  XOR2_X1 U457 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n407) );
  XNOR2_X1 U458 ( .A(n408), .B(n407), .ZN(n427) );
  XOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n410) );
  XNOR2_X1 U460 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n426) );
  XOR2_X1 U462 ( .A(G85GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G141GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U465 ( .A(G57GAT), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G120GAT), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U468 ( .A(n416), .B(n415), .Z(n424) );
  XOR2_X1 U469 ( .A(G155GAT), .B(KEYINPUT2), .Z(n418) );
  XNOR2_X1 U470 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n438) );
  XOR2_X1 U472 ( .A(n438), .B(KEYINPUT5), .Z(n420) );
  NAND2_X1 U473 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U477 ( .A(n426), .B(n425), .Z(n508) );
  NAND2_X1 U478 ( .A1(n427), .A2(n508), .ZN(n564) );
  XOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n429) );
  XNOR2_X1 U480 ( .A(G50GAT), .B(G106GAT), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U482 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n443) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n435) );
  XNOR2_X1 U486 ( .A(KEYINPUT23), .B(KEYINPUT84), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U488 ( .A(n437), .B(n436), .Z(n441) );
  XNOR2_X1 U489 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U490 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U491 ( .A(n443), .B(n442), .ZN(n457) );
  NOR2_X1 U492 ( .A1(n564), .A2(n457), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n444), .B(KEYINPUT55), .ZN(n445) );
  NOR2_X1 U494 ( .A1(n522), .A2(n445), .ZN(n446) );
  XOR2_X1 U495 ( .A(KEYINPUT121), .B(n446), .Z(n560) );
  NAND2_X1 U496 ( .A1(n548), .A2(n289), .ZN(n451) );
  XOR2_X1 U497 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n448) );
  XNOR2_X1 U498 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  NOR2_X1 U500 ( .A1(n552), .A2(n570), .ZN(n482) );
  XNOR2_X1 U501 ( .A(KEYINPUT27), .B(n511), .ZN(n460) );
  NOR2_X1 U502 ( .A1(n508), .A2(n460), .ZN(n539) );
  XNOR2_X1 U503 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n452), .B(n457), .ZN(n517) );
  NAND2_X1 U505 ( .A1(n539), .A2(n517), .ZN(n521) );
  XNOR2_X1 U506 ( .A(n521), .B(KEYINPUT93), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n453), .A2(n522), .ZN(n466) );
  XOR2_X1 U508 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n456) );
  NOR2_X1 U509 ( .A1(n522), .A2(n511), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n457), .A2(n454), .ZN(n455) );
  XNOR2_X1 U511 ( .A(n456), .B(n455), .ZN(n462) );
  XOR2_X1 U512 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n459) );
  NAND2_X1 U513 ( .A1(n522), .A2(n457), .ZN(n458) );
  XOR2_X1 U514 ( .A(n459), .B(n458), .Z(n563) );
  OR2_X1 U515 ( .A1(n563), .A2(n460), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U517 ( .A(KEYINPUT96), .B(n463), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n464), .A2(n508), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n478) );
  NAND2_X1 U520 ( .A1(n536), .A2(n573), .ZN(n467) );
  XOR2_X1 U521 ( .A(KEYINPUT16), .B(n467), .Z(n468) );
  AND2_X1 U522 ( .A1(n478), .A2(n468), .ZN(n496) );
  NAND2_X1 U523 ( .A1(n482), .A2(n496), .ZN(n475) );
  NOR2_X1 U524 ( .A1(n508), .A2(n475), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT34), .B(n469), .Z(n470) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(n470), .ZN(G1324GAT) );
  NOR2_X1 U527 ( .A1(n511), .A2(n475), .ZN(n472) );
  XNOR2_X1 U528 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(G1325GAT) );
  NOR2_X1 U530 ( .A1(n522), .A2(n475), .ZN(n474) );
  XNOR2_X1 U531 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U533 ( .A1(n517), .A2(n475), .ZN(n476) );
  XOR2_X1 U534 ( .A(KEYINPUT98), .B(n476), .Z(n477) );
  XNOR2_X1 U535 ( .A(G22GAT), .B(n477), .ZN(G1327GAT) );
  INV_X1 U536 ( .A(n573), .ZN(n531) );
  NAND2_X1 U537 ( .A1(n531), .A2(n478), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT99), .B(n479), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n480), .A2(n575), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n481), .ZN(n507) );
  NAND2_X1 U541 ( .A1(n507), .A2(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n491) );
  NOR2_X1 U544 ( .A1(n508), .A2(n491), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT39), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U547 ( .A(G29GAT), .B(n487), .Z(G1328GAT) );
  NOR2_X1 U548 ( .A1(n511), .A2(n491), .ZN(n488) );
  XOR2_X1 U549 ( .A(G36GAT), .B(n488), .Z(G1329GAT) );
  NOR2_X1 U550 ( .A1(n522), .A2(n491), .ZN(n489) );
  XOR2_X1 U551 ( .A(KEYINPUT40), .B(n489), .Z(n490) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  NOR2_X1 U553 ( .A1(n517), .A2(n491), .ZN(n493) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  INV_X1 U557 ( .A(n290), .ZN(n527) );
  NOR2_X1 U558 ( .A1(n527), .A2(n565), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n495), .B(KEYINPUT104), .ZN(n506) );
  NAND2_X1 U560 ( .A1(n496), .A2(n506), .ZN(n503) );
  NOR2_X1 U561 ( .A1(n508), .A2(n503), .ZN(n497) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n497), .Z(n498) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(n498), .ZN(G1332GAT) );
  NOR2_X1 U564 ( .A1(n511), .A2(n503), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n499) );
  XNOR2_X1 U566 ( .A(n500), .B(n499), .ZN(G1333GAT) );
  NOR2_X1 U567 ( .A1(n522), .A2(n503), .ZN(n501) );
  XOR2_X1 U568 ( .A(KEYINPUT106), .B(n501), .Z(n502) );
  XNOR2_X1 U569 ( .A(G71GAT), .B(n502), .ZN(G1334GAT) );
  NOR2_X1 U570 ( .A1(n517), .A2(n503), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n506), .ZN(n516) );
  NOR2_X1 U574 ( .A1(n508), .A2(n516), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1336GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n516), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(n514), .ZN(G1337GAT) );
  NOR2_X1 U581 ( .A1(n522), .A2(n516), .ZN(n515) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n515), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n519) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n520), .Z(G1339GAT) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U588 ( .A1(n540), .A2(n523), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n552), .A2(n535), .ZN(n525) );
  XNOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n526), .ZN(G1340GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n535), .ZN(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n535), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n538) );
  XNOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U605 ( .A1(n563), .A2(n541), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n565), .A2(n549), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n544) );
  NAND2_X1 U610 ( .A1(n549), .A2(n290), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n549), .A2(n573), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U615 ( .A(G162GAT), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  INV_X1 U618 ( .A(n552), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n289), .A2(n553), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n554), .ZN(G1348GAT) );
  NAND2_X1 U621 ( .A1(n289), .A2(n290), .ZN(n557) );
  XOR2_X1 U622 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT123), .Z(n562) );
  NAND2_X1 U627 ( .A1(n289), .A2(n573), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .Z(n567) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  NAND2_X1 U631 ( .A1(n576), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT59), .B(KEYINPUT127), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n576), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT62), .ZN(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

