//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT65), .B1(new_n187), .B2(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT64), .A2(G146), .ZN(new_n190));
  NOR2_X1   g004(.A1(KEYINPUT64), .A2(G146), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n189), .B1(new_n192), .B2(G143), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n194), .B(new_n187), .C1(new_n190), .C2(new_n191), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n192), .B2(G143), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT68), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT68), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n193), .B(new_n195), .C1(new_n197), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT64), .A2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G143), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n187), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n201), .A2(new_n202), .A3(new_n211), .ZN(new_n212));
  XOR2_X1   g026(.A(KEYINPUT0), .B(G128), .Z(new_n213));
  AOI21_X1  g027(.A(G143), .B1(new_n205), .B2(new_n206), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n195), .B(new_n213), .C1(new_n214), .C2(new_n188), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n207), .A2(KEYINPUT0), .A3(G128), .A4(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT90), .B(G224), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT91), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n220), .A2(new_n221), .A3(G953), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n221), .B1(new_n220), .B2(G953), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT92), .B(KEYINPUT7), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT93), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n230), .A3(new_n224), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n231), .A2(KEYINPUT7), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT93), .B1(new_n223), .B2(new_n225), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n232), .A2(new_n218), .A3(new_n212), .A4(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT8), .ZN(new_n236));
  INV_X1    g050(.A(G101), .ZN(new_n237));
  INV_X1    g051(.A(G107), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G104), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n238), .A2(KEYINPUT85), .A3(G104), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n238), .A2(KEYINPUT85), .A3(KEYINPUT3), .A4(G104), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n241), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G101), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n242), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G116), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(G119), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT5), .ZN(new_n259));
  XNOR2_X1  g073(.A(G116), .B(G119), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n255), .A2(new_n259), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n250), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n250), .A2(new_n265), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n236), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n229), .A2(new_n234), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n247), .A2(new_n249), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n248), .B1(new_n245), .B2(new_n246), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n271), .B(KEYINPUT4), .C1(new_n237), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n260), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT2), .B(G113), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n264), .A2(new_n260), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT69), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  INV_X1    g093(.A(new_n277), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n264), .A2(new_n260), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n240), .A2(G107), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT3), .B1(new_n283), .B2(KEYINPUT85), .ZN(new_n284));
  INV_X1    g098(.A(new_n246), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n241), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G101), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n273), .A2(new_n278), .A3(new_n282), .A4(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT88), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n266), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n250), .A2(KEYINPUT88), .A3(new_n265), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .A4(new_n235), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n270), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n235), .A2(KEYINPUT6), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n250), .A2(KEYINPUT88), .A3(new_n265), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT88), .B1(new_n250), .B2(new_n265), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g113(.A(KEYINPUT89), .B(new_n296), .C1(new_n299), .C2(new_n289), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT89), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n271), .A2(KEYINPUT4), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n272), .A2(new_n237), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n288), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n282), .A2(new_n278), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n291), .B(new_n292), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n293), .A2(KEYINPUT6), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n235), .B1(new_n299), .B2(new_n289), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n300), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n219), .B(new_n226), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n294), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G210), .B1(G237), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n317));
  INV_X1    g131(.A(new_n235), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n306), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT6), .A3(new_n293), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n311), .C1(new_n300), .C2(new_n307), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n294), .A3(new_n314), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n317), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n314), .B1(new_n321), .B2(new_n294), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT94), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT95), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT95), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n329), .A3(new_n324), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT9), .B(G234), .ZN(new_n332));
  OAI21_X1  g146(.A(G221), .B1(new_n332), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n215), .A2(new_n216), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n273), .A3(new_n288), .ZN(new_n336));
  INV_X1    g150(.A(G134), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT11), .B1(new_n337), .B2(G137), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  INV_X1    g153(.A(G137), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G134), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n337), .A2(G137), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n338), .A2(new_n341), .B1(new_n337), .B2(G137), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n343), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n242), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n207), .A2(new_n208), .B1(G128), .B2(new_n352), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n271), .B(new_n350), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n195), .B1(new_n214), .B2(new_n188), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n200), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n211), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n355), .B(new_n242), .C1(new_n247), .C2(new_n249), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n336), .A2(new_n349), .A3(new_n356), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT86), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n354), .A2(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT86), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n336), .A4(new_n349), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n354), .B1(new_n359), .B2(new_n250), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n349), .A2(KEYINPUT87), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT12), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G140), .ZN(new_n376));
  INV_X1    g190(.A(G953), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(G227), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n376), .B(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n363), .B2(new_n366), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n364), .A2(new_n336), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n347), .B(new_n343), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n375), .A2(new_n379), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G469), .B1(new_n384), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(G469), .ZN(new_n386));
  INV_X1    g200(.A(G902), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n380), .A2(new_n374), .ZN(new_n388));
  INV_X1    g202(.A(new_n379), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n367), .B2(new_n383), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n334), .B1(new_n385), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G217), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n332), .A2(new_n393), .A3(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G116), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n238), .B1(new_n397), .B2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n252), .A2(G122), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  OR2_X1    g215(.A1(KEYINPUT68), .A2(G128), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT68), .A2(G128), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G143), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n187), .A2(G128), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n405), .B1(new_n404), .B2(new_n406), .ZN(new_n408));
  OAI21_X1  g222(.A(G134), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n198), .A2(new_n199), .A3(new_n187), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n209), .A2(G143), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT98), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n337), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n401), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n411), .A2(KEYINPUT13), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n404), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n400), .A2(G107), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G122), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n238), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n419), .A2(G134), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n395), .B1(new_n415), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n401), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n407), .A2(new_n408), .A3(G134), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n337), .B1(new_n412), .B2(new_n413), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n414), .A2(new_n423), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n394), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n387), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n433), .B(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G952), .A3(new_n377), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT16), .ZN(new_n446));
  INV_X1    g260(.A(G140), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G125), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT80), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n202), .B2(KEYINPUT78), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n447), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n450), .B(G140), .C1(new_n202), .C2(KEYINPUT78), .ZN(new_n453));
  NAND3_X1  g267(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(KEYINPUT16), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n204), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n455), .A3(G146), .ZN(new_n458));
  NOR2_X1   g272(.A1(G237), .A2(G953), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(G143), .A3(G214), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(G143), .B1(new_n459), .B2(G214), .ZN(new_n462));
  OAI21_X1  g276(.A(G131), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n463), .A2(KEYINPUT17), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(G214), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n187), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n343), .A3(new_n460), .ZN(new_n467));
  AOI21_X1  g281(.A(KEYINPUT17), .B1(new_n463), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n457), .B(new_n458), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT18), .B(G131), .C1(new_n461), .C2(new_n462), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n466), .A2(new_n460), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n451), .B2(new_n447), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n204), .B1(new_n476), .B2(new_n453), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT96), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n202), .A2(new_n447), .ZN(new_n479));
  NOR2_X1   g293(.A1(G125), .A2(G140), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n205), .A2(new_n206), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT78), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT79), .B1(new_n485), .B2(G125), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n454), .B1(new_n486), .B2(G140), .ZN(new_n487));
  INV_X1    g301(.A(new_n453), .ZN(new_n488));
  OAI21_X1  g302(.A(G146), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n192), .B1(new_n479), .B2(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT96), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n474), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(G113), .B(G122), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n240), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n469), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n469), .B2(new_n492), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n387), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G475), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT20), .ZN(new_n499));
  INV_X1    g313(.A(new_n494), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT19), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(new_n503), .C1(new_n479), .C2(new_n480), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n487), .A2(new_n488), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n192), .B(new_n504), .C1(new_n505), .C2(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n463), .A2(new_n467), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(new_n458), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n478), .B1(new_n477), .B2(new_n483), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n489), .A2(KEYINPUT96), .A3(new_n490), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n473), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n500), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n469), .A2(new_n492), .A3(new_n494), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n499), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n515), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT20), .B(new_n517), .C1(new_n512), .C2(new_n513), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n498), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n438), .A2(new_n445), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n392), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n331), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT99), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n393), .B1(G234), .B2(new_n387), .ZN(new_n525));
  NOR2_X1   g339(.A1(KEYINPUT83), .A2(KEYINPUT25), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT75), .B1(new_n209), .B2(G119), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n528), .B1(new_n200), .B2(G119), .ZN(new_n529));
  NOR4_X1   g343(.A1(new_n198), .A2(new_n199), .A3(KEYINPUT75), .A4(new_n256), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT76), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT24), .B(G110), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT77), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n402), .A2(G119), .A3(new_n403), .ZN(new_n534));
  INV_X1    g348(.A(new_n528), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT75), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n200), .A2(new_n537), .A3(G119), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n531), .A2(new_n533), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n209), .A2(G119), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n402), .A2(KEYINPUT23), .A3(G119), .A4(new_n403), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G110), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n449), .A2(new_n455), .A3(G146), .ZN(new_n549));
  AOI21_X1  g363(.A(G146), .B1(new_n449), .B2(new_n455), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n458), .A2(new_n490), .ZN(new_n553));
  INV_X1    g367(.A(new_n533), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n539), .B1(new_n536), .B2(new_n538), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n544), .A2(new_n545), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT81), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n553), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT82), .B1(new_n552), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n559), .B(KEYINPUT81), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n533), .B1(new_n531), .B2(new_n540), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n458), .B(new_n490), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n541), .B(new_n547), .C1(new_n549), .C2(new_n550), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n377), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n566), .A2(new_n568), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT82), .A3(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n527), .B1(new_n577), .B2(new_n387), .ZN(new_n578));
  AOI211_X1 g392(.A(G902), .B(new_n526), .C1(new_n574), .C2(new_n576), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n525), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n525), .A2(G902), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n574), .A2(KEYINPUT84), .A3(new_n576), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT66), .B1(new_n340), .B2(G134), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT66), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n337), .A3(G137), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n340), .A2(G134), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT67), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(G131), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n345), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n591), .B2(G131), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT70), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n591), .A2(G131), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT67), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT70), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n345), .A4(new_n593), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n600), .A3(new_n359), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n216), .B(new_n215), .C1(new_n346), .C2(new_n348), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n305), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT28), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT28), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n305), .A4(new_n602), .ZN(new_n606));
  INV_X1    g420(.A(new_n305), .ZN(new_n607));
  INV_X1    g421(.A(new_n359), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n598), .A2(new_n345), .A3(new_n593), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n604), .A2(new_n606), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n459), .A2(G210), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT27), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT26), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT72), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n603), .A2(new_n615), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT71), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT30), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n621), .B1(new_n335), .B2(new_n382), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  AND4_X1   g438(.A1(new_n620), .A2(new_n622), .A3(new_n624), .A4(new_n607), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n305), .B1(new_n610), .B2(new_n621), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n620), .B1(new_n626), .B2(new_n624), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n619), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT31), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n594), .A2(new_n595), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n631), .A2(new_n359), .B1(new_n335), .B2(new_n382), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n607), .B1(new_n632), .B2(KEYINPUT30), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n602), .A2(KEYINPUT30), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n609), .A2(KEYINPUT70), .B1(new_n201), .B2(new_n211), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n600), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT71), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n626), .A2(new_n620), .A3(new_n624), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(KEYINPUT31), .A3(new_n619), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n617), .B1(new_n630), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(G472), .A2(G902), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT32), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n617), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT31), .B1(new_n639), .B2(new_n619), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n629), .B(new_n618), .C1(new_n637), .C2(new_n638), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT32), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n603), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n637), .B2(new_n638), .ZN(new_n653));
  OAI21_X1  g467(.A(KEYINPUT73), .B1(new_n653), .B2(new_n615), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n603), .B1(new_n625), .B2(new_n627), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT73), .ZN(new_n656));
  INV_X1    g470(.A(new_n615), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT29), .B1(new_n611), .B2(new_n616), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n604), .A2(new_n606), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n601), .A2(new_n602), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n607), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n615), .A2(KEYINPUT29), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT74), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT74), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n661), .A2(new_n667), .A3(new_n663), .A4(new_n664), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G472), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n586), .B1(new_n651), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n331), .A2(new_n673), .A3(new_n522), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n524), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT100), .B(G101), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G3));
  OAI21_X1  g491(.A(G472), .B1(new_n641), .B2(G902), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n678), .B1(new_n641), .B2(new_n643), .ZN(new_n679));
  INV_X1    g493(.A(new_n392), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n586), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n445), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n321), .A2(new_n294), .A3(new_n314), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n324), .B1(new_n683), .B2(new_n325), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT101), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n415), .B2(new_n424), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT33), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n432), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n425), .A2(new_n687), .A3(new_n431), .A4(KEYINPUT33), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n434), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n432), .A2(new_n434), .A3(new_n387), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n434), .A2(new_n387), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n519), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n519), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n702), .B(new_n324), .C1(new_n683), .C2(new_n325), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n682), .A2(new_n685), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n681), .A2(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT34), .B(G104), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G6));
  NOR2_X1   g521(.A1(new_n519), .A2(new_n437), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n682), .A2(new_n685), .A3(new_n703), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n681), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT104), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT35), .B(G107), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G9));
  NOR2_X1   g527(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n575), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n583), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n580), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n679), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n524), .A2(new_n674), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(KEYINPUT105), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT37), .B(G110), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G12));
  NAND2_X1  g537(.A1(new_n651), .A2(new_n671), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n685), .A2(new_n703), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n717), .A2(new_n392), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT106), .B(G900), .Z(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n443), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n440), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n708), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n724), .A2(new_n726), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G128), .ZN(G30));
  NAND2_X1  g548(.A1(new_n323), .A2(new_n326), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT38), .Z(new_n736));
  INV_X1    g550(.A(new_n628), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n616), .B1(new_n663), .B2(new_n603), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n387), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(G472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n651), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n324), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n514), .A2(new_n515), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT20), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n514), .A2(new_n499), .A3(new_n515), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n744), .A2(new_n745), .B1(G475), .B2(new_n497), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n717), .A2(new_n742), .A3(new_n437), .A4(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n736), .A2(new_n741), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n730), .B(KEYINPUT39), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n392), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT40), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G143), .ZN(G45));
  NAND3_X1  g570(.A1(new_n696), .A2(new_n519), .A3(new_n730), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n696), .A2(new_n519), .A3(KEYINPUT108), .A4(new_n730), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n724), .A2(new_n726), .A3(new_n727), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G146), .ZN(G48));
  NAND2_X1  g577(.A1(new_n367), .A2(new_n383), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n764), .A2(new_n379), .B1(new_n380), .B2(new_n374), .ZN(new_n765));
  OAI21_X1  g579(.A(G469), .B1(new_n765), .B2(G902), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n333), .A3(new_n391), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n769), .A3(new_n391), .A4(new_n333), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n672), .A2(new_n704), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT41), .B(G113), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT110), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n772), .B(new_n774), .ZN(G15));
  NAND3_X1  g589(.A1(new_n672), .A2(new_n709), .A3(new_n771), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G116), .ZN(G18));
  AND2_X1   g591(.A1(new_n717), .A2(new_n520), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n771), .A2(new_n724), .A3(new_n726), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G119), .ZN(G21));
  NOR2_X1   g594(.A1(new_n746), .A2(new_n437), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n682), .A2(new_n685), .A3(new_n703), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n580), .B2(new_n585), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n580), .A2(new_n783), .A3(new_n585), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n642), .B(KEYINPUT111), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n646), .A2(new_n647), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n616), .B1(new_n661), .B2(new_n663), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n678), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n782), .A2(new_n771), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G122), .ZN(G24));
  AND4_X1   g608(.A1(new_n703), .A2(new_n768), .A3(new_n685), .A4(new_n770), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n678), .A2(new_n717), .A3(new_n791), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n759), .A2(new_n760), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G125), .ZN(G27));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n765), .A2(G469), .A3(G902), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n367), .A2(new_n389), .A3(new_n383), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n368), .A2(new_n369), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT12), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n371), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n366), .B2(new_n363), .ZN(new_n807));
  OAI211_X1 g621(.A(G469), .B(new_n803), .C1(new_n807), .C2(new_n389), .ZN(new_n808));
  NAND2_X1  g622(.A1(G469), .A2(G902), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT113), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n801), .B1(new_n802), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n391), .A2(KEYINPUT114), .A3(new_n808), .A4(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n333), .A2(new_n324), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n323), .B2(new_n326), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n797), .A2(KEYINPUT42), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n672), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n761), .A3(new_n816), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n580), .A2(new_n783), .A3(new_n585), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n784), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n644), .A2(new_n650), .B1(new_n670), .B2(G472), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT42), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n343), .ZN(G33));
  NAND3_X1  g641(.A1(new_n817), .A2(new_n672), .A3(new_n732), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G134), .ZN(G36));
  OR2_X1    g643(.A1(new_n384), .A2(KEYINPUT45), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n384), .A2(KEYINPUT45), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(G469), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT46), .B1(new_n832), .B2(new_n810), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n802), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(KEYINPUT46), .A3(new_n810), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n334), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n752), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT44), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n519), .A2(KEYINPUT43), .A3(new_n691), .A4(new_n695), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(new_n696), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n839), .B1(new_n842), .B2(KEYINPUT43), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n679), .A3(new_n717), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n837), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n735), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n742), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n844), .B2(new_n838), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(KEYINPUT116), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n340), .ZN(G39));
  OR2_X1    g666(.A1(new_n836), .A2(KEYINPUT47), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n836), .A2(KEYINPUT47), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n823), .A2(new_n847), .A3(new_n586), .A4(new_n761), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  INV_X1    g672(.A(new_n736), .ZN(new_n859));
  INV_X1    g673(.A(new_n741), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n766), .A2(new_n391), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT49), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n815), .A3(new_n842), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n859), .A2(new_n860), .A3(new_n787), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n817), .A2(new_n672), .A3(new_n732), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n678), .A2(new_n717), .A3(new_n791), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n761), .A3(new_n814), .A4(new_n816), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n746), .A2(new_n437), .A3(new_n730), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n742), .B(new_n869), .C1(new_n323), .C2(new_n326), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n641), .A2(KEYINPUT32), .A3(new_n643), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n649), .B1(new_n648), .B2(new_n642), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(G472), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n660), .B2(new_n669), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n870), .B(new_n727), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT117), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n828), .A2(new_n879), .A3(new_n868), .A4(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n772), .A2(new_n793), .A3(new_n776), .A4(new_n779), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n826), .ZN(new_n883));
  INV_X1    g697(.A(new_n708), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n445), .B1(new_n884), .B2(new_n697), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n681), .A2(new_n331), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n673), .B1(new_n331), .B2(new_n522), .ZN(new_n887));
  AOI211_X1 g701(.A(KEYINPUT99), .B(new_n521), .C1(new_n328), .C2(new_n330), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n886), .B1(new_n889), .B2(new_n672), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n881), .A2(new_n883), .A3(new_n720), .A4(new_n890), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n725), .A2(new_n718), .A3(new_n680), .A4(new_n731), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n892), .A2(new_n724), .B1(new_n795), .B2(new_n798), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n894));
  INV_X1    g708(.A(new_n730), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n717), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n333), .A3(new_n814), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n580), .A2(KEYINPUT118), .A3(new_n716), .A4(new_n730), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n685), .A3(new_n703), .A4(new_n781), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n741), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n893), .A2(new_n901), .A3(KEYINPUT52), .A4(new_n762), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT52), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n799), .A2(new_n733), .A3(new_n762), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n860), .A2(new_n897), .A3(new_n899), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n865), .B1(new_n891), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n822), .A2(new_n823), .ZN(new_n909));
  INV_X1    g723(.A(new_n820), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n825), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n817), .A2(new_n672), .A3(new_n818), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n793), .A2(new_n772), .A3(new_n779), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(new_n776), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n681), .A2(new_n331), .A3(new_n885), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n675), .A2(new_n720), .A3(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n902), .A2(new_n906), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n881), .ZN(new_n920));
  INV_X1    g734(.A(new_n893), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT53), .B1(new_n921), .B2(KEYINPUT52), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n908), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n865), .B1(new_n921), .B2(KEYINPUT52), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n918), .A2(new_n919), .A3(new_n881), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n908), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n771), .A2(new_n847), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n843), .A2(new_n441), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n909), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT48), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n377), .A2(G952), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n787), .A2(new_n792), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n931), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n934), .B1(new_n937), .B2(new_n795), .ZN(new_n938));
  INV_X1    g752(.A(new_n701), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n741), .A2(new_n586), .A3(new_n440), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n930), .A2(new_n940), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n933), .B(new_n938), .C1(new_n939), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n859), .A2(new_n742), .A3(new_n771), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n937), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT50), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(KEYINPUT50), .A3(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(KEYINPUT51), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n930), .A2(new_n931), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(new_n796), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n941), .A2(new_n519), .A3(new_n696), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n853), .B(new_n854), .C1(new_n333), .C2(new_n861), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n936), .A2(new_n742), .A3(new_n846), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n951), .B(new_n952), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n942), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n946), .A2(KEYINPUT120), .A3(new_n947), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n960), .B2(KEYINPUT51), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n929), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(G952), .A2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n864), .B1(new_n962), .B2(new_n963), .ZN(G75));
  NOR2_X1   g778(.A1(new_n377), .A2(G952), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n387), .B1(new_n908), .B2(new_n926), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT56), .B1(new_n967), .B2(G210), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n310), .A2(new_n312), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n321), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n966), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n968), .B2(new_n972), .ZN(G51));
  XOR2_X1   g788(.A(new_n810), .B(KEYINPUT57), .Z(new_n975));
  AND2_X1   g789(.A1(new_n927), .A2(new_n928), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n927), .A2(new_n928), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n765), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n832), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n967), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n965), .B1(new_n980), .B2(new_n982), .ZN(G54));
  AND2_X1   g797(.A1(KEYINPUT58), .A2(G475), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n967), .A2(new_n514), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n514), .B1(new_n967), .B2(new_n984), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n986), .A3(new_n965), .ZN(G60));
  AND2_X1   g801(.A1(new_n689), .A2(new_n690), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n693), .B(KEYINPUT59), .Z(new_n989));
  OAI211_X1 g803(.A(new_n988), .B(new_n989), .C1(new_n976), .C2(new_n977), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n966), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n929), .B2(new_n989), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(new_n992), .ZN(G63));
  NAND2_X1  g807(.A1(G217), .A2(G902), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT60), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n715), .B(KEYINPUT121), .Z(new_n997));
  NAND3_X1  g811(.A1(new_n927), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT122), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g814(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n995), .B1(new_n908), .B2(new_n926), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n582), .A2(new_n584), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n966), .B(new_n1001), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(KEYINPUT122), .A3(new_n997), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1000), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n927), .A2(new_n996), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1003), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n966), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT123), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1009), .A2(new_n966), .A3(new_n998), .A4(new_n1001), .ZN(new_n1013));
  AOI22_X1  g827(.A1(new_n1007), .A2(new_n1012), .B1(KEYINPUT61), .B2(new_n1013), .ZN(G66));
  NOR2_X1   g828(.A1(new_n917), .A2(new_n882), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(G953), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT124), .ZN(new_n1017));
  OAI21_X1  g831(.A(G953), .B1(new_n220), .B2(new_n444), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n310), .B1(G898), .B2(new_n377), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1020), .B(KEYINPUT125), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1019), .B(new_n1021), .ZN(G69));
  NAND2_X1  g836(.A1(new_n622), .A2(new_n624), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n504), .B1(new_n505), .B2(new_n501), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1024), .B(KEYINPUT126), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1023), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n857), .B1(new_n849), .B2(new_n850), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n909), .A2(new_n726), .A3(new_n781), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n913), .B(new_n828), .C1(new_n837), .C2(new_n1028), .ZN(new_n1029));
  NOR4_X1   g843(.A1(new_n1027), .A2(new_n1029), .A3(G953), .A4(new_n904), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G900), .A2(G953), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1026), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G227), .A2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(G953), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n755), .A2(new_n762), .A3(new_n893), .ZN(new_n1036));
  OR2_X1    g850(.A1(new_n1036), .A2(KEYINPUT62), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1027), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n884), .A2(new_n697), .ZN(new_n1039));
  AND4_X1   g853(.A1(new_n672), .A2(new_n753), .A3(new_n847), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1040), .B1(new_n1036), .B2(KEYINPUT62), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1026), .A2(G953), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1033), .A2(new_n1035), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1035), .B1(new_n1033), .B2(new_n1044), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1045), .A2(new_n1046), .ZN(G72));
  NAND4_X1  g861(.A1(new_n1037), .A2(new_n1038), .A3(new_n1041), .A4(new_n1015), .ZN(new_n1048));
  XNOR2_X1  g862(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1049));
  NOR2_X1   g863(.A1(new_n874), .A2(new_n387), .ZN(new_n1050));
  XOR2_X1   g864(.A(new_n1049), .B(new_n1050), .Z(new_n1051));
  AOI211_X1 g865(.A(new_n657), .B(new_n653), .C1(new_n1048), .C2(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1051), .ZN(new_n1053));
  NOR3_X1   g867(.A1(new_n1027), .A2(new_n904), .A3(new_n1029), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n1015), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n653), .A2(new_n657), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n966), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n654), .A2(new_n658), .A3(new_n628), .ZN(new_n1058));
  AND3_X1   g872(.A1(new_n923), .A2(new_n1051), .A3(new_n1058), .ZN(new_n1059));
  NOR3_X1   g873(.A1(new_n1052), .A2(new_n1057), .A3(new_n1059), .ZN(G57));
endmodule


