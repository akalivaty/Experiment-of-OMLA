//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT64), .A2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G143), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT92), .A4(new_n191), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n187), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n191), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT92), .B1(new_n197), .B2(new_n189), .ZN(new_n198));
  OAI211_X1 g012(.A(KEYINPUT18), .B(G131), .C1(new_n194), .C2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n199), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n197), .A2(new_n189), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT92), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n193), .A4(new_n192), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n216), .A3(new_n193), .A4(new_n192), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT93), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n194), .A2(new_n198), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n220), .C1(new_n216), .C2(new_n214), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n210), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT94), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT94), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n210), .A2(new_n218), .A3(new_n224), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(KEYINPUT17), .B(G131), .C1(new_n194), .C2(new_n198), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n204), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  OAI211_X1 g046(.A(G146), .B(new_n229), .C1(new_n204), .C2(new_n230), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n194), .B2(new_n198), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n215), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n227), .B(new_n234), .C1(KEYINPUT17), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G113), .B(G122), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT95), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n238), .B2(new_n243), .ZN(new_n246));
  OR2_X1    g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n238), .A2(new_n241), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n206), .B(KEYINPUT19), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n207), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n236), .A2(new_n233), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n242), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n223), .B2(new_n225), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT20), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n242), .B1(new_n226), .B2(new_n237), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n255), .ZN(new_n261));
  AOI22_X1  g075(.A1(G475), .A2(new_n247), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G143), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT97), .B1(new_n263), .B2(G128), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT97), .ZN(new_n265));
  INV_X1    g079(.A(G128), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n190), .A2(G128), .A3(new_n191), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT66), .B(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n272), .A2(G122), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(G122), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G107), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n268), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n269), .A2(new_n278), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT96), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n269), .A2(KEYINPUT96), .A3(new_n278), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G134), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n271), .B(new_n277), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n268), .A2(new_n269), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n271), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT14), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n275), .B(G107), .C1(new_n294), .C2(new_n274), .ZN(new_n295));
  OAI21_X1  g109(.A(G107), .B1(new_n274), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n274), .B2(new_n273), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n293), .A2(new_n298), .A3(KEYINPUT98), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT98), .B1(new_n293), .B2(new_n298), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n286), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  INV_X1    g117(.A(G217), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(new_n304), .A3(G953), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n286), .B(new_n305), .C1(new_n300), .C2(new_n301), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G478), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT15), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n309), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n262), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G140), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n188), .A2(G227), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G101), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n276), .A2(G104), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n240), .A2(G107), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n321), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n240), .A2(G107), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT85), .B(KEYINPUT3), .C1(new_n240), .C2(G107), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n322), .B1(new_n329), .B2(new_n319), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n190), .A2(G146), .A3(new_n191), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n263), .A2(G146), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n331), .A2(G128), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n207), .B1(new_n195), .B2(new_n196), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n266), .B1(new_n336), .B2(KEYINPUT1), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n333), .B1(new_n197), .B2(G146), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND4_X1   g158(.A1(KEYINPUT0), .A2(new_n331), .A3(G128), .A4(new_n334), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n336), .B1(G143), .B2(new_n207), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT0), .B(G128), .Z(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(KEYINPUT65), .A3(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n207), .A2(G143), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n190), .A2(new_n191), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n350), .B1(new_n351), .B2(new_n207), .ZN(new_n352));
  INV_X1    g166(.A(new_n347), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n349), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n345), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n276), .A2(G104), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n326), .B2(new_n325), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT85), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(new_n328), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G101), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n357), .B(new_n319), .C1(new_n358), .C2(new_n359), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n364), .A3(G101), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n355), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G128), .B1(new_n332), .B2(new_n333), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n335), .B1(new_n368), .B2(new_n352), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n330), .A3(KEYINPUT10), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n340), .A2(KEYINPUT86), .A3(new_n341), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n344), .A2(new_n366), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n288), .A2(new_n290), .A3(G137), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT67), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT11), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n375), .A2(new_n285), .A3(G137), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT67), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n288), .A2(new_n290), .A3(new_n379), .A4(G137), .ZN(new_n380));
  AOI21_X1  g194(.A(G137), .B1(new_n288), .B2(new_n290), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n381), .B2(KEYINPUT11), .ZN(new_n382));
  OAI21_X1  g196(.A(G131), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n376), .B1(new_n373), .B2(KEYINPUT67), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n375), .B1(new_n270), .B2(G137), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n384), .A2(new_n214), .A3(new_n380), .A4(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT72), .B1(new_n383), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n318), .B1(new_n372), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n392));
  INV_X1    g206(.A(G137), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT11), .B1(new_n291), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n380), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n214), .B1(new_n396), .B2(new_n384), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n214), .A2(new_n384), .A3(new_n380), .A4(new_n385), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n392), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n386), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n332), .A2(G128), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n346), .A2(new_n367), .B1(new_n338), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n322), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n362), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n399), .A2(new_n400), .B1(new_n340), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT87), .B1(new_n406), .B2(KEYINPUT12), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n340), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n408), .B(new_n409), .C1(new_n389), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n410), .B(KEYINPUT12), .C1(new_n398), .C2(new_n397), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n391), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n372), .A2(new_n390), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n366), .A2(new_n370), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n417), .A2(new_n389), .A3(new_n344), .A4(new_n371), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n318), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n314), .B(new_n245), .C1(new_n415), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n391), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n416), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n372), .A2(new_n390), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n423), .B1(new_n413), .B2(new_n414), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(G469), .C1(new_n424), .C2(new_n318), .ZN(new_n425));
  NAND2_X1  g239(.A1(G469), .A2(G902), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT2), .A2(G113), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT2), .A2(G113), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(KEYINPUT71), .A2(KEYINPUT2), .A3(G113), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G119), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G113), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n272), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G119), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n272), .A2(G119), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT5), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n330), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n363), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n437), .A2(new_n438), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n439), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n365), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n450), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT6), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(KEYINPUT6), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n327), .A2(new_n328), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n319), .B1(new_n461), .B2(new_n357), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n462), .A2(new_n364), .B1(new_n452), .B2(new_n439), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n463), .A2(new_n363), .B1(new_n330), .B2(new_n449), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n460), .B1(new_n464), .B2(new_n457), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n457), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n402), .A2(new_n202), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n355), .B2(new_n202), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n188), .A2(G224), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n469), .B(new_n470), .Z(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n457), .B(KEYINPUT8), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n362), .A2(new_n403), .B1(new_n439), .B2(new_n448), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n447), .A2(KEYINPUT89), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n443), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n447), .A2(KEYINPUT89), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n439), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI22_X1  g292(.A1(new_n474), .A2(KEYINPUT90), .B1(new_n478), .B2(new_n404), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n330), .A2(new_n449), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n473), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n470), .A2(KEYINPUT7), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n469), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n483), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n468), .B(new_n485), .C1(new_n355), .C2(new_n202), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n464), .A2(new_n457), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n482), .A2(new_n484), .A3(KEYINPUT91), .A4(new_n486), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n472), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G210), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n472), .A2(new_n492), .A3(new_n494), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n431), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G952), .ZN(new_n499));
  AOI211_X1 g313(.A(G953), .B(new_n499), .C1(G234), .C2(G237), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n245), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT21), .B(G898), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n313), .A2(new_n429), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n355), .B1(new_n387), .B2(new_n388), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n393), .A2(G134), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n508), .B(G131), .C1(new_n381), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n509), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n270), .B2(G137), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n508), .B1(new_n513), .B2(G131), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n386), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G131), .B1(new_n381), .B2(new_n509), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT68), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT73), .A3(new_n386), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n521), .A3(new_n369), .ZN(new_n522));
  INV_X1    g336(.A(new_n453), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n507), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT74), .B(KEYINPUT27), .Z(new_n525));
  NAND3_X1  g339(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT26), .B(G101), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n527), .B(new_n528), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n507), .B2(new_n522), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT70), .B1(new_n515), .B2(new_n402), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n355), .B1(new_n397), .B2(new_n398), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT70), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n520), .A2(new_n537), .A3(new_n369), .A4(new_n386), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n533), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n453), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n524), .A2(KEYINPUT75), .A3(new_n529), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT31), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n524), .A2(KEYINPUT28), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n507), .A2(new_n522), .A3(new_n545), .A4(new_n523), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n453), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n529), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT31), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n532), .A2(new_n540), .A3(new_n553), .A4(new_n541), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n543), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(G472), .A2(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n523), .B1(new_n507), .B2(new_n522), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n547), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n551), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n540), .A2(new_n524), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n551), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT76), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n547), .A2(new_n569), .A3(new_n529), .A4(new_n549), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n547), .A2(new_n529), .A3(new_n549), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n572), .A2(KEYINPUT76), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n566), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  INV_X1    g389(.A(new_n556), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n558), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n555), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT77), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n555), .A2(KEYINPUT77), .A3(new_n577), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n559), .A2(new_n575), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n304), .B1(G234), .B2(new_n245), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n266), .A2(G119), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT79), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n444), .A2(G128), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT23), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n266), .A2(KEYINPUT79), .A3(G119), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G110), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT78), .ZN(new_n592));
  NAND2_X1  g406(.A1(KEYINPUT23), .A2(G119), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n592), .B1(new_n593), .B2(G128), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n266), .A2(KEYINPUT78), .A3(KEYINPUT23), .A4(G119), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(KEYINPUT81), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT81), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n590), .A2(new_n599), .A3(new_n591), .A4(new_n596), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n587), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT24), .B(G110), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n233), .B(new_n208), .C1(new_n598), .C2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT82), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n601), .A2(new_n602), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n590), .A2(new_n596), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(G110), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n232), .A2(new_n233), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT80), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n611), .B1(new_n609), .B2(new_n610), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n605), .B(new_n606), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT22), .B(G137), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n615), .B(new_n616), .Z(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n605), .B1(new_n612), .B2(new_n613), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n614), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n622), .B2(new_n617), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT25), .B1(new_n623), .B2(new_n245), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n618), .B1(new_n621), .B2(new_n614), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  NOR4_X1   g440(.A1(new_n625), .A2(new_n619), .A3(new_n626), .A4(G902), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n583), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n623), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n583), .A2(G902), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT83), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT84), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT84), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n628), .A2(new_n636), .A3(new_n633), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n506), .A2(new_n582), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(G101), .ZN(G3));
  OAI21_X1  g454(.A(G475), .B1(new_n244), .B2(new_n246), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n260), .B1(new_n259), .B2(new_n255), .ZN(new_n642));
  INV_X1    g456(.A(new_n255), .ZN(new_n643));
  NOR4_X1   g457(.A1(new_n258), .A2(KEYINPUT20), .A3(new_n253), .A4(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n310), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n307), .A2(new_n308), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(KEYINPUT33), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n307), .B2(new_n308), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n245), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(G478), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT100), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n309), .A2(new_n656), .A3(new_n653), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n651), .B(KEYINPUT101), .C1(new_n655), .C2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n652), .A2(KEYINPUT100), .A3(new_n654), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n656), .B1(new_n309), .B2(new_n653), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(KEYINPUT101), .B1(new_n662), .B2(new_n651), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n645), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT102), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n645), .B(new_n666), .C1(new_n659), .C2(new_n663), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n505), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n429), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n555), .A2(new_n245), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n670), .A2(G472), .B1(new_n556), .B2(new_n555), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n668), .A2(new_n638), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  NOR2_X1   g488(.A1(new_n645), .A2(new_n312), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n505), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n638), .A3(new_n669), .A4(new_n671), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  XNOR2_X1  g494(.A(new_n620), .B(KEYINPUT103), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n618), .A2(KEYINPUT36), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n631), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n628), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n529), .B1(new_n547), .B2(new_n549), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n532), .A2(new_n540), .A3(new_n541), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n687), .B1(new_n688), .B2(new_n553), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n543), .ZN(new_n690));
  INV_X1    g504(.A(G472), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n557), .B(new_n686), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT104), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n671), .A2(new_n694), .A3(new_n686), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n695), .A3(new_n506), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT105), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n696), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(new_n500), .ZN(new_n700));
  INV_X1    g514(.A(new_n501), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(G900), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n675), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n686), .A2(new_n427), .A3(new_n498), .A4(new_n428), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n582), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n702), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n669), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n496), .A2(new_n497), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT38), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR4_X1   g528(.A1(new_n714), .A2(new_n312), .A3(new_n262), .A4(new_n431), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n710), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n580), .A2(new_n581), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n529), .B1(new_n561), .B2(new_n524), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n245), .B1(new_n688), .B2(new_n718), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n557), .A2(new_n558), .B1(G472), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n686), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n197), .ZN(G45));
  OAI211_X1 g539(.A(new_n645), .B(new_n702), .C1(new_n659), .C2(new_n663), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n704), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n582), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT106), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n582), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND2_X1  g547(.A1(new_n635), .A2(new_n637), .ZN(new_n734));
  AOI22_X1  g548(.A1(G472), .A2(new_n574), .B1(new_n557), .B2(new_n558), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n717), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n415), .A2(new_n419), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n428), .A3(new_n420), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n736), .A2(new_n668), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT107), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n741), .B(new_n743), .ZN(G15));
  NAND4_X1  g558(.A1(new_n582), .A2(new_n677), .A3(new_n638), .A4(new_n740), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT108), .B(G116), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G18));
  AND2_X1   g561(.A1(new_n740), .A2(new_n498), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n313), .A2(new_n503), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n582), .A3(new_n686), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  INV_X1    g565(.A(new_n554), .ZN(new_n752));
  AOI22_X1  g566(.A1(new_n542), .A2(KEYINPUT31), .B1(new_n562), .B2(new_n551), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n753), .B2(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n562), .A2(new_n551), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n543), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT109), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n576), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n690), .B2(new_n691), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n670), .A2(KEYINPUT110), .A3(G472), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n634), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n262), .A2(new_n312), .A3(new_n503), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n763), .A2(new_n764), .A3(new_n748), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  INV_X1    g581(.A(new_n726), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n763), .A2(new_n686), .A3(new_n768), .A4(new_n748), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  AND3_X1   g584(.A1(new_n472), .A2(new_n492), .A3(new_n494), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n494), .B1(new_n472), .B2(new_n492), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n771), .A2(new_n772), .A3(new_n431), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n427), .A3(new_n428), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(KEYINPUT111), .ZN(new_n778));
  AND4_X1   g592(.A1(KEYINPUT42), .A2(new_n777), .A3(new_n768), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n575), .A2(new_n559), .A3(new_n578), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n764), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT112), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n780), .B2(new_n764), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n779), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n774), .B(new_n776), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n736), .A2(new_n786), .A3(new_n768), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND4_X1  g605(.A1(new_n736), .A2(new_n675), .A3(new_n702), .A4(new_n786), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  INV_X1    g607(.A(new_n420), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n413), .A2(new_n414), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n418), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n796), .A2(new_n317), .B1(new_n416), .B2(new_n421), .ZN(new_n797));
  OAI21_X1  g611(.A(G469), .B1(new_n797), .B2(KEYINPUT45), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(KEYINPUT45), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT113), .B(G469), .C1(new_n797), .C2(KEYINPUT45), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n426), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n794), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(KEYINPUT46), .A3(new_n426), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n428), .A3(new_n708), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n428), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n806), .B2(new_n807), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(KEYINPUT114), .A3(new_n708), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n262), .B1(new_n663), .B2(new_n659), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT43), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT43), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n671), .A2(new_n722), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n815), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n823), .A3(KEYINPUT44), .A4(new_n821), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n773), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  INV_X1    g643(.A(new_n773), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n582), .A2(new_n638), .A3(new_n726), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n813), .A2(KEYINPUT47), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT47), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n833), .B(new_n812), .C1(new_n806), .C2(new_n807), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G140), .ZN(G42));
  NAND2_X1  g650(.A1(new_n808), .A2(new_n428), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n813), .A2(KEYINPUT47), .ZN(new_n839));
  INV_X1    g653(.A(new_n738), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n794), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n812), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n763), .A2(new_n764), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n822), .A2(new_n844), .A3(new_n700), .A4(new_n830), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n721), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n739), .A2(new_n830), .A3(new_n700), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n638), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  OR3_X1    g664(.A1(new_n645), .A2(new_n659), .A3(new_n663), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n820), .A2(new_n821), .A3(new_n848), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n763), .A2(new_n686), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT121), .ZN(new_n855));
  OAI21_X1  g669(.A(KEYINPUT121), .B1(new_n853), .B2(new_n854), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n820), .A2(new_n500), .A3(new_n821), .ZN(new_n859));
  INV_X1    g673(.A(new_n844), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n714), .A2(new_n431), .A3(new_n740), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT50), .A4(new_n861), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n858), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n846), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n859), .A2(new_n860), .A3(new_n748), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n665), .A2(new_n667), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n847), .A2(new_n849), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(G952), .A3(new_n188), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n781), .B(KEYINPUT112), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n820), .A3(new_n821), .A4(new_n848), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n873), .A2(KEYINPUT48), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(KEYINPUT48), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n857), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n843), .B2(new_n845), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n864), .A2(KEYINPUT120), .A3(new_n865), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT120), .B1(new_n864), .B2(new_n865), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n867), .B(new_n876), .C1(new_n882), .C2(KEYINPUT51), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n505), .A2(new_n664), .A3(new_n429), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n638), .A3(new_n671), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n639), .A2(new_n885), .A3(KEYINPUT116), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT116), .B1(new_n639), .B2(new_n885), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n696), .A2(new_n678), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n786), .A2(new_n763), .A3(new_n686), .A4(new_n768), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n262), .A2(new_n312), .A3(new_n702), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n582), .A2(new_n686), .A3(new_n775), .A4(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n792), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n741), .A2(new_n766), .A3(new_n745), .A4(new_n750), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n889), .A2(new_n790), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n582), .A2(new_n727), .A3(new_n730), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n730), .B1(new_n582), .B2(new_n727), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n769), .B(new_n706), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n312), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n498), .A2(new_n900), .A3(new_n645), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n702), .B(KEYINPUT117), .Z(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n429), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n721), .A2(new_n903), .A3(new_n722), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT52), .B1(new_n899), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n705), .A2(new_n582), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n729), .B2(new_n731), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n769), .A4(new_n904), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n896), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n910), .ZN(new_n913));
  XOR2_X1   g727(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n914));
  NOR3_X1   g728(.A1(new_n895), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT54), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n639), .A2(new_n885), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT116), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n888), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n639), .A2(new_n885), .A3(KEYINPUT116), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT53), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n792), .A2(new_n890), .A3(new_n892), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n872), .A2(new_n779), .B1(new_n787), .B2(new_n788), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n741), .A2(new_n745), .A3(new_n750), .A4(new_n766), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT119), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT119), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n790), .A2(new_n894), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n911), .A2(new_n925), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT54), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n914), .B1(new_n895), .B2(new_n913), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n883), .A2(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n764), .A2(new_n714), .A3(new_n430), .A4(new_n428), .ZN(new_n937));
  INV_X1    g751(.A(new_n841), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT49), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n816), .B1(new_n938), .B2(KEYINPUT49), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n847), .A2(new_n937), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n936), .A2(new_n941), .ZN(G75));
  NAND2_X1  g756(.A1(new_n931), .A2(new_n933), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(G210), .A3(G902), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT56), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n467), .B(new_n471), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT55), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n944), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n188), .A2(G952), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(G51));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  INV_X1    g766(.A(new_n803), .ZN(new_n953));
  AND4_X1   g767(.A1(new_n952), .A2(new_n943), .A3(G902), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n245), .B1(new_n931), .B2(new_n933), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n955), .B2(new_n953), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n426), .B(KEYINPUT57), .Z(new_n958));
  AND3_X1   g772(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n737), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n950), .B1(new_n957), .B2(new_n963), .ZN(G54));
  NAND3_X1  g778(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n258), .B2(new_n253), .ZN(new_n966));
  INV_X1    g780(.A(new_n950), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n955), .A2(KEYINPUT58), .A3(G475), .A4(new_n259), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(G60));
  NOR2_X1   g783(.A1(new_n648), .A2(new_n650), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT59), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n973), .C1(new_n959), .C2(new_n960), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n967), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n971), .B1(new_n935), .B2(new_n973), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G63));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n931), .B2(new_n933), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n683), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n967), .B1(new_n981), .B2(new_n623), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n978), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n981), .A2(new_n623), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G66));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n989));
  INV_X1    g803(.A(new_n502), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(G224), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n991), .B2(G953), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n922), .A2(new_n927), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n993), .A2(G953), .ZN(new_n994));
  MUX2_X1   g808(.A(new_n992), .B(new_n989), .S(new_n994), .Z(new_n995));
  INV_X1    g809(.A(new_n467), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(G898), .B2(new_n188), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n995), .B(new_n998), .ZN(G69));
  AND2_X1   g813(.A1(new_n828), .A2(new_n835), .ZN(new_n1000));
  INV_X1    g814(.A(new_n899), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n1001), .B(KEYINPUT62), .C1(new_n723), .C2(new_n716), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT62), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1003), .B1(new_n724), .B2(new_n899), .ZN(new_n1004));
  AOI211_X1 g818(.A(new_n830), .B(new_n709), .C1(new_n664), .C2(new_n676), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1002), .A2(new_n1004), .B1(new_n736), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(G953), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n534), .A2(new_n539), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n249), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(KEYINPUT125), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1009), .B1(G900), .B2(G953), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n872), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1015), .A2(new_n901), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n811), .A2(new_n1016), .A3(new_n814), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n790), .A2(new_n1001), .A3(new_n792), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n828), .A2(new_n1017), .A3(new_n835), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1014), .B1(new_n1019), .B2(new_n188), .ZN(new_n1020));
  OR3_X1    g834(.A1(new_n1011), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1012), .B1(new_n1011), .B2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(G72));
  NAND3_X1  g837(.A1(new_n1000), .A2(new_n993), .A3(new_n1006), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n551), .B1(new_n540), .B2(new_n524), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1025), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1027), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n568), .B2(new_n542), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n912), .B2(new_n915), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1019), .B2(new_n993), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n567), .A2(new_n529), .ZN(new_n1037));
  XNOR2_X1  g851(.A(new_n1037), .B(KEYINPUT127), .ZN(new_n1038));
  OAI211_X1 g852(.A(new_n967), .B(new_n1035), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1032), .A2(new_n1039), .ZN(G57));
endmodule


