//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n466), .A2(G137), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n461), .A2(new_n470), .A3(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n466), .A2(G2105), .A3(new_n469), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(G136), .B2(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n466), .A2(G138), .A3(new_n467), .A4(new_n469), .ZN(new_n486));
  INV_X1    g061(.A(new_n473), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n488), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n489));
  AOI22_X1  g064(.A1(new_n486), .A2(KEYINPUT4), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n490), .A2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT6), .A3(G651), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n496), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G50), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n496), .B1(new_n504), .B2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n509), .B2(new_n498), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n499), .A2(new_n501), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n512), .B1(new_n508), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n510), .B1(G88), .B2(new_n515), .ZN(G166));
  NAND2_X1  g091(.A1(new_n515), .A2(G89), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n500), .A2(KEYINPUT6), .A3(G651), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT6), .B1(new_n500), .B2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n502), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  AND3_X1   g102(.A1(new_n505), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT73), .B1(new_n505), .B2(new_n507), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n517), .A2(new_n525), .A3(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  NAND2_X1  g109(.A1(new_n515), .A2(G90), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n524), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n530), .A2(G64), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n498), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n528), .A2(new_n529), .A3(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(G68), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n524), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n508), .A2(new_n511), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT72), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n508), .A2(new_n511), .A3(new_n512), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G81), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT75), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n548), .A2(G91), .A3(new_n549), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT76), .B(G65), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n508), .A2(new_n560), .B1(G78), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n498), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT9), .B1(new_n520), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n502), .A2(new_n565), .A3(G53), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n559), .A2(new_n562), .A3(new_n567), .ZN(G299));
  AND2_X1   g143(.A1(new_n538), .A2(new_n539), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n536), .B(new_n535), .C1(new_n569), .C2(new_n498), .ZN(G301));
  NAND2_X1  g145(.A1(G75), .A2(G543), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n505), .A2(new_n507), .ZN(new_n572));
  INV_X1    g147(.A(G62), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n548), .A2(new_n549), .ZN(new_n576));
  INV_X1    g151(.A(G88), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n503), .C1(new_n576), .C2(new_n577), .ZN(G303));
  NAND2_X1  g153(.A1(new_n515), .A2(G87), .ZN(new_n579));
  INV_X1    g154(.A(G74), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n528), .B2(new_n529), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G49), .B2(new_n502), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT77), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n572), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(G48), .B2(new_n502), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n515), .A2(KEYINPUT78), .A3(G86), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT78), .B1(new_n515), .B2(G86), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n530), .A2(G60), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n498), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n548), .A2(G85), .A3(new_n549), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n502), .A2(new_n522), .ZN(new_n597));
  AOI211_X1 g172(.A(KEYINPUT74), .B(new_n496), .C1(new_n499), .C2(new_n501), .ZN(new_n598));
  OAI21_X1  g173(.A(G47), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n596), .A2(new_n599), .A3(KEYINPUT79), .ZN(new_n600));
  AOI21_X1  g175(.A(KEYINPUT79), .B1(new_n596), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n576), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n572), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n524), .A2(G54), .B1(new_n611), .B2(G651), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n603), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n603), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND3_X1  g197(.A1(new_n608), .A2(new_n621), .A3(new_n612), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(G111), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n627), .A2(KEYINPUT81), .B1(new_n628), .B2(G2105), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(KEYINPUT81), .B2(new_n627), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n480), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n632), .B1(G135), .B2(new_n484), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n487), .A2(new_n459), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT13), .B(G2100), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2084), .B(G2090), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT83), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n661), .A2(new_n662), .ZN(new_n665));
  AOI21_X1  g240(.A(KEYINPUT18), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  NOR2_X1   g242(.A1(G2072), .A2(G2078), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n663), .B2(KEYINPUT18), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2096), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT19), .Z(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT84), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(new_n674), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n675), .A2(new_n676), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n686), .A3(new_n678), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n683), .A2(new_n684), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT86), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n690), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT87), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  INV_X1    g276(.A(new_n588), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n515), .A2(G86), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT78), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n515), .A2(KEYINPUT78), .A3(G86), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n701), .B1(new_n707), .B2(new_n700), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT32), .B(G1981), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G23), .B(new_n583), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT89), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n716));
  NAND2_X1  g291(.A1(G303), .A2(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G22), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1971), .ZN(new_n723));
  INV_X1    g298(.A(G1971), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n720), .A2(new_n724), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n715), .A2(new_n716), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n716), .B1(new_n715), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n699), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n715), .A2(new_n726), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(KEYINPUT91), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n715), .A2(new_n716), .A3(new_n726), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G24), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n596), .A2(new_n599), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT79), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n596), .A2(new_n599), .A3(KEYINPUT79), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n594), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(G16), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(G1986), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n484), .A2(G131), .ZN(new_n742));
  INV_X1    g317(.A(G119), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n480), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(G107), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT88), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n742), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G25), .B(new_n749), .S(G29), .Z(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n741), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G1986), .B2(new_n740), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n729), .A2(new_n733), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n757), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n729), .A2(new_n733), .A3(new_n759), .A4(new_n755), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n614), .A2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G4), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT93), .B(G1348), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G29), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G33), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n484), .A2(G139), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT25), .ZN(new_n769));
  NAND2_X1  g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(G127), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n473), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n769), .B1(G2105), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n767), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(new_n765), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n775), .A2(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(G2072), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(KEYINPUT24), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(KEYINPUT24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n765), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G160), .B2(new_n765), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G2084), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n776), .A2(new_n777), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n700), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n765), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n634), .B2(new_n765), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G2084), .B2(new_n782), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n784), .A2(new_n788), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n765), .A2(G27), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G164), .B2(new_n765), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n764), .B(new_n795), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n796), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n765), .A2(G35), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n765), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT29), .Z(new_n804));
  INV_X1    g379(.A(G2090), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI211_X1 g381(.A(new_n801), .B(new_n806), .C1(new_n763), .C2(new_n762), .ZN(new_n807));
  NOR2_X1   g382(.A1(G5), .A2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT94), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G301), .B2(new_n700), .ZN(new_n810));
  INV_X1    g385(.A(G1961), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n700), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n700), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n810), .A2(new_n811), .B1(new_n813), .B2(G1966), .ZN(new_n814));
  INV_X1    g389(.A(G1341), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n552), .A2(G16), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G16), .B2(G19), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n814), .B1(new_n815), .B2(new_n817), .C1(G1966), .C2(new_n813), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n765), .A2(G26), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT28), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n484), .A2(G140), .ZN(new_n821));
  INV_X1    g396(.A(G128), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n467), .A2(G116), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n480), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n820), .B1(new_n826), .B2(new_n765), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2067), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n817), .A2(new_n815), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n811), .B2(new_n810), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n818), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n800), .A2(new_n807), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n765), .A2(G32), .ZN(new_n833));
  NAND3_X1  g408(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT26), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n836), .A2(new_n837), .B1(G105), .B2(new_n459), .ZN(new_n838));
  INV_X1    g413(.A(G129), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n480), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G141), .B2(new_n484), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n833), .B1(new_n841), .B2(new_n765), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT27), .ZN(new_n843));
  INV_X1    g418(.A(G1996), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n804), .A2(new_n805), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT96), .Z(new_n847));
  NOR3_X1   g422(.A1(new_n832), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n758), .A2(new_n760), .A3(new_n848), .ZN(G311));
  NAND3_X1  g424(.A1(new_n758), .A2(new_n848), .A3(new_n760), .ZN(G150));
  INV_X1    g425(.A(G67), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n528), .A2(new_n529), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(G80), .A2(G543), .ZN(new_n853));
  OAI21_X1  g428(.A(G651), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n524), .A2(G55), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n548), .A2(G93), .A3(new_n549), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n621), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n515), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n515), .A2(G93), .B1(new_n524), .B2(G55), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n545), .A4(new_n854), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n551), .A2(new_n857), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n859), .B1(new_n870), .B2(new_n872), .ZN(G145));
  INV_X1    g448(.A(G130), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n467), .A2(KEYINPUT98), .A3(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT98), .B1(new_n467), .B2(G118), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(G2104), .A3(new_n877), .ZN(new_n878));
  OAI22_X1  g453(.A1(new_n480), .A2(new_n874), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G142), .B2(new_n484), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(new_n749), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n749), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n639), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n639), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n841), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n826), .A2(G164), .ZN(new_n889));
  OAI22_X1  g464(.A1(new_n821), .A2(new_n825), .B1(new_n490), .B2(new_n494), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n888), .A3(new_n890), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n774), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n774), .ZN(new_n895));
  INV_X1    g470(.A(new_n893), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n887), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(G162), .B(new_n633), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G160), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT100), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n897), .A2(new_n894), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n902), .B1(new_n897), .B2(new_n894), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n887), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(KEYINPUT101), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n901), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n887), .A2(new_n897), .A3(new_n894), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n909), .B2(new_n898), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT99), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT99), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n912), .B(new_n900), .C1(new_n909), .C2(new_n898), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n908), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n908), .B2(new_n914), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(G395));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n583), .A2(G166), .ZN(new_n920));
  NAND3_X1  g495(.A1(G303), .A2(new_n579), .A3(new_n582), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n739), .A2(G305), .ZN(new_n924));
  NOR2_X1   g499(.A1(G290), .A2(new_n707), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n739), .A2(G305), .ZN(new_n927));
  NAND2_X1  g502(.A1(G290), .A2(new_n707), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n922), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G299), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n608), .A2(new_n931), .A3(new_n612), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n608), .B2(new_n612), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n623), .A2(new_n866), .A3(new_n865), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n623), .B1(new_n866), .B2(new_n865), .ZN(new_n936));
  OR3_X1    g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n932), .B2(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n613), .A2(G299), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n608), .A2(new_n931), .A3(new_n612), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n940), .B(new_n944), .C1(new_n935), .C2(new_n936), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n937), .A2(new_n938), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n937), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n930), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n937), .A2(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g525(.A(new_n930), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n937), .A2(new_n938), .A3(new_n945), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G868), .ZN(new_n955));
  INV_X1    g530(.A(new_n857), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G868), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n919), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n617), .B1(new_n948), .B2(new_n953), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n960), .A2(KEYINPUT104), .A3(new_n957), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(G295));
  OR3_X1    g537(.A1(new_n960), .A2(KEYINPUT105), .A3(new_n957), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT105), .B1(new_n960), .B2(new_n957), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n927), .A2(new_n928), .A3(new_n922), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n922), .B1(new_n927), .B2(new_n928), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n926), .A2(KEYINPUT106), .A3(new_n929), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n551), .A2(new_n857), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n551), .A2(new_n857), .ZN(new_n974));
  OAI21_X1  g549(.A(G171), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n865), .A2(new_n866), .A3(G301), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(G168), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n865), .A2(new_n866), .A3(G301), .ZN(new_n978));
  AOI21_X1  g553(.A(G301), .B1(new_n865), .B2(new_n866), .ZN(new_n979));
  OAI21_X1  g554(.A(G286), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n934), .A2(new_n939), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n941), .A2(new_n943), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n942), .ZN(new_n983));
  AND4_X1   g558(.A1(new_n977), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n980), .B2(new_n977), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n972), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G37), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n978), .A2(new_n979), .A3(G286), .ZN(new_n988));
  AOI21_X1  g563(.A(G168), .B1(new_n975), .B2(new_n976), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n934), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n940), .A2(new_n944), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n980), .A3(new_n977), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n930), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n987), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n966), .B1(new_n994), .B2(KEYINPUT43), .ZN(new_n995));
  INV_X1    g570(.A(new_n992), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n972), .B1(new_n996), .B2(new_n985), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT43), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n987), .A4(new_n993), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n995), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n993), .A2(new_n987), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n990), .A2(new_n992), .B1(new_n970), .B2(new_n971), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT43), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n986), .A2(new_n998), .A3(new_n987), .A4(new_n993), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1004), .B1(new_n1009), .B2(new_n966), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1003), .B1(new_n1010), .B2(new_n1011), .ZN(G397));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n490), .B2(new_n494), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n461), .A2(new_n476), .A3(new_n470), .A4(G40), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n826), .B(G2067), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n888), .A2(G1996), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(KEYINPUT109), .A3(new_n844), .A4(new_n841), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1018), .A2(new_n844), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n888), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1022), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n749), .B(new_n751), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  OR2_X1    g604(.A1(G290), .A2(G1986), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G290), .A2(G1986), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1019), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1033), .B(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G286), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1015), .A2(G1384), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n490), .B2(new_n494), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n1038), .C1(new_n490), .C2(new_n494), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1017), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1966), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1017), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n1013), .C1(new_n490), .C2(new_n494), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT115), .B(G2084), .ZN(new_n1050));
  AND4_X1   g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1037), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT51), .B1(new_n1037), .B2(new_n1054), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1053), .A2(new_n1036), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1053), .B2(new_n1036), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1052), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n1052), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G303), .A2(G8), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT55), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1971), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n805), .A2(new_n1047), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1064), .B(G8), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1063), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1070));
  INV_X1    g645(.A(G1976), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n583), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT111), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1075), .B(KEYINPUT52), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G288), .A2(new_n1071), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1070), .A2(new_n1072), .A3(KEYINPUT52), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1074), .A2(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT49), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G305), .A2(G1981), .ZN(new_n1081));
  INV_X1    g656(.A(G1981), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1082), .B1(new_n703), .B2(new_n588), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n707), .A2(new_n1082), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1083), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(KEYINPUT49), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1070), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1067), .A2(new_n1069), .A3(new_n1079), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1044), .A2(new_n796), .A3(new_n1039), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1047), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n811), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1043), .A2(new_n1044), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1059), .A2(new_n1061), .A3(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1068), .A2(new_n1063), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1101), .A2(new_n1079), .A3(new_n1089), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1084), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT112), .B1(G288), .B2(G1976), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT77), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n583), .B(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1071), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1085), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT113), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1070), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(KEYINPUT113), .B(new_n1085), .C1(new_n1103), .C2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1102), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1069), .A2(new_n1079), .A3(new_n1089), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1069), .A2(new_n1079), .A3(KEYINPUT117), .A4(new_n1089), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  OAI211_X1 g694(.A(G8), .B(G168), .C1(new_n1045), .C2(new_n1051), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1101), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1090), .B2(new_n1120), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1100), .A2(new_n1114), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1090), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G301), .B(KEYINPUT54), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1017), .B(KEYINPUT124), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1129), .A2(new_n1039), .A3(new_n1095), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1130), .B2(new_n1016), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1131), .A2(new_n1094), .B1(new_n1097), .B2(new_n1128), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1058), .A2(new_n1127), .A3(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1014), .A2(G2067), .A3(new_n1017), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1093), .B2(new_n763), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n614), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(new_n815), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1016), .A2(new_n1046), .A3(new_n844), .A4(new_n1039), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT121), .B(new_n1139), .C1(new_n1014), .C2(new_n1017), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1145), .A2(new_n1146), .A3(new_n552), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1146), .B1(new_n1145), .B2(new_n552), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1137), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1135), .A2(new_n613), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n613), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1136), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT56), .B(G2072), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1044), .A2(new_n1039), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(G1956), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1093), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1044), .A2(KEYINPUT119), .A3(new_n1039), .A4(new_n1155), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT57), .B1(new_n567), .B2(KEYINPUT118), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(G299), .Z(new_n1164));
  AND2_X1   g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1154), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT122), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1162), .A2(new_n1168), .A3(new_n1164), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT61), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1153), .B(new_n1167), .C1(new_n1169), .C2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1166), .A2(new_n1150), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1173), .A2(new_n1165), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1133), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1035), .B1(new_n1126), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1030), .A2(new_n1019), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1025), .B(KEYINPUT46), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT47), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1020), .A2(new_n841), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1018), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1180), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1029), .A2(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n742), .A2(new_n744), .A3(new_n751), .A4(new_n748), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT125), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1027), .A2(new_n1187), .ZN(new_n1188));
  OR3_X1    g763(.A1(new_n821), .A2(G2067), .A3(new_n825), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1019), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OR3_X1    g765(.A1(new_n1185), .A2(new_n1190), .A3(KEYINPUT126), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n1185), .B2(new_n1190), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g769(.A(G319), .B1(new_n657), .B2(new_n658), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G227), .A2(new_n1196), .ZN(new_n1197));
  OR2_X1    g771(.A1(new_n1197), .A2(KEYINPUT127), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1197), .A2(KEYINPUT127), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n697), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n908), .B2(new_n914), .ZN(new_n1201));
  AND2_X1   g775(.A1(new_n1201), .A2(new_n1009), .ZN(G308));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1009), .ZN(G225));
endmodule


