

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830;

  XNOR2_X1 U377 ( .A(n477), .B(n608), .ZN(n830) );
  AND2_X1 U378 ( .A1(n599), .A2(n768), .ZN(n773) );
  XNOR2_X1 U379 ( .A(n496), .B(G953), .ZN(n500) );
  BUF_X1 U380 ( .A(n500), .Z(n550) );
  NAND2_X1 U381 ( .A1(n619), .A2(n799), .ZN(n477) );
  XNOR2_X1 U382 ( .A(n614), .B(n446), .ZN(n467) );
  XOR2_X1 U383 ( .A(n600), .B(KEYINPUT103), .Z(n354) );
  AND2_X1 U384 ( .A1(n433), .A2(n467), .ZN(n355) );
  XNOR2_X1 U385 ( .A(n660), .B(KEYINPUT33), .ZN(n356) );
  XNOR2_X1 U386 ( .A(n543), .B(G472), .ZN(n357) );
  AND2_X4 U387 ( .A1(n689), .A2(n688), .ZN(n737) );
  XNOR2_X2 U388 ( .A(n566), .B(n824), .ZN(n740) );
  XNOR2_X2 U389 ( .A(n386), .B(n576), .ZN(n622) );
  AND2_X2 U390 ( .A1(n359), .A2(n646), .ZN(n686) );
  NOR2_X2 U391 ( .A1(n690), .A2(G902), .ZN(n544) );
  NOR2_X1 U392 ( .A1(G953), .A2(G237), .ZN(n583) );
  NAND2_X1 U393 ( .A1(G234), .A2(G237), .ZN(n518) );
  XNOR2_X1 U394 ( .A(n604), .B(n374), .ZN(n659) );
  BUF_X1 U395 ( .A(n550), .Z(n707) );
  XNOR2_X1 U396 ( .A(n704), .B(G146), .ZN(n529) );
  NOR2_X1 U397 ( .A1(n766), .A2(n639), .ZN(n414) );
  AND2_X1 U398 ( .A1(n402), .A2(n400), .ZN(n399) );
  AND2_X1 U399 ( .A1(n398), .A2(n397), .ZN(n396) );
  INV_X1 U400 ( .A(n403), .ZN(n407) );
  AND2_X1 U401 ( .A1(n638), .A2(n373), .ZN(n766) );
  NOR2_X1 U402 ( .A1(n753), .A2(n627), .ZN(n639) );
  XNOR2_X1 U403 ( .A(n410), .B(n356), .ZN(n790) );
  NAND2_X1 U404 ( .A1(n440), .A2(n441), .ZN(n406) );
  NAND2_X1 U405 ( .A1(n443), .A2(n442), .ZN(n403) );
  NOR2_X1 U406 ( .A1(n659), .A2(n358), .ZN(n371) );
  OR2_X1 U407 ( .A1(n771), .A2(n358), .ZN(n672) );
  AND2_X1 U408 ( .A1(n652), .A2(n405), .ZN(n404) );
  INV_X1 U409 ( .A(n771), .ZN(n409) );
  NAND2_X1 U410 ( .A1(n622), .A2(n621), .ZN(n760) );
  NAND2_X1 U411 ( .A1(n622), .A2(n612), .ZN(n593) );
  XNOR2_X1 U412 ( .A(n559), .B(n498), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n501), .B(n417), .ZN(n502) );
  INV_X1 U414 ( .A(KEYINPUT101), .ZN(n385) );
  INV_X1 U415 ( .A(KEYINPUT34), .ZN(n376) );
  INV_X1 U416 ( .A(KEYINPUT8), .ZN(n417) );
  INV_X1 U417 ( .A(KEYINPUT1), .ZN(n374) );
  XNOR2_X1 U418 ( .A(n408), .B(n683), .ZN(n805) );
  NAND2_X1 U419 ( .A1(n388), .A2(n665), .ZN(n387) );
  AND2_X1 U420 ( .A1(n391), .A2(n682), .ZN(n390) );
  XNOR2_X1 U421 ( .A(n686), .B(KEYINPUT86), .ZN(n424) );
  XNOR2_X1 U422 ( .A(n484), .B(n487), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n436), .B(KEYINPUT88), .ZN(n666) );
  NAND2_X1 U424 ( .A1(n700), .A2(n701), .ZN(n436) );
  NAND2_X1 U425 ( .A1(n437), .A2(n462), .ZN(n701) );
  NAND2_X1 U426 ( .A1(n439), .A2(n438), .ZN(n700) );
  XNOR2_X1 U427 ( .A(n663), .B(n662), .ZN(n729) );
  AND2_X1 U428 ( .A1(n454), .A2(n457), .ZN(n439) );
  XNOR2_X1 U429 ( .A(n469), .B(G131), .ZN(G33) );
  XNOR2_X1 U430 ( .A(n377), .B(n376), .ZN(n375) );
  AND2_X2 U431 ( .A1(n473), .A2(n470), .ZN(n469) );
  NAND2_X1 U432 ( .A1(n467), .A2(n466), .ZN(n415) );
  NAND2_X2 U433 ( .A1(n399), .A2(n396), .ZN(n657) );
  NAND2_X1 U434 ( .A1(n472), .A2(n471), .ZN(n470) );
  AND2_X1 U435 ( .A1(n475), .A2(n474), .ZN(n473) );
  AND2_X1 U436 ( .A1(n625), .A2(n624), .ZN(n466) );
  NAND2_X1 U437 ( .A1(n394), .A2(n406), .ZN(n398) );
  NAND2_X1 U438 ( .A1(n404), .A2(n403), .ZN(n402) );
  AND2_X1 U439 ( .A1(n443), .A2(n395), .ZN(n394) );
  NOR2_X1 U440 ( .A1(n782), .A2(n781), .ZN(n787) );
  NOR2_X1 U441 ( .A1(n606), .A2(n605), .ZN(n619) );
  AND2_X1 U442 ( .A1(n549), .A2(n548), .ZN(n609) );
  NOR2_X1 U443 ( .A1(n677), .A2(n409), .ZN(n678) );
  BUF_X1 U444 ( .A(n659), .Z(n370) );
  XNOR2_X1 U445 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U446 ( .A(n360), .B(G469), .ZN(n637) );
  INV_X1 U447 ( .A(n773), .ZN(n358) );
  XNOR2_X1 U448 ( .A(n721), .B(n723), .ZN(n724) );
  INV_X1 U449 ( .A(n760), .ZN(n757) );
  AND2_X1 U450 ( .A1(n442), .A2(n491), .ZN(n395) );
  NOR2_X1 U451 ( .A1(n622), .A2(n612), .ZN(n661) );
  XNOR2_X1 U452 ( .A(n361), .B(n529), .ZN(n720) );
  XNOR2_X1 U453 ( .A(n542), .B(n541), .ZN(n690) );
  AND2_X1 U454 ( .A1(n447), .A2(n520), .ZN(n521) );
  XNOR2_X1 U455 ( .A(n715), .B(KEYINPUT59), .ZN(n716) );
  XNOR2_X1 U456 ( .A(n382), .B(n379), .ZN(n572) );
  NAND2_X1 U457 ( .A1(n429), .A2(n482), .ZN(n435) );
  XNOR2_X1 U458 ( .A(n384), .B(n383), .ZN(n382) );
  XNOR2_X1 U459 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U460 ( .A(n535), .B(KEYINPUT74), .ZN(n495) );
  XNOR2_X1 U461 ( .A(n385), .B(G122), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n555), .B(G134), .ZN(n573) );
  XNOR2_X1 U463 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U464 ( .A(n393), .B(KEYINPUT23), .ZN(n504) );
  XNOR2_X1 U465 ( .A(KEYINPUT16), .B(G122), .ZN(n564) );
  XNOR2_X1 U466 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n380) );
  XNOR2_X1 U467 ( .A(G902), .B(KEYINPUT15), .ZN(n684) );
  XNOR2_X1 U468 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n381) );
  XNOR2_X1 U469 ( .A(G128), .B(G119), .ZN(n393) );
  INV_X1 U470 ( .A(KEYINPUT76), .ZN(n416) );
  XNOR2_X1 U471 ( .A(G116), .B(G107), .ZN(n383) );
  XNOR2_X1 U472 ( .A(G128), .B(G143), .ZN(n555) );
  NOR2_X1 U473 ( .A1(n693), .A2(n743), .ZN(n695) );
  NOR2_X1 U474 ( .A1(n726), .A2(n743), .ZN(n727) );
  NOR2_X1 U475 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U476 ( .A1(n718), .A2(n743), .ZN(n719) );
  XNOR2_X1 U477 ( .A(n424), .B(KEYINPUT76), .ZN(n366) );
  NAND2_X1 U478 ( .A1(n720), .A2(n588), .ZN(n360) );
  NAND2_X1 U479 ( .A1(n362), .A2(n368), .ZN(n689) );
  NAND2_X1 U480 ( .A1(n364), .A2(n363), .ZN(n362) );
  NAND2_X1 U481 ( .A1(n365), .A2(KEYINPUT84), .ZN(n363) );
  NAND2_X1 U482 ( .A1(n366), .A2(n367), .ZN(n364) );
  XNOR2_X1 U483 ( .A(n702), .B(n416), .ZN(n365) );
  INV_X1 U484 ( .A(n483), .ZN(n367) );
  NAND2_X1 U485 ( .A1(n369), .A2(n479), .ZN(n368) );
  OR2_X1 U486 ( .A1(n805), .A2(n435), .ZN(n369) );
  OR2_X1 U487 ( .A1(n659), .A2(n354), .ZN(n372) );
  AND2_X1 U488 ( .A1(n370), .A2(n358), .ZN(n774) );
  NOR2_X1 U489 ( .A1(n370), .A2(n672), .ZN(n777) );
  AND2_X1 U490 ( .A1(n354), .A2(n370), .ZN(n670) );
  INV_X1 U491 ( .A(n370), .ZN(n373) );
  NAND2_X1 U492 ( .A1(n375), .A2(n661), .ZN(n663) );
  NAND2_X1 U493 ( .A1(n790), .A2(n679), .ZN(n377) );
  NAND2_X1 U494 ( .A1(n378), .A2(n419), .ZN(n421) );
  INV_X1 U495 ( .A(n495), .ZN(n378) );
  XNOR2_X2 U496 ( .A(n492), .B(G101), .ZN(n535) );
  NAND2_X1 U497 ( .A1(n735), .A2(n588), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n390), .A2(n387), .ZN(n408) );
  NAND2_X1 U499 ( .A1(n389), .A2(n664), .ZN(n388) );
  NAND2_X1 U500 ( .A1(n666), .A2(KEYINPUT66), .ZN(n389) );
  NAND2_X1 U501 ( .A1(n392), .A2(n669), .ZN(n391) );
  INV_X1 U502 ( .A(n666), .ZN(n392) );
  NAND2_X1 U503 ( .A1(n407), .A2(n406), .ZN(n679) );
  OR2_X1 U504 ( .A1(n652), .A2(n405), .ZN(n397) );
  NAND2_X1 U505 ( .A1(n404), .A2(n401), .ZN(n400) );
  INV_X1 U506 ( .A(n406), .ZN(n401) );
  INV_X1 U507 ( .A(n491), .ZN(n405) );
  NOR2_X1 U508 ( .A1(n771), .A2(n781), .ZN(n547) );
  NAND2_X1 U509 ( .A1(n601), .A2(n409), .ZN(n603) );
  XNOR2_X2 U510 ( .A(n544), .B(n357), .ZN(n771) );
  NAND2_X1 U511 ( .A1(n654), .A2(n371), .ZN(n410) );
  NAND2_X1 U512 ( .A1(n412), .A2(n411), .ZN(n486) );
  NAND2_X1 U513 ( .A1(n355), .A2(n414), .ZN(n411) );
  NAND2_X1 U514 ( .A1(n413), .A2(n415), .ZN(n412) );
  AND2_X1 U515 ( .A1(n414), .A2(KEYINPUT81), .ZN(n413) );
  INV_X1 U516 ( .A(n805), .ZN(n480) );
  NAND2_X1 U517 ( .A1(n502), .A2(G217), .ZN(n574) );
  BUF_X1 U518 ( .A(n631), .Z(n418) );
  NAND2_X1 U519 ( .A1(n495), .A2(n494), .ZN(n420) );
  NAND2_X1 U520 ( .A1(n420), .A2(n421), .ZN(n559) );
  INV_X1 U521 ( .A(n494), .ZN(n419) );
  XNOR2_X1 U522 ( .A(n535), .B(KEYINPUT74), .ZN(n422) );
  BUF_X1 U523 ( .A(n737), .Z(n734) );
  NOR2_X1 U524 ( .A1(n731), .A2(G902), .ZN(n445) );
  INV_X1 U525 ( .A(n472), .ZN(n423) );
  XNOR2_X1 U526 ( .A(n422), .B(n494), .ZN(n425) );
  XNOR2_X1 U527 ( .A(n686), .B(KEYINPUT86), .ZN(n702) );
  BUF_X1 U528 ( .A(n637), .Z(n604) );
  NOR2_X1 U529 ( .A1(n460), .A2(KEYINPUT68), .ZN(n459) );
  NAND2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n490) );
  XNOR2_X1 U531 ( .A(KEYINPUT4), .B(G131), .ZN(n499) );
  XNOR2_X1 U532 ( .A(G137), .B(G140), .ZN(n507) );
  INV_X1 U533 ( .A(KEYINPUT48), .ZN(n487) );
  NAND2_X1 U534 ( .A1(n372), .A2(n465), .ZN(n464) );
  INV_X1 U535 ( .A(KEYINPUT0), .ZN(n444) );
  XOR2_X1 U536 ( .A(G113), .B(KEYINPUT73), .Z(n533) );
  XNOR2_X1 U537 ( .A(G119), .B(G116), .ZN(n532) );
  INV_X1 U538 ( .A(n811), .ZN(n688) );
  NAND2_X1 U539 ( .A1(n760), .A2(n476), .ZN(n474) );
  NOR2_X1 U540 ( .A1(n372), .A2(n465), .ZN(n463) );
  NAND2_X1 U541 ( .A1(n464), .A2(n428), .ZN(n461) );
  NOR2_X1 U542 ( .A1(n656), .A2(n478), .ZN(n458) );
  NOR2_X1 U543 ( .A1(n707), .A2(G952), .ZN(n743) );
  NAND2_X1 U544 ( .A1(n482), .A2(KEYINPUT84), .ZN(n481) );
  NAND2_X1 U545 ( .A1(n429), .A2(KEYINPUT84), .ZN(n479) );
  INV_X1 U546 ( .A(G237), .ZN(n545) );
  INV_X1 U547 ( .A(KEYINPUT38), .ZN(n451) );
  INV_X1 U548 ( .A(G902), .ZN(n588) );
  XNOR2_X1 U549 ( .A(G110), .B(KEYINPUT24), .ZN(n503) );
  XOR2_X1 U550 ( .A(G104), .B(G143), .Z(n578) );
  XNOR2_X1 U551 ( .A(G113), .B(G131), .ZN(n577) );
  XNOR2_X1 U552 ( .A(G122), .B(G140), .ZN(n579) );
  XNOR2_X1 U553 ( .A(n603), .B(n602), .ZN(n606) );
  XNOR2_X1 U554 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n602) );
  XNOR2_X1 U555 ( .A(n690), .B(KEYINPUT62), .ZN(n691) );
  INV_X1 U556 ( .A(G953), .ZN(n818) );
  NAND2_X1 U557 ( .A1(n645), .A2(n452), .ZN(n696) );
  NOR2_X1 U558 ( .A1(n760), .A2(n476), .ZN(n471) );
  NAND2_X1 U559 ( .A1(n453), .A2(n461), .ZN(n437) );
  INV_X1 U560 ( .A(KEYINPUT109), .ZN(n446) );
  NAND2_X1 U561 ( .A1(n456), .A2(KEYINPUT68), .ZN(n438) );
  NOR2_X1 U562 ( .A1(n458), .A2(n600), .ZN(n457) );
  XNOR2_X1 U563 ( .A(n450), .B(n449), .ZN(n736) );
  INV_X1 U564 ( .A(n735), .ZN(n449) );
  NAND2_X1 U565 ( .A1(n734), .A2(G478), .ZN(n450) );
  XNOR2_X1 U566 ( .A(n651), .B(KEYINPUT95), .ZN(n426) );
  AND2_X1 U567 ( .A1(n624), .A2(n488), .ZN(n427) );
  XOR2_X1 U568 ( .A(n655), .B(KEYINPUT32), .Z(n428) );
  NAND2_X1 U569 ( .A1(n685), .A2(KEYINPUT2), .ZN(n429) );
  XOR2_X1 U570 ( .A(n568), .B(KEYINPUT92), .Z(n430) );
  XOR2_X1 U571 ( .A(n514), .B(n513), .Z(n431) );
  NAND2_X1 U572 ( .A1(n657), .A2(n658), .ZN(n432) );
  XNOR2_X1 U573 ( .A(n617), .B(n616), .ZN(n618) );
  AND2_X1 U574 ( .A1(n625), .A2(n427), .ZN(n433) );
  AND2_X1 U575 ( .A1(n464), .A2(n658), .ZN(n434) );
  INV_X1 U576 ( .A(KEYINPUT68), .ZN(n478) );
  INV_X1 U577 ( .A(n428), .ZN(n465) );
  INV_X1 U578 ( .A(KEYINPUT81), .ZN(n488) );
  INV_X1 U579 ( .A(n618), .ZN(n440) );
  NOR2_X1 U580 ( .A1(n426), .A2(n444), .ZN(n441) );
  NAND2_X1 U581 ( .A1(n426), .A2(n444), .ZN(n442) );
  NAND2_X1 U582 ( .A1(n618), .A2(n444), .ZN(n443) );
  XNOR2_X1 U583 ( .A(n445), .B(n431), .ZN(n599) );
  INV_X1 U584 ( .A(n830), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n490), .B(n489), .ZN(n485) );
  INV_X1 U586 ( .A(n467), .ZN(n730) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT104), .ZN(n447) );
  XNOR2_X1 U588 ( .A(n448), .B(n598), .ZN(n630) );
  NOR2_X1 U589 ( .A1(n596), .A2(n597), .ZN(n448) );
  NOR2_X1 U590 ( .A1(n524), .A2(n650), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n631), .B(n451), .ZN(n591) );
  INV_X1 U592 ( .A(n418), .ZN(n452) );
  XNOR2_X2 U593 ( .A(n569), .B(n430), .ZN(n631) );
  NAND2_X1 U594 ( .A1(n657), .A2(n434), .ZN(n453) );
  NAND2_X1 U595 ( .A1(n657), .A2(n459), .ZN(n454) );
  NAND2_X1 U596 ( .A1(n657), .A2(n455), .ZN(n462) );
  AND2_X1 U597 ( .A1(n463), .A2(n658), .ZN(n455) );
  INV_X1 U598 ( .A(n657), .ZN(n456) );
  INV_X1 U599 ( .A(n656), .ZN(n460) );
  INV_X1 U600 ( .A(n640), .ZN(n472) );
  NAND2_X1 U601 ( .A1(n640), .A2(n476), .ZN(n475) );
  INV_X1 U602 ( .A(KEYINPUT40), .ZN(n476) );
  XNOR2_X2 U603 ( .A(n571), .B(n570), .ZN(n640) );
  XNOR2_X2 U604 ( .A(n594), .B(n595), .ZN(n799) );
  NAND2_X1 U605 ( .A1(n486), .A2(n485), .ZN(n484) );
  NOR2_X1 U606 ( .A1(n805), .A2(n481), .ZN(n483) );
  INV_X1 U607 ( .A(n684), .ZN(n482) );
  INV_X1 U608 ( .A(KEYINPUT46), .ZN(n489) );
  XOR2_X1 U609 ( .A(n653), .B(KEYINPUT22), .Z(n491) );
  INV_X1 U610 ( .A(KEYINPUT63), .ZN(n694) );
  XNOR2_X2 U611 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n492) );
  XNOR2_X1 U612 ( .A(G104), .B(G110), .ZN(n493) );
  XNOR2_X1 U613 ( .A(n493), .B(G107), .ZN(n823) );
  INV_X1 U614 ( .A(n823), .ZN(n494) );
  INV_X2 U615 ( .A(KEYINPUT64), .ZN(n496) );
  NAND2_X1 U616 ( .A1(n707), .A2(G227), .ZN(n497) );
  XNOR2_X1 U617 ( .A(n497), .B(n507), .ZN(n498) );
  XNOR2_X2 U618 ( .A(n573), .B(n499), .ZN(n704) );
  NAND2_X1 U619 ( .A1(n500), .A2(G234), .ZN(n501) );
  NAND2_X1 U620 ( .A1(n502), .A2(G221), .ZN(n506) );
  XNOR2_X1 U621 ( .A(n506), .B(n505), .ZN(n508) );
  XNOR2_X1 U622 ( .A(G146), .B(G125), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n554), .B(KEYINPUT10), .ZN(n585) );
  XNOR2_X1 U624 ( .A(n585), .B(n507), .ZN(n706) );
  XNOR2_X1 U625 ( .A(n508), .B(n706), .ZN(n731) );
  NAND2_X1 U626 ( .A1(n684), .A2(G234), .ZN(n510) );
  INV_X1 U627 ( .A(KEYINPUT20), .ZN(n509) );
  XNOR2_X1 U628 ( .A(n510), .B(n509), .ZN(n516) );
  INV_X1 U629 ( .A(n516), .ZN(n511) );
  NAND2_X1 U630 ( .A1(n511), .A2(G217), .ZN(n514) );
  XNOR2_X1 U631 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n512) );
  XNOR2_X1 U632 ( .A(n512), .B(KEYINPUT25), .ZN(n513) );
  INV_X1 U633 ( .A(G221), .ZN(n515) );
  OR2_X1 U634 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U635 ( .A(n517), .B(KEYINPUT21), .ZN(n597) );
  INV_X1 U636 ( .A(n597), .ZN(n768) );
  NAND2_X1 U637 ( .A1(n637), .A2(n773), .ZN(n676) );
  XNOR2_X1 U638 ( .A(n676), .B(KEYINPUT107), .ZN(n527) );
  XNOR2_X1 U639 ( .A(n518), .B(KEYINPUT14), .ZN(n522) );
  NAND2_X1 U640 ( .A1(n522), .A2(G902), .ZN(n647) );
  NOR2_X1 U641 ( .A1(n647), .A2(n550), .ZN(n519) );
  INV_X1 U642 ( .A(G900), .ZN(n520) );
  XOR2_X1 U643 ( .A(KEYINPUT105), .B(n521), .Z(n524) );
  NAND2_X1 U644 ( .A1(n522), .A2(G952), .ZN(n523) );
  XNOR2_X1 U645 ( .A(n523), .B(KEYINPUT94), .ZN(n797) );
  NOR2_X1 U646 ( .A1(G953), .A2(n797), .ZN(n650) );
  XNOR2_X1 U647 ( .A(n525), .B(KEYINPUT80), .ZN(n596) );
  INV_X1 U648 ( .A(n596), .ZN(n526) );
  NAND2_X1 U649 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U650 ( .A(n528), .B(KEYINPUT77), .ZN(n549) );
  INV_X1 U651 ( .A(n529), .ZN(n542) );
  INV_X1 U652 ( .A(KEYINPUT91), .ZN(n530) );
  XNOR2_X1 U653 ( .A(n530), .B(KEYINPUT3), .ZN(n531) );
  XNOR2_X1 U654 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U655 ( .A(n534), .B(n533), .ZN(n565) );
  NAND2_X1 U656 ( .A1(n583), .A2(G210), .ZN(n536) );
  XNOR2_X1 U657 ( .A(n536), .B(KEYINPUT96), .ZN(n538) );
  XNOR2_X1 U658 ( .A(G137), .B(KEYINPUT5), .ZN(n537) );
  XNOR2_X1 U659 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U660 ( .A(n535), .B(n539), .ZN(n540) );
  XNOR2_X1 U661 ( .A(n565), .B(n540), .ZN(n541) );
  INV_X1 U662 ( .A(KEYINPUT97), .ZN(n543) );
  NAND2_X1 U663 ( .A1(n588), .A2(n545), .ZN(n567) );
  NAND2_X1 U664 ( .A1(n567), .A2(G214), .ZN(n546) );
  XNOR2_X1 U665 ( .A(n546), .B(KEYINPUT93), .ZN(n781) );
  INV_X1 U666 ( .A(n781), .ZN(n615) );
  XNOR2_X1 U667 ( .A(n547), .B(KEYINPUT30), .ZN(n548) );
  NAND2_X1 U668 ( .A1(n550), .A2(G224), .ZN(n553) );
  XNOR2_X1 U669 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n551) );
  XNOR2_X1 U670 ( .A(n551), .B(KEYINPUT4), .ZN(n552) );
  XNOR2_X1 U671 ( .A(n553), .B(n552), .ZN(n557) );
  XNOR2_X1 U672 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U673 ( .A(n557), .B(n556), .ZN(n560) );
  INV_X1 U674 ( .A(n560), .ZN(n558) );
  NAND2_X1 U675 ( .A1(n558), .A2(n425), .ZN(n563) );
  INV_X1 U676 ( .A(n425), .ZN(n561) );
  NAND2_X1 U677 ( .A1(n560), .A2(n561), .ZN(n562) );
  NAND2_X1 U678 ( .A1(n563), .A2(n562), .ZN(n566) );
  XNOR2_X1 U679 ( .A(n565), .B(n564), .ZN(n824) );
  NAND2_X1 U680 ( .A1(n740), .A2(n684), .ZN(n569) );
  NAND2_X1 U681 ( .A1(n567), .A2(G210), .ZN(n568) );
  NAND2_X1 U682 ( .A1(n609), .A2(n591), .ZN(n571) );
  INV_X1 U683 ( .A(KEYINPUT39), .ZN(n570) );
  XNOR2_X1 U684 ( .A(n573), .B(n572), .ZN(n575) );
  XNOR2_X1 U685 ( .A(n575), .B(n574), .ZN(n735) );
  INV_X1 U686 ( .A(G478), .ZN(n576) );
  XNOR2_X1 U687 ( .A(n578), .B(n577), .ZN(n582) );
  XOR2_X1 U688 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n580) );
  XNOR2_X1 U689 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U690 ( .A(n582), .B(n581), .Z(n587) );
  AND2_X1 U691 ( .A1(n583), .A2(G214), .ZN(n584) );
  XNOR2_X1 U692 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U693 ( .A(n587), .B(n586), .ZN(n715) );
  NAND2_X1 U694 ( .A1(n715), .A2(n588), .ZN(n590) );
  XNOR2_X1 U695 ( .A(KEYINPUT13), .B(G475), .ZN(n589) );
  XNOR2_X1 U696 ( .A(n590), .B(n589), .ZN(n612) );
  INV_X1 U697 ( .A(n612), .ZN(n621) );
  XOR2_X1 U698 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n595) );
  INV_X1 U699 ( .A(n591), .ZN(n782) );
  INV_X1 U700 ( .A(KEYINPUT102), .ZN(n592) );
  XNOR2_X1 U701 ( .A(n593), .B(n592), .ZN(n784) );
  NAND2_X1 U702 ( .A1(n787), .A2(n784), .ZN(n594) );
  INV_X1 U703 ( .A(KEYINPUT72), .ZN(n598) );
  BUF_X1 U704 ( .A(n599), .Z(n600) );
  NOR2_X1 U705 ( .A1(n630), .A2(n600), .ZN(n601) );
  INV_X1 U706 ( .A(n604), .ZN(n605) );
  INV_X1 U707 ( .A(KEYINPUT112), .ZN(n607) );
  XNOR2_X1 U708 ( .A(n607), .B(KEYINPUT42), .ZN(n608) );
  NAND2_X1 U709 ( .A1(n609), .A2(n418), .ZN(n611) );
  INV_X1 U710 ( .A(KEYINPUT108), .ZN(n610) );
  XNOR2_X1 U711 ( .A(n611), .B(n610), .ZN(n613) );
  NAND2_X1 U712 ( .A1(n613), .A2(n661), .ZN(n614) );
  NAND2_X1 U713 ( .A1(n631), .A2(n615), .ZN(n617) );
  INV_X1 U714 ( .A(KEYINPUT19), .ZN(n616) );
  NAND2_X1 U715 ( .A1(n619), .A2(n440), .ZN(n753) );
  NAND2_X1 U716 ( .A1(n753), .A2(KEYINPUT47), .ZN(n620) );
  XNOR2_X1 U717 ( .A(n620), .B(KEYINPUT82), .ZN(n625) );
  OR2_X1 U718 ( .A1(n622), .A2(n621), .ZN(n762) );
  NAND2_X1 U719 ( .A1(n760), .A2(n762), .ZN(n786) );
  INV_X1 U720 ( .A(n786), .ZN(n623) );
  NAND2_X1 U721 ( .A1(n623), .A2(KEYINPUT47), .ZN(n624) );
  INV_X1 U722 ( .A(KEYINPUT47), .ZN(n626) );
  NAND2_X1 U723 ( .A1(n786), .A2(n626), .ZN(n627) );
  NOR2_X1 U724 ( .A1(n600), .A2(n781), .ZN(n628) );
  NAND2_X1 U725 ( .A1(n757), .A2(n628), .ZN(n629) );
  NOR2_X1 U726 ( .A1(n630), .A2(n629), .ZN(n641) );
  AND2_X1 U727 ( .A1(n418), .A2(n641), .ZN(n632) );
  XNOR2_X1 U728 ( .A(n771), .B(KEYINPUT6), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n632), .A2(n654), .ZN(n636) );
  XNOR2_X1 U730 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n634) );
  INV_X1 U731 ( .A(KEYINPUT113), .ZN(n633) );
  XNOR2_X1 U732 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U733 ( .A(n636), .B(n635), .ZN(n638) );
  OR2_X1 U734 ( .A1(n423), .A2(n762), .ZN(n698) );
  AND2_X1 U735 ( .A1(n654), .A2(n641), .ZN(n642) );
  NAND2_X1 U736 ( .A1(n642), .A2(n659), .ZN(n644) );
  XNOR2_X1 U737 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n643) );
  XNOR2_X1 U738 ( .A(n644), .B(n643), .ZN(n645) );
  AND2_X1 U739 ( .A1(n698), .A2(n696), .ZN(n646) );
  INV_X1 U740 ( .A(n647), .ZN(n648) );
  NOR2_X1 U741 ( .A1(G898), .A2(n818), .ZN(n827) );
  AND2_X1 U742 ( .A1(n648), .A2(n827), .ZN(n649) );
  OR2_X1 U743 ( .A1(n650), .A2(n649), .ZN(n651) );
  AND2_X1 U744 ( .A1(n784), .A2(n768), .ZN(n652) );
  INV_X1 U745 ( .A(KEYINPUT69), .ZN(n653) );
  INV_X1 U746 ( .A(n654), .ZN(n658) );
  INV_X1 U747 ( .A(KEYINPUT67), .ZN(n655) );
  AND2_X1 U748 ( .A1(n659), .A2(n771), .ZN(n656) );
  INV_X1 U749 ( .A(KEYINPUT75), .ZN(n660) );
  INV_X1 U750 ( .A(KEYINPUT35), .ZN(n662) );
  AND2_X1 U751 ( .A1(n729), .A2(KEYINPUT44), .ZN(n664) );
  INV_X1 U752 ( .A(KEYINPUT44), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n667), .A2(KEYINPUT66), .ZN(n665) );
  NAND2_X1 U754 ( .A1(n729), .A2(n667), .ZN(n668) );
  NAND2_X1 U755 ( .A1(n668), .A2(KEYINPUT66), .ZN(n669) );
  XNOR2_X1 U756 ( .A(n432), .B(KEYINPUT87), .ZN(n671) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n746) );
  NAND2_X1 U758 ( .A1(n679), .A2(n777), .ZN(n675) );
  INV_X1 U759 ( .A(KEYINPUT98), .ZN(n673) );
  XNOR2_X1 U760 ( .A(n673), .B(KEYINPUT31), .ZN(n674) );
  XNOR2_X1 U761 ( .A(n675), .B(n674), .ZN(n763) );
  BUF_X1 U762 ( .A(n676), .Z(n677) );
  NAND2_X1 U763 ( .A1(n679), .A2(n678), .ZN(n750) );
  NAND2_X1 U764 ( .A1(n763), .A2(n750), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n680), .A2(n786), .ZN(n681) );
  AND2_X1 U766 ( .A1(n746), .A2(n681), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n683) );
  XNOR2_X1 U768 ( .A(n684), .B(KEYINPUT85), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n686), .A2(KEYINPUT2), .ZN(n687) );
  NOR2_X1 U770 ( .A1(n805), .A2(n687), .ZN(n811) );
  NAND2_X1 U771 ( .A1(n737), .A2(G472), .ZN(n692) );
  XNOR2_X1 U772 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U773 ( .A(n695), .B(n694), .ZN(G57) );
  XNOR2_X1 U774 ( .A(n696), .B(G140), .ZN(G42) );
  XOR2_X1 U775 ( .A(G134), .B(KEYINPUT117), .Z(n697) );
  XNOR2_X1 U776 ( .A(n698), .B(n697), .ZN(G36) );
  XOR2_X1 U777 ( .A(G110), .B(KEYINPUT115), .Z(n699) );
  XNOR2_X1 U778 ( .A(n700), .B(n699), .ZN(G12) );
  XNOR2_X1 U779 ( .A(n701), .B(G119), .ZN(G21) );
  BUF_X1 U780 ( .A(n424), .Z(n703) );
  XNOR2_X1 U781 ( .A(n704), .B(KEYINPUT125), .ZN(n705) );
  XOR2_X1 U782 ( .A(n706), .B(n705), .Z(n709) );
  XNOR2_X1 U783 ( .A(n703), .B(n709), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n708), .A2(n707), .ZN(n714) );
  XOR2_X1 U785 ( .A(n709), .B(KEYINPUT126), .Z(n710) );
  XNOR2_X1 U786 ( .A(G227), .B(n710), .ZN(n711) );
  NAND2_X1 U787 ( .A1(G900), .A2(n711), .ZN(n712) );
  NAND2_X1 U788 ( .A1(n712), .A2(G953), .ZN(n713) );
  NAND2_X1 U789 ( .A1(n714), .A2(n713), .ZN(G72) );
  NAND2_X1 U790 ( .A1(n737), .A2(G475), .ZN(n717) );
  XNOR2_X1 U791 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U792 ( .A(n719), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U793 ( .A1(n737), .A2(G469), .ZN(n725) );
  BUF_X1 U794 ( .A(n720), .Z(n721) );
  XOR2_X1 U795 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n722) );
  XNOR2_X1 U796 ( .A(n722), .B(KEYINPUT58), .ZN(n723) );
  XNOR2_X1 U797 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U798 ( .A(n727), .B(KEYINPUT124), .ZN(G54) );
  XOR2_X1 U799 ( .A(G122), .B(KEYINPUT127), .Z(n728) );
  XNOR2_X1 U800 ( .A(n729), .B(n728), .ZN(G24) );
  XOR2_X1 U801 ( .A(n730), .B(G143), .Z(G45) );
  NAND2_X1 U802 ( .A1(n734), .A2(G217), .ZN(n732) );
  XNOR2_X1 U803 ( .A(n731), .B(n732), .ZN(n733) );
  NOR2_X1 U804 ( .A1(n733), .A2(n743), .ZN(G66) );
  NOR2_X1 U805 ( .A1(n736), .A2(n743), .ZN(G63) );
  NAND2_X1 U806 ( .A1(n737), .A2(G210), .ZN(n742) );
  XNOR2_X1 U807 ( .A(KEYINPUT90), .B(KEYINPUT54), .ZN(n738) );
  XNOR2_X1 U808 ( .A(n738), .B(KEYINPUT55), .ZN(n739) );
  XNOR2_X1 U809 ( .A(n742), .B(n741), .ZN(n744) );
  XNOR2_X1 U810 ( .A(n745), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U811 ( .A(G101), .B(n746), .ZN(G3) );
  NOR2_X1 U812 ( .A1(n750), .A2(n760), .ZN(n747) );
  XOR2_X1 U813 ( .A(G104), .B(n747), .Z(G6) );
  XOR2_X1 U814 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n749) );
  XNOR2_X1 U815 ( .A(G107), .B(KEYINPUT114), .ZN(n748) );
  XNOR2_X1 U816 ( .A(n749), .B(n748), .ZN(n752) );
  NOR2_X1 U817 ( .A1(n750), .A2(n762), .ZN(n751) );
  XOR2_X1 U818 ( .A(n752), .B(n751), .Z(G9) );
  XOR2_X1 U819 ( .A(G128), .B(KEYINPUT29), .Z(n756) );
  INV_X1 U820 ( .A(n753), .ZN(n758) );
  INV_X1 U821 ( .A(n762), .ZN(n754) );
  NAND2_X1 U822 ( .A1(n758), .A2(n754), .ZN(n755) );
  XNOR2_X1 U823 ( .A(n756), .B(n755), .ZN(G30) );
  NAND2_X1 U824 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U825 ( .A(n759), .B(G146), .ZN(G48) );
  NOR2_X1 U826 ( .A1(n763), .A2(n760), .ZN(n761) );
  XOR2_X1 U827 ( .A(G113), .B(n761), .Z(G15) );
  NOR2_X1 U828 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U829 ( .A(KEYINPUT116), .B(n764), .Z(n765) );
  XNOR2_X1 U830 ( .A(G116), .B(n765), .ZN(G18) );
  XNOR2_X1 U831 ( .A(G125), .B(n766), .ZN(n767) );
  XNOR2_X1 U832 ( .A(n767), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U833 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n817) );
  NOR2_X1 U834 ( .A1(n354), .A2(n768), .ZN(n769) );
  XNOR2_X1 U835 ( .A(n769), .B(KEYINPUT49), .ZN(n770) );
  XNOR2_X1 U836 ( .A(n770), .B(KEYINPUT118), .ZN(n772) );
  NAND2_X1 U837 ( .A1(n772), .A2(n771), .ZN(n776) );
  XNOR2_X1 U838 ( .A(n774), .B(KEYINPUT50), .ZN(n775) );
  NOR2_X1 U839 ( .A1(n776), .A2(n775), .ZN(n778) );
  OR2_X1 U840 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U841 ( .A(KEYINPUT51), .B(n779), .Z(n780) );
  NAND2_X1 U842 ( .A1(n799), .A2(n780), .ZN(n793) );
  NAND2_X1 U843 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U844 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U845 ( .A(KEYINPUT119), .B(n785), .Z(n789) );
  NAND2_X1 U846 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U847 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U848 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U849 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U850 ( .A(n794), .B(KEYINPUT52), .Z(n795) );
  XNOR2_X1 U851 ( .A(KEYINPUT120), .B(n795), .ZN(n796) );
  NOR2_X1 U852 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U853 ( .A(n798), .B(KEYINPUT121), .ZN(n801) );
  NAND2_X1 U854 ( .A1(n799), .A2(n790), .ZN(n800) );
  NAND2_X1 U855 ( .A1(n801), .A2(n800), .ZN(n814) );
  INV_X1 U856 ( .A(n703), .ZN(n802) );
  NOR2_X1 U857 ( .A1(n802), .A2(n805), .ZN(n803) );
  NOR2_X1 U858 ( .A1(n803), .A2(KEYINPUT2), .ZN(n804) );
  NOR2_X1 U859 ( .A1(n804), .A2(KEYINPUT83), .ZN(n810) );
  INV_X1 U860 ( .A(KEYINPUT83), .ZN(n806) );
  NOR2_X1 U861 ( .A1(n806), .A2(KEYINPUT2), .ZN(n807) );
  NAND2_X1 U862 ( .A1(n480), .A2(n807), .ZN(n808) );
  NOR2_X1 U863 ( .A1(n703), .A2(n808), .ZN(n809) );
  NOR2_X1 U864 ( .A1(n810), .A2(n809), .ZN(n812) );
  NOR2_X1 U865 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U866 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U867 ( .A1(n815), .A2(n818), .ZN(n816) );
  XNOR2_X1 U868 ( .A(n817), .B(n816), .ZN(G75) );
  NAND2_X1 U869 ( .A1(n480), .A2(n818), .ZN(n822) );
  NAND2_X1 U870 ( .A1(G953), .A2(G224), .ZN(n819) );
  XNOR2_X1 U871 ( .A(KEYINPUT61), .B(n819), .ZN(n820) );
  NAND2_X1 U872 ( .A1(n820), .A2(G898), .ZN(n821) );
  NAND2_X1 U873 ( .A1(n822), .A2(n821), .ZN(n829) );
  XNOR2_X1 U874 ( .A(G101), .B(n823), .ZN(n825) );
  XNOR2_X1 U875 ( .A(n825), .B(n824), .ZN(n826) );
  NOR2_X1 U876 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U877 ( .A(n829), .B(n828), .ZN(G69) );
  XOR2_X1 U878 ( .A(G137), .B(n830), .Z(G39) );
endmodule

