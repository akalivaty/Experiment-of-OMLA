

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U326 ( .A(n346), .B(n358), .ZN(n502) );
  XOR2_X1 U327 ( .A(KEYINPUT38), .B(n453), .Z(n294) );
  NOR2_X1 U328 ( .A1(n549), .A2(n406), .ZN(n407) );
  INV_X1 U329 ( .A(KEYINPUT77), .ZN(n438) );
  XNOR2_X1 U330 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U331 ( .A(n439), .B(n438), .ZN(n448) );
  XOR2_X1 U332 ( .A(G15GAT), .B(G127GAT), .Z(n331) );
  XNOR2_X1 U333 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U334 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n412), .B(KEYINPUT103), .ZN(n413) );
  XNOR2_X1 U336 ( .A(n414), .B(n413), .ZN(n520) );
  NOR2_X1 U337 ( .A1(n502), .A2(n475), .ZN(n565) );
  XNOR2_X1 U338 ( .A(KEYINPUT41), .B(n574), .ZN(n557) );
  INV_X1 U339 ( .A(n502), .ZN(n532) );
  XNOR2_X1 U340 ( .A(n479), .B(G176GAT), .ZN(n480) );
  XNOR2_X1 U341 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n454) );
  XNOR2_X1 U342 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  XNOR2_X1 U343 ( .A(n455), .B(n454), .ZN(G1328GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT82), .B(KEYINPUT10), .Z(n296) );
  XNOR2_X1 U345 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U347 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n298) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(KEYINPUT9), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(n299), .B(G218GAT), .Z(n301) );
  XOR2_X1 U351 ( .A(G43GAT), .B(G134GAT), .Z(n334) );
  XNOR2_X1 U352 ( .A(G190GAT), .B(n334), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U354 ( .A(G85GAT), .B(G92GAT), .Z(n433) );
  XOR2_X1 U355 ( .A(n433), .B(KEYINPUT65), .Z(n303) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(n305), .B(n304), .Z(n311) );
  XOR2_X1 U359 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n307) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U362 ( .A(KEYINPUT7), .B(n308), .Z(n431) );
  INV_X1 U363 ( .A(n431), .ZN(n309) );
  XOR2_X1 U364 ( .A(G50GAT), .B(G162GAT), .Z(n387) );
  XOR2_X1 U365 ( .A(n309), .B(n387), .Z(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n564) );
  XOR2_X1 U368 ( .A(n564), .B(KEYINPUT36), .Z(n583) );
  XNOR2_X1 U369 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n314) );
  XNOR2_X1 U370 ( .A(n314), .B(KEYINPUT13), .ZN(n434) );
  XOR2_X1 U371 ( .A(KEYINPUT83), .B(n434), .Z(n316) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(G22GAT), .B(G155GAT), .Z(n386) );
  XOR2_X1 U375 ( .A(n317), .B(n386), .Z(n320) );
  XNOR2_X1 U376 ( .A(G8GAT), .B(G1GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n318), .B(KEYINPUT71), .ZN(n423) );
  XNOR2_X1 U378 ( .A(n423), .B(n331), .ZN(n319) );
  XNOR2_X1 U379 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U380 ( .A(G211GAT), .B(G78GAT), .Z(n322) );
  XNOR2_X1 U381 ( .A(G183GAT), .B(G71GAT), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U383 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n324) );
  XNOR2_X1 U384 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U387 ( .A(n328), .B(n327), .Z(n579) );
  INV_X1 U388 ( .A(n579), .ZN(n462) );
  XOR2_X1 U389 ( .A(KEYINPUT86), .B(KEYINPUT0), .Z(n330) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n377) );
  XNOR2_X1 U392 ( .A(n331), .B(KEYINPUT20), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n332), .B(KEYINPUT87), .ZN(n336) );
  AND2_X1 U394 ( .A1(G227GAT), .A2(G233GAT), .ZN(n333) );
  XOR2_X1 U395 ( .A(n377), .B(n337), .Z(n339) );
  XOR2_X1 U396 ( .A(G99GAT), .B(G71GAT), .Z(n338) );
  XOR2_X1 U397 ( .A(G120GAT), .B(n338), .Z(n437) );
  XNOR2_X1 U398 ( .A(n339), .B(n437), .ZN(n346) );
  XOR2_X1 U399 ( .A(G176GAT), .B(G183GAT), .Z(n341) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U402 ( .A(KEYINPUT17), .B(KEYINPUT88), .Z(n343) );
  XNOR2_X1 U403 ( .A(G190GAT), .B(KEYINPUT18), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U405 ( .A(n345), .B(n344), .Z(n358) );
  XNOR2_X1 U406 ( .A(n532), .B(KEYINPUT89), .ZN(n401) );
  XOR2_X1 U407 ( .A(G204GAT), .B(KEYINPUT98), .Z(n348) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n351) );
  XNOR2_X1 U410 ( .A(G36GAT), .B(G92GAT), .ZN(n349) );
  XOR2_X1 U411 ( .A(KEYINPUT79), .B(G64GAT), .Z(n444) );
  XNOR2_X1 U412 ( .A(n349), .B(n444), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U414 ( .A(KEYINPUT90), .B(G218GAT), .Z(n353) );
  XNOR2_X1 U415 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U417 ( .A(G197GAT), .B(n354), .Z(n385) );
  XNOR2_X1 U418 ( .A(G8GAT), .B(n385), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U420 ( .A(n358), .B(n357), .Z(n523) );
  XOR2_X1 U421 ( .A(KEYINPUT27), .B(n523), .Z(n403) );
  XOR2_X1 U422 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n360) );
  XNOR2_X1 U423 ( .A(G1GAT), .B(G57GAT), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U425 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n362) );
  XNOR2_X1 U426 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U428 ( .A(n364), .B(n363), .Z(n369) );
  XOR2_X1 U429 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n366) );
  NAND2_X1 U430 ( .A1(G225GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U432 ( .A(KEYINPUT1), .B(n367), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U434 ( .A(G85GAT), .B(G162GAT), .Z(n371) );
  XNOR2_X1 U435 ( .A(G29GAT), .B(G134GAT), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U437 ( .A(G155GAT), .B(G148GAT), .Z(n373) );
  XNOR2_X1 U438 ( .A(G120GAT), .B(G127GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U440 ( .A(n375), .B(n374), .Z(n379) );
  XNOR2_X1 U441 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n376), .B(KEYINPUT2), .ZN(n391) );
  XNOR2_X1 U443 ( .A(n377), .B(n391), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n521) );
  XOR2_X1 U446 ( .A(G148GAT), .B(G106GAT), .Z(n383) );
  XNOR2_X1 U447 ( .A(G204GAT), .B(G78GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U449 ( .A(KEYINPUT78), .B(n384), .ZN(n451) );
  XOR2_X1 U450 ( .A(n451), .B(n385), .Z(n398) );
  XOR2_X1 U451 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n389) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U454 ( .A(n390), .B(KEYINPUT23), .Z(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT24), .B(n391), .Z(n393) );
  NAND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n394), .B(KEYINPUT91), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n473) );
  XOR2_X1 U461 ( .A(n473), .B(KEYINPUT66), .Z(n399) );
  XOR2_X1 U462 ( .A(KEYINPUT28), .B(n399), .Z(n528) );
  INV_X1 U463 ( .A(n528), .ZN(n505) );
  NAND2_X1 U464 ( .A1(n521), .A2(n505), .ZN(n400) );
  NOR2_X1 U465 ( .A1(n403), .A2(n400), .ZN(n533) );
  NAND2_X1 U466 ( .A1(n401), .A2(n533), .ZN(n410) );
  NAND2_X1 U467 ( .A1(n473), .A2(n502), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n402), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U469 ( .A1(n569), .A2(n403), .ZN(n549) );
  INV_X1 U470 ( .A(n523), .ZN(n498) );
  NOR2_X1 U471 ( .A1(n502), .A2(n498), .ZN(n404) );
  NOR2_X1 U472 ( .A1(n473), .A2(n404), .ZN(n405) );
  XOR2_X1 U473 ( .A(KEYINPUT25), .B(n405), .Z(n406) );
  XNOR2_X1 U474 ( .A(KEYINPUT99), .B(n407), .ZN(n408) );
  INV_X1 U475 ( .A(n521), .ZN(n546) );
  NAND2_X1 U476 ( .A1(n408), .A2(n546), .ZN(n409) );
  NAND2_X1 U477 ( .A1(n410), .A2(n409), .ZN(n485) );
  NAND2_X1 U478 ( .A1(n462), .A2(n485), .ZN(n411) );
  NOR2_X1 U479 ( .A1(n583), .A2(n411), .ZN(n414) );
  INV_X1 U480 ( .A(KEYINPUT37), .ZN(n412) );
  XOR2_X1 U481 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n416) );
  XNOR2_X1 U482 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n430) );
  XOR2_X1 U484 ( .A(G113GAT), .B(G197GAT), .Z(n418) );
  XNOR2_X1 U485 ( .A(G22GAT), .B(G141GAT), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U487 ( .A(KEYINPUT72), .B(KEYINPUT30), .Z(n420) );
  XNOR2_X1 U488 ( .A(G169GAT), .B(G15GAT), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U490 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U491 ( .A(G43GAT), .B(n423), .Z(n425) );
  NAND2_X1 U492 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U493 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U494 ( .A(G50GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U496 ( .A(n430), .B(n429), .Z(n432) );
  XOR2_X1 U497 ( .A(n432), .B(n431), .Z(n507) );
  INV_X1 U498 ( .A(n507), .ZN(n570) );
  XOR2_X1 U499 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n450) );
  XNOR2_X1 U502 ( .A(n437), .B(KEYINPUT31), .ZN(n439) );
  XOR2_X1 U503 ( .A(KEYINPUT75), .B(KEYINPUT74), .Z(n441) );
  XNOR2_X1 U504 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n443) );
  INV_X1 U506 ( .A(KEYINPUT33), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n443), .B(n442), .ZN(n446) );
  XNOR2_X1 U508 ( .A(G176GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n574) );
  NAND2_X1 U512 ( .A1(n570), .A2(n574), .ZN(n487) );
  NOR2_X1 U513 ( .A1(n520), .A2(n487), .ZN(n453) );
  NOR2_X1 U514 ( .A1(n294), .A2(n546), .ZN(n455) );
  XNOR2_X1 U515 ( .A(KEYINPUT47), .B(KEYINPUT112), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n557), .A2(n570), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT46), .ZN(n457) );
  NAND2_X1 U518 ( .A1(n457), .A2(n462), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT111), .ZN(n459) );
  INV_X1 U520 ( .A(n564), .ZN(n482) );
  NAND2_X1 U521 ( .A1(n459), .A2(n482), .ZN(n460) );
  XNOR2_X1 U522 ( .A(n461), .B(n460), .ZN(n469) );
  XOR2_X1 U523 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n464) );
  NOR2_X1 U524 ( .A1(n462), .A2(n583), .ZN(n463) );
  XOR2_X1 U525 ( .A(n464), .B(n463), .Z(n465) );
  NAND2_X1 U526 ( .A1(n574), .A2(n465), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n570), .A2(n466), .ZN(n467) );
  XOR2_X1 U528 ( .A(KEYINPUT113), .B(n467), .Z(n468) );
  NOR2_X1 U529 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT48), .ZN(n547) );
  NOR2_X1 U531 ( .A1(n498), .A2(n547), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n471), .B(KEYINPUT54), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n546), .ZN(n568) );
  NOR2_X1 U534 ( .A1(n473), .A2(n568), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n565), .A2(n570), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n476) );
  XNOR2_X1 U538 ( .A(n476), .B(G169GAT), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(G1348GAT) );
  NAND2_X1 U540 ( .A1(n565), .A2(n557), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n484) );
  NAND2_X1 U543 ( .A1(n579), .A2(n482), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n508) );
  NOR2_X1 U546 ( .A1(n487), .A2(n508), .ZN(n496) );
  NAND2_X1 U547 ( .A1(n521), .A2(n496), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT100), .ZN(n489) );
  XOR2_X1 U549 ( .A(n489), .B(KEYINPUT101), .Z(n491) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1324GAT) );
  NAND2_X1 U552 ( .A1(n496), .A2(n523), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n492), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U555 ( .A1(n496), .A2(n532), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U558 ( .A1(n496), .A2(n528), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U560 ( .A1(n294), .A2(n498), .ZN(n499) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(n504) );
  NOR2_X1 U565 ( .A1(n502), .A2(n294), .ZN(n503) );
  XOR2_X1 U566 ( .A(n504), .B(n503), .Z(G1330GAT) );
  NOR2_X1 U567 ( .A1(n294), .A2(n505), .ZN(n506) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n506), .Z(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  NAND2_X1 U570 ( .A1(n507), .A2(n557), .ZN(n519) );
  NOR2_X1 U571 ( .A1(n519), .A2(n508), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n515), .A2(n521), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n515), .A2(n523), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT106), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U578 ( .A1(n515), .A2(n532), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n528), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n529), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n522), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n525) );
  NAND2_X1 U588 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n532), .A2(n529), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n536) );
  NAND2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U598 ( .A1(n547), .A2(n534), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n541), .A2(n570), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U602 ( .A1(n541), .A2(n557), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n541), .A2(n579), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n564), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT115), .Z(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n552) );
  NOR2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT117), .B(n550), .ZN(n561) );
  NAND2_X1 U616 ( .A1(n561), .A2(n570), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT52), .B(n556), .Z(n559) );
  NAND2_X1 U623 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n579), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n564), .A2(n561), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n579), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n580), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n580), .ZN(n582) );
  NOR2_X1 U640 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

