//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G107), .A2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(G50), .B2(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G116), .ZN(new_n222));
  INV_X1    g0022(.A(G270), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(G20), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(G58), .A2(G68), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n210), .B(new_n229), .C1(new_n232), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n223), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT66), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  OR2_X1    g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G222), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n256), .B(new_n258), .C1(new_n259), .C2(new_n257), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n225), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n260), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT68), .B1(new_n262), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g0072(.A(G226), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n269), .B(G274), .C1(G41), .C2(G45), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT67), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n268), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n268), .A2(new_n273), .A3(KEYINPUT69), .A4(new_n275), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n269), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G50), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n230), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n231), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n295));
  INV_X1    g0095(.A(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n231), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G150), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n295), .A2(new_n231), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n291), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n285), .A2(new_n286), .ZN(new_n301));
  INV_X1    g0101(.A(new_n291), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n231), .A2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n301), .A2(new_n302), .A3(G50), .A4(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n289), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n278), .A2(new_n279), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n282), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT71), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n280), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n307), .A2(KEYINPUT71), .A3(G190), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n306), .B(KEYINPUT9), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n278), .A2(G200), .A3(new_n279), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT71), .B1(new_n307), .B2(G190), .ZN(new_n323));
  AOI211_X1 g0123(.A(new_n312), .B(new_n313), .C1(new_n278), .C2(new_n279), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(KEYINPUT10), .B1(new_n325), .B2(new_n320), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n311), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n262), .A2(G232), .A3(new_n270), .ZN(new_n328));
  INV_X1    g0128(.A(G226), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n254), .A2(new_n255), .B1(new_n329), .B2(G1698), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n259), .A2(new_n257), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n330), .A2(new_n331), .B1(G33), .B2(G87), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n275), .B(new_n328), .C1(new_n332), .C2(new_n262), .ZN(new_n333));
  INV_X1    g0133(.A(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n331), .B1(G226), .B2(new_n257), .C1(new_n264), .C2(new_n265), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G33), .A2(G87), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n263), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n339), .A2(new_n313), .A3(new_n275), .A4(new_n328), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n291), .B1(new_n285), .B2(new_n286), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n292), .B1(new_n341), .B2(new_n304), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n301), .A2(new_n292), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT75), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT75), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n303), .B(new_n291), .C1(new_n285), .C2(new_n286), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(new_n343), .C1(new_n347), .C2(new_n292), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n335), .A2(new_n340), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n254), .A2(new_n231), .A3(new_n255), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT74), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n231), .A4(new_n255), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n354), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(G68), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n216), .A2(new_n212), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n233), .ZN(new_n360));
  INV_X1    g0160(.A(new_n297), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G159), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n212), .B1(new_n352), .B2(new_n354), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n366), .B1(new_n367), .B2(new_n363), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n365), .A2(new_n291), .A3(new_n368), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n349), .A2(KEYINPUT77), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT77), .B1(new_n349), .B2(new_n369), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT17), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n345), .A2(new_n348), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n335), .A2(new_n340), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(KEYINPUT17), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n333), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n281), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n333), .A2(new_n308), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT76), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(G179), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n382), .B(new_n383), .C1(new_n281), .C2(new_n378), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n369), .A2(new_n373), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT18), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(KEYINPUT18), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n372), .A2(new_n377), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n327), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n257), .A2(G232), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n256), .B(new_n393), .C1(new_n213), .C2(new_n257), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n394), .B(new_n263), .C1(G107), .C2(new_n256), .ZN(new_n395));
  OAI21_X1  g0195(.A(G244), .B1(new_n271), .B2(new_n272), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(new_n275), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n281), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n347), .A2(G77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n287), .A2(new_n225), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n292), .A2(new_n297), .B1(new_n231), .B2(new_n225), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT15), .B(G87), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n293), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n291), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n398), .B(new_n405), .C1(G179), .C2(new_n397), .ZN(new_n406));
  OAI21_X1  g0206(.A(G238), .B1(new_n271), .B2(new_n272), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n329), .A2(new_n257), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n217), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n409), .C1(new_n264), .C2(new_n265), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G97), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n263), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n413), .A3(new_n275), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT72), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT13), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n407), .A2(new_n413), .A3(new_n417), .A4(new_n275), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(G169), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT14), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n415), .A2(new_n418), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G179), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n419), .A2(new_n425), .A3(G169), .A4(new_n420), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n287), .A2(new_n212), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT12), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n347), .A2(G68), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n293), .A2(new_n225), .B1(new_n231), .B2(G68), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n297), .A2(new_n288), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n291), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g0233(.A(new_n433), .B(KEYINPUT11), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n419), .A2(G200), .A3(new_n420), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(KEYINPUT73), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n435), .B1(new_n423), .B2(G190), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(KEYINPUT73), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n397), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n405), .B1(new_n442), .B2(G190), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n397), .A2(G200), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n436), .A2(new_n441), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n391), .A2(new_n392), .A3(new_n406), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n327), .A2(new_n390), .A3(new_n406), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT78), .B1(new_n449), .B2(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n269), .A2(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n341), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n301), .A2(G97), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT7), .B1(new_n266), .B2(new_n231), .ZN(new_n459));
  OAI21_X1  g0259(.A(G107), .B1(new_n459), .B2(new_n356), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT6), .ZN(new_n461));
  AND2_X1   g0261(.A1(G97), .A2(G107), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n202), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(KEYINPUT6), .A3(G97), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(G20), .B1(G77), .B2(new_n361), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT79), .B1(new_n468), .B2(new_n291), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT79), .ZN(new_n470));
  AOI211_X1 g0270(.A(new_n470), .B(new_n302), .C1(new_n460), .C2(new_n467), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n456), .B(new_n458), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT4), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n474), .B(G244), .C1(new_n265), .C2(new_n264), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n226), .B1(new_n254), .B2(new_n255), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(G250), .B1(new_n264), .B2(new_n265), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n257), .B1(new_n479), .B2(KEYINPUT4), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n263), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT80), .B1(new_n482), .B2(G41), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n269), .A2(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n263), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n269), .B(G45), .C1(new_n485), .C2(KEYINPUT5), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n483), .B2(new_n486), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n491), .A2(G257), .B1(G274), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(G169), .B1(new_n481), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n481), .A2(new_n494), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n308), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n472), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n464), .A2(KEYINPUT6), .A3(G97), .ZN(new_n499));
  XNOR2_X1  g0299(.A(G97), .B(G107), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n461), .ZN(new_n501));
  OAI22_X1  g0301(.A1(new_n501), .A2(new_n231), .B1(new_n225), .B2(new_n297), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n464), .B1(new_n352), .B2(new_n354), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n291), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n470), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n468), .A2(KEYINPUT79), .A3(new_n291), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n457), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n481), .A2(new_n494), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n334), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n481), .A2(new_n313), .A3(new_n494), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n507), .A2(new_n511), .A3(new_n456), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT19), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n293), .B2(new_n454), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n231), .B1(new_n411), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(G87), .B2(new_n203), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n231), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n519));
  OAI211_X1 g0319(.A(KEYINPUT82), .B(new_n513), .C1(new_n293), .C2(new_n454), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n291), .ZN(new_n522));
  INV_X1    g0322(.A(new_n402), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n341), .A2(new_n523), .A3(new_n452), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n287), .A2(new_n402), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(G45), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n221), .B1(new_n527), .B2(G1), .ZN(new_n528));
  INV_X1    g0328(.A(G274), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n269), .A2(new_n529), .A3(G45), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n262), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT81), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT81), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n262), .A2(new_n528), .A3(new_n530), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n213), .A2(new_n257), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n226), .A2(G1698), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n535), .B(new_n536), .C1(new_n264), .C2(new_n265), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n532), .A2(new_n534), .B1(new_n539), .B2(new_n263), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n308), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n532), .A2(new_n534), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n263), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n281), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n526), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(G200), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n341), .A2(G87), .A3(new_n452), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n521), .A2(new_n291), .B1(new_n287), .B2(new_n402), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n543), .A3(G190), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n491), .A2(G264), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n221), .A2(new_n257), .ZN(new_n555));
  INV_X1    g0355(.A(G257), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G1698), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n555), .B(new_n557), .C1(new_n264), .C2(new_n265), .ZN(new_n558));
  INV_X1    g0358(.A(G294), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n296), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n263), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n493), .A2(G274), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n554), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n334), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(G190), .B2(new_n563), .ZN(new_n565));
  XNOR2_X1  g0365(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n256), .A2(new_n566), .A3(new_n231), .A4(G87), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n231), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(KEYINPUT22), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n231), .A2(G33), .A3(G116), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n231), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n464), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n567), .A2(new_n571), .A3(new_n572), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT84), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n568), .A2(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(KEYINPUT84), .A3(new_n567), .A4(new_n572), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(KEYINPUT24), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n577), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n291), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n287), .A2(new_n464), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n453), .A2(new_n464), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n287), .B2(new_n464), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n565), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n498), .A2(new_n512), .A3(new_n553), .A4(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n301), .A2(new_n302), .A3(G116), .A4(new_n452), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n285), .A2(new_n222), .A3(new_n286), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n290), .A2(new_n230), .B1(G20), .B2(new_n222), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n476), .B(new_n231), .C1(G33), .C2(new_n454), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(KEYINPUT20), .A3(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n595), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n487), .A2(new_n490), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G270), .A3(new_n262), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G264), .A2(G1698), .ZN(new_n604));
  OAI221_X1 g0404(.A(new_n604), .B1(new_n556), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n605));
  INV_X1    g0405(.A(G303), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n266), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n607), .A3(new_n263), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n603), .A2(new_n608), .A3(new_n562), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n601), .A2(G169), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(G200), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n491), .A2(G270), .B1(G274), .B2(new_n493), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(G190), .A3(new_n608), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n596), .B1(new_n600), .B2(new_n599), .ZN(new_n616));
  INV_X1    g0416(.A(new_n595), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n613), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n601), .A2(G179), .A3(new_n608), .A4(new_n614), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n601), .A2(KEYINPUT21), .A3(new_n609), .A4(G169), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n612), .A2(new_n619), .A3(new_n620), .A4(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n585), .A2(new_n592), .ZN(new_n624));
  AOI22_X1  g0424(.A1(G264), .A2(new_n491), .B1(new_n560), .B2(new_n263), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT86), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(G179), .A4(new_n562), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT86), .B1(new_n563), .B2(G169), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n563), .A2(new_n308), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n594), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n451), .A2(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n436), .A2(new_n406), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n372), .A2(new_n377), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n441), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n382), .B1(new_n281), .B2(new_n378), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n385), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT18), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n317), .B1(new_n316), .B2(new_n321), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n325), .A2(KEYINPUT10), .A3(new_n320), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n311), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n451), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n546), .B(KEYINPUT87), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n612), .A2(new_n620), .A3(new_n621), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n624), .B2(new_n630), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n594), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n481), .A2(new_n308), .A3(new_n494), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n496), .B2(G169), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n456), .B2(new_n507), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT26), .B1(new_n655), .B2(new_n553), .ZN(new_n656));
  AOI211_X1 g0456(.A(new_n455), .B(new_n457), .C1(new_n505), .C2(new_n506), .ZN(new_n657));
  XNOR2_X1  g0457(.A(KEYINPUT88), .B(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR4_X1   g0459(.A1(new_n657), .A2(new_n552), .A3(new_n654), .A4(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n647), .B1(new_n648), .B2(new_n662), .ZN(G369));
  AND3_X1   g0463(.A1(new_n565), .A2(new_n585), .A3(new_n592), .ZN(new_n664));
  INV_X1    g0464(.A(G13), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G20), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OR3_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .A3(G1), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT27), .B1(new_n667), .B2(G1), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n585), .B2(new_n592), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n631), .B1(new_n664), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n624), .A2(new_n630), .A3(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT89), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n650), .A2(new_n673), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n673), .A2(new_n618), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n650), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n622), .B2(new_n685), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(G330), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n683), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n235), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n673), .B1(new_n652), .B2(new_n661), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n655), .A2(new_n553), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n658), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(KEYINPUT26), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n673), .B1(new_n701), .B2(new_n652), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n625), .A2(G179), .A3(new_n608), .A4(new_n614), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n481), .A2(new_n494), .A3(new_n540), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT91), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n707), .A2(new_n708), .A3(new_n706), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n609), .A2(new_n544), .A3(new_n308), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT90), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT90), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n609), .A2(new_n544), .A3(new_n714), .A4(new_n308), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n508), .A3(new_n563), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT91), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n717), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n710), .A2(new_n711), .A3(new_n716), .A4(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(KEYINPUT31), .B1(new_n719), .B2(new_n672), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n633), .B2(new_n673), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n711), .A2(new_n716), .A3(new_n709), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n705), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n696), .B1(new_n727), .B2(G1), .ZN(G364));
  AOI21_X1  g0528(.A(new_n230), .B1(G20), .B2(new_n281), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n231), .A2(new_n308), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(G190), .A3(new_n334), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n313), .A2(new_n334), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n231), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n732), .A2(G58), .B1(new_n736), .B2(G87), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n334), .A2(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n737), .B1(new_n464), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G159), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT32), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n231), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n454), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n730), .A2(new_n738), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n256), .B1(new_n749), .B2(new_n212), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n745), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n730), .A2(new_n733), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT92), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n751), .B1(new_n288), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n730), .A2(new_n741), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n740), .B(new_n758), .C1(G77), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI22_X1  g0563(.A1(new_n762), .A2(new_n731), .B1(new_n763), .B2(new_n749), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n735), .B(KEYINPUT93), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n747), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G303), .B1(G294), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n757), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G326), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n760), .A2(G311), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n256), .B1(new_n743), .B2(G329), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n739), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n765), .B(new_n774), .C1(G283), .C2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n729), .B1(new_n761), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n690), .A2(new_n266), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G355), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n690), .A2(new_n256), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n235), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n252), .A2(G45), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n779), .B1(G116), .B2(new_n207), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n729), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n269), .B1(new_n666), .B2(G45), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n691), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n786), .B(KEYINPUT95), .Z(new_n792));
  OAI211_X1 g0592(.A(new_n686), .B(new_n792), .C1(new_n622), .C2(new_n685), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n777), .A2(new_n788), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n791), .B1(new_n687), .B2(G330), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G330), .B2(new_n687), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n794), .A2(new_n796), .ZN(G396));
  INV_X1    g0597(.A(G137), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n757), .A2(new_n798), .B1(new_n298), .B2(new_n749), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT96), .Z(new_n800));
  INV_X1    g0600(.A(G143), .ZN(new_n801));
  INV_X1    g0601(.A(G159), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n731), .A2(new_n801), .B1(new_n759), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT34), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n805), .A2(new_n806), .B1(G68), .B2(new_n775), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n216), .B2(new_n747), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n766), .A2(new_n288), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n742), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n256), .B1(new_n805), .B2(new_n806), .ZN(new_n812));
  NOR4_X1   g0612(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G283), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n766), .A2(new_n464), .B1(new_n814), .B2(new_n749), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n256), .B(new_n815), .C1(G294), .C2(new_n732), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n606), .B2(new_n757), .C1(new_n817), .C2(new_n742), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n739), .A2(new_n220), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n759), .A2(new_n222), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n818), .A2(new_n748), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n729), .B1(new_n813), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n822), .A2(new_n791), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n729), .A2(new_n784), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n405), .A2(new_n672), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n445), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n406), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n406), .A2(new_n672), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n823), .B1(G77), .B2(new_n825), .C1(new_n785), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n697), .A2(new_n831), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n832), .B(new_n673), .C1(new_n652), .C2(new_n661), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(new_n725), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(new_n791), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT40), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n343), .B1(new_n347), .B2(new_n292), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n365), .A2(new_n291), .ZN(new_n842));
  AOI21_X1  g0642(.A(KEYINPUT16), .B1(new_n358), .B2(new_n364), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n638), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(KEYINPUT100), .C1(new_n370), .C2(new_n371), .ZN(new_n846));
  INV_X1    g0646(.A(new_n670), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT77), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n375), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n349), .A2(KEYINPUT77), .A3(new_n369), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT100), .B1(new_n853), .B2(new_n845), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n385), .A2(new_n847), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n386), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n388), .A2(new_n389), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n848), .B1(new_n636), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(KEYINPUT38), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n856), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n376), .B1(new_n853), .B2(KEYINPUT17), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n869), .B1(new_n870), .B2(new_n640), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n639), .A2(new_n856), .A3(new_n375), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n857), .A2(new_n859), .B1(new_n872), .B2(new_n858), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n840), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n435), .A2(new_n672), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n436), .A2(new_n441), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n427), .A2(new_n435), .A3(new_n672), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n831), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n498), .A2(new_n512), .A3(new_n553), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n622), .B1(new_n624), .B2(new_n630), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n882), .A2(new_n593), .A3(new_n883), .A4(new_n673), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n719), .A2(new_n672), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT31), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT104), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n721), .A2(KEYINPUT104), .A3(new_n888), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n881), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n876), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT104), .B1(new_n721), .B2(new_n888), .ZN(new_n895));
  AND4_X1   g0695(.A1(KEYINPUT104), .A2(new_n884), .A3(new_n887), .A4(new_n888), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n880), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT38), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n845), .B1(new_n370), .B2(new_n371), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT100), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n846), .A3(new_n848), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n860), .B1(new_n902), .B2(KEYINPUT37), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n898), .B1(new_n903), .B2(new_n864), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n897), .B1(new_n866), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(G330), .B(new_n894), .C1(new_n905), .C2(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n891), .A2(new_n892), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n451), .A2(G330), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n866), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n893), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n910), .A2(new_n840), .B1(new_n893), .B2(new_n876), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n448), .A2(new_n450), .B1(new_n891), .B2(new_n892), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n906), .A2(new_n908), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n913), .B(KEYINPUT103), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n451), .A2(new_n704), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n647), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n914), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n640), .A2(new_n670), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n835), .A2(new_n830), .B1(new_n878), .B2(new_n879), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n904), .A2(new_n866), .A3(KEYINPUT39), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n864), .B1(new_n855), .B2(new_n861), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n874), .B1(new_n923), .B2(KEYINPUT38), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n922), .B1(KEYINPUT39), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n427), .A2(new_n435), .A3(new_n673), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT101), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n919), .B(new_n921), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n918), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n269), .B2(new_n666), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n235), .A2(new_n225), .A3(new_n359), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT99), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(G50), .B2(new_n212), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(G1), .A3(new_n665), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n501), .B(KEYINPUT97), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n222), .B1(new_n935), .B2(KEYINPUT35), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n936), .B(new_n232), .C1(KEYINPUT35), .C2(new_n935), .ZN(new_n937));
  XOR2_X1   g0737(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n938));
  XNOR2_X1  g0738(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n930), .A2(new_n934), .A3(new_n939), .ZN(G367));
  OAI211_X1 g0740(.A(new_n498), .B(new_n512), .C1(new_n657), .C2(new_n673), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n681), .A2(KEYINPUT42), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n676), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n655), .A2(new_n673), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT42), .B1(new_n681), .B2(new_n941), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n549), .A2(new_n548), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n672), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n649), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n553), .A2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n946), .A2(KEYINPUT43), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n655), .A2(new_n672), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n941), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n688), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n946), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n952), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n956), .B1(new_n952), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n691), .B(new_n964), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n681), .A2(new_n676), .A3(new_n954), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT44), .B1(new_n683), .B2(new_n954), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT44), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n682), .A2(new_n971), .A3(new_n955), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n688), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n684), .A2(new_n680), .B1(G330), .B2(new_n687), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT106), .B1(new_n684), .B2(new_n680), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(new_n726), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n969), .A2(new_n970), .A3(new_n688), .A4(new_n972), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n966), .B1(new_n981), .B2(new_n727), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n963), .B1(new_n982), .B2(new_n790), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n814), .A2(new_n759), .B1(new_n749), .B2(new_n559), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT46), .B1(new_n766), .B2(new_n222), .ZN(new_n985));
  OR3_X1    g0785(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n222), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n256), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n987), .B1(new_n464), .B2(new_n747), .C1(new_n988), .C2(new_n742), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n984), .B(new_n989), .C1(G311), .C2(new_n770), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n454), .B2(new_n739), .C1(new_n606), .C2(new_n731), .ZN(new_n991));
  INV_X1    g0791(.A(new_n749), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G159), .A2(new_n992), .B1(new_n760), .B2(G50), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n216), .B2(new_n735), .C1(new_n798), .C2(new_n742), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n739), .A2(new_n225), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n994), .A2(new_n266), .A3(new_n995), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n747), .A2(new_n212), .B1(new_n731), .B2(new_n298), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT107), .Z(new_n998));
  OAI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(new_n801), .C2(new_n757), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n991), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n729), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n949), .A2(new_n792), .A3(new_n950), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n780), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n787), .B1(new_n207), .B2(new_n402), .C1(new_n244), .C2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n791), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT108), .Z(new_n1007));
  NAND2_X1  g0807(.A1(new_n983), .A2(new_n1007), .ZN(G387));
  AOI21_X1  g0808(.A(new_n692), .B1(new_n978), .B2(new_n726), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n726), .B2(new_n978), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n684), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n792), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G77), .A2(new_n736), .B1(new_n743), .B2(G150), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n256), .B(new_n1013), .C1(new_n757), .C2(new_n802), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n747), .A2(new_n402), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n731), .A2(new_n288), .B1(new_n749), .B2(new_n292), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n759), .A2(new_n212), .B1(new_n739), .B2(new_n454), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT110), .Z(new_n1019));
  AOI22_X1  g0819(.A1(new_n732), .A2(G317), .B1(new_n760), .B2(G303), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n757), .A2(new_n762), .B1(new_n817), .B2(new_n749), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n814), .B2(new_n747), .C1(new_n559), .C2(new_n735), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT49), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n775), .A2(G116), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n743), .A2(G326), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1028), .A2(new_n266), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n729), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1004), .B1(new_n241), .B2(G45), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n693), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n778), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n292), .A2(G50), .ZN(new_n1038));
  XOR2_X1   g0838(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n693), .B(new_n527), .C1(new_n212), .C2(new_n225), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1037), .A2(new_n1042), .B1(G107), .B2(new_n207), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n787), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1034), .A2(new_n791), .A3(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1010), .B1(new_n789), .B2(new_n978), .C1(new_n1012), .C2(new_n1045), .ZN(G393));
  INV_X1    g0846(.A(KEYINPUT112), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n975), .A2(new_n1047), .A3(new_n980), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n980), .A2(new_n1047), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n691), .B(new_n981), .C1(new_n1050), .C2(new_n979), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n780), .A2(new_n248), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n787), .C1(new_n454), .C2(new_n207), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n759), .A2(new_n292), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n757), .A2(new_n298), .B1(new_n802), .B2(new_n731), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT51), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n747), .A2(new_n225), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n819), .B(new_n1057), .C1(G50), .C2(new_n992), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n256), .A3(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1054), .B(new_n1059), .C1(G143), .C2(new_n743), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n736), .A2(G68), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n736), .A2(G283), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n757), .A2(new_n988), .B1(new_n817), .B2(new_n731), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n992), .A2(G303), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n759), .A2(new_n559), .B1(new_n739), .B2(new_n464), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G116), .B2(new_n768), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1064), .A2(new_n266), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G322), .B2(new_n743), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1060), .A2(new_n1061), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT113), .Z(new_n1071));
  INV_X1    g0871(.A(new_n729), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n791), .B(new_n1053), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n786), .B2(new_n955), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1050), .B2(new_n790), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1051), .A2(new_n1075), .ZN(G390));
  NAND2_X1  g0876(.A1(new_n824), .A2(new_n292), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n757), .A2(new_n1078), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n256), .B1(new_n739), .B2(new_n288), .C1(new_n798), .C2(new_n749), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT54), .B(G143), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n760), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n732), .A2(G132), .B1(new_n743), .B2(G125), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n735), .A2(new_n298), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT53), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1079), .B(new_n1086), .C1(G159), .C2(new_n768), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n770), .A2(G283), .B1(G107), .B2(new_n992), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n454), .B2(new_n759), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT117), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n766), .A2(new_n220), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n266), .B1(new_n742), .B2(new_n559), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n731), .A2(new_n222), .B1(new_n739), .B2(new_n212), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n1091), .A2(new_n1057), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1087), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT118), .Z(new_n1096));
  OAI211_X1 g0896(.A(new_n791), .B(new_n1077), .C1(new_n1096), .C2(new_n1072), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n925), .B2(new_n784), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT119), .Z(new_n1099));
  INV_X1    g0899(.A(KEYINPUT114), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n927), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n920), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n835), .A2(new_n830), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n878), .A2(new_n879), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(KEYINPUT114), .A3(new_n927), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n904), .A2(new_n866), .A3(KEYINPUT39), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT39), .B1(new_n866), .B2(new_n875), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1102), .B(new_n1106), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n673), .B(new_n828), .C1(new_n701), .C2(new_n652), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1110), .A2(new_n830), .B1(new_n878), .B2(new_n879), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n924), .A2(new_n1111), .A3(new_n1101), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n725), .A2(new_n881), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1109), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT114), .B1(new_n1105), .B2(new_n927), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n920), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1112), .B1(new_n1119), .B2(new_n925), .ZN(new_n1120));
  INV_X1    g0920(.A(G330), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n891), .B2(new_n892), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n880), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1099), .B1(new_n789), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n912), .A2(KEYINPUT115), .A3(G330), .ZN(new_n1126));
  AOI21_X1  g0926(.A(KEYINPUT115), .B1(new_n912), .B2(G330), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n917), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1104), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n832), .B1(new_n1122), .B2(KEYINPUT116), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n907), .A2(KEYINPUT116), .A3(G330), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1115), .A2(new_n830), .A3(new_n1110), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1130), .B1(new_n725), .B2(new_n831), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1103), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1124), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1114), .B(new_n1112), .C1(new_n1119), .C2(new_n925), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1123), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1133), .A2(new_n1134), .B1(new_n1103), .B2(new_n1137), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(new_n1128), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n692), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1125), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(G378));
  OAI21_X1  g0949(.A(new_n791), .B1(G50), .B2(new_n825), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n288), .B1(new_n264), .B2(G41), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n775), .A2(G58), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n464), .B2(new_n731), .C1(new_n757), .C2(new_n222), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n485), .B(new_n266), .C1(new_n735), .C2(new_n225), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT120), .Z(new_n1155));
  AOI22_X1  g0955(.A1(new_n768), .A2(G68), .B1(new_n760), .B2(new_n523), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n814), .C2(new_n742), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G97), .C2(new_n992), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT58), .Z(new_n1159));
  AOI22_X1  g0959(.A1(new_n770), .A2(G125), .B1(G150), .B2(new_n768), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT121), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n992), .A2(G132), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n736), .A2(new_n1081), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n732), .A2(G128), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G137), .B2(new_n760), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  OR2_X1    g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n775), .A2(G159), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G33), .B1(new_n743), .B2(G124), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1168), .A2(new_n485), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1151), .B(new_n1159), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1150), .B1(new_n1173), .B2(new_n729), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n327), .B(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n306), .A2(new_n847), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1174), .B1(new_n1178), .B2(new_n785), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n906), .A2(new_n1178), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n910), .A2(new_n840), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1178), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(G330), .A4(new_n894), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1181), .A2(new_n928), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n928), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT122), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n928), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n911), .B2(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT122), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1187), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1180), .B1(new_n1194), .B2(new_n790), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1129), .B1(new_n1124), .B2(new_n1145), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1181), .A2(new_n928), .A3(new_n1184), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1196), .A3(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n691), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1197), .B2(new_n1201), .ZN(G375));
  OAI21_X1  g1002(.A(new_n791), .B1(G68), .B2(new_n825), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1130), .A2(new_n784), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT123), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n256), .B1(new_n742), .B2(new_n1078), .C1(new_n747), .C2(new_n288), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1152), .B1(new_n766), .B2(new_n802), .C1(new_n757), .C2(new_n810), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n992), .C2(new_n1081), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n798), .B2(new_n731), .C1(new_n298), .C2(new_n759), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n766), .A2(new_n454), .B1(new_n606), .B2(new_n742), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT124), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n256), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n732), .A2(G283), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n770), .A2(G294), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n995), .B(new_n1015), .C1(G107), .C2(new_n760), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n749), .A2(new_n222), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1209), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n1203), .B(new_n1205), .C1(new_n729), .C2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n1139), .B2(new_n790), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1140), .A2(new_n965), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1220), .B1(new_n1221), .B2(new_n1222), .ZN(G381));
  NAND2_X1  g1023(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT122), .B1(new_n1224), .B2(new_n1188), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1199), .B2(KEYINPUT122), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1179), .B1(new_n1226), .B2(new_n789), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1128), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1201), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1148), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G381), .A2(G384), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n983), .A2(new_n1051), .A3(new_n1007), .A4(new_n1075), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1236), .A2(G396), .A3(G393), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(G407));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(G343), .C2(new_n1233), .ZN(G409));
  NAND2_X1  g1039(.A1(new_n671), .A2(G213), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1192), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n965), .B(new_n1196), .C1(new_n1241), .C2(new_n1225), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1199), .A2(new_n790), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1148), .A2(new_n1242), .A3(new_n1179), .A4(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1240), .B(new_n1244), .C1(new_n1232), .C2(new_n1148), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1222), .A2(KEYINPUT60), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1145), .A2(new_n1128), .A3(KEYINPUT60), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1140), .A2(new_n691), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1220), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n838), .A3(new_n833), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G384), .B(new_n1220), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1240), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G2897), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1250), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1245), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1229), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n691), .B(new_n1200), .C1(new_n1258), .C2(KEYINPUT57), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1148), .B1(new_n1259), .B2(new_n1195), .ZN(new_n1260));
  AND4_X1   g1060(.A1(new_n1148), .A2(new_n1242), .A3(new_n1179), .A4(new_n1243), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1262));
  NOR4_X1   g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1252), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1257), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G375), .A2(G378), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1262), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1240), .A4(new_n1244), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1266), .B1(new_n1269), .B2(KEYINPUT62), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  XOR2_X1   g1071(.A(G393), .B(G396), .Z(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1236), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1274), .B2(new_n1236), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1273), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1277), .A2(new_n1273), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1263), .A2(KEYINPUT63), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT63), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1269), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1257), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1245), .A2(new_n1256), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1271), .A2(new_n1281), .B1(new_n1286), .B2(new_n1290), .ZN(G405));
  XNOR2_X1  g1091(.A(new_n1262), .B(KEYINPUT127), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1234), .B2(new_n1260), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT127), .ZN(new_n1294));
  XNOR2_X1  g1094(.A(new_n1262), .B(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1295), .A2(new_n1233), .A3(new_n1267), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1280), .A2(new_n1293), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1280), .B1(new_n1296), .B2(new_n1293), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


