//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n202), .A2(G1gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G43gat), .A2(G50gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT15), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT14), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G29gat), .B2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT88), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT88), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n213), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n216), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n213), .A2(new_n219), .A3(new_n217), .A4(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT15), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(KEYINPUT89), .A2(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT89), .A2(G50gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G43gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n224), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n218), .A2(G29gat), .A3(G36gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT14), .B1(new_n214), .B2(new_n215), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n221), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n223), .A3(new_n225), .ZN(new_n240));
  INV_X1    g039(.A(new_n213), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT89), .B(G50gat), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n227), .B(new_n210), .C1(new_n243), .C2(G43gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n220), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n213), .A3(new_n245), .A4(new_n225), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT90), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n209), .B1(new_n236), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G229gat), .A2(G233gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n235), .B1(new_n224), .B2(new_n234), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(KEYINPUT90), .A3(new_n246), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT17), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n207), .B(G8gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n242), .A2(KEYINPUT17), .A3(new_n246), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n248), .B(new_n249), .C1(new_n252), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(KEYINPUT18), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n249), .B(KEYINPUT13), .Z(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n253), .A2(new_n251), .A3(new_n250), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n263), .B1(new_n248), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(G197gat), .ZN(new_n269));
  XOR2_X1   g068(.A(KEYINPUT11), .B(G169gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT12), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n259), .A2(new_n272), .A3(new_n261), .A4(new_n266), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G64gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G57gat), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n278), .A2(KEYINPUT93), .ZN(new_n279));
  NOR2_X1   g078(.A1(G71gat), .A2(G78gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT9), .ZN(new_n281));
  NAND2_X1  g080(.A1(G71gat), .A2(G78gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G57gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G64gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n278), .A3(KEYINPUT93), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n279), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n282), .B1(new_n280), .B2(KEYINPUT92), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n282), .A2(KEYINPUT92), .ZN(new_n289));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n288), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT21), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G231gat), .A2(G233gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(G127gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n287), .A2(new_n292), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT95), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT95), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n287), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(KEYINPUT21), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n253), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n302), .ZN(new_n304));
  XNOR2_X1  g103(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT94), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n306), .B(G155gat), .ZN(new_n307));
  XOR2_X1   g106(.A(G183gat), .B(G211gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n303), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n303), .B2(new_n304), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n250), .A2(new_n251), .ZN(new_n314));
  XNOR2_X1  g113(.A(G99gat), .B(G106gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT8), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(G99gat), .B2(G106gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(KEYINPUT96), .A2(G85gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G92gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G85gat), .A2(G92gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT7), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n320), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(new_n322), .A3(new_n318), .ZN(new_n328));
  INV_X1    g127(.A(new_n317), .ZN(new_n329));
  AND4_X1   g128(.A1(new_n315), .A2(new_n325), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT41), .ZN(new_n333));
  NAND2_X1  g132(.A1(G232gat), .A2(G233gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n254), .B1(new_n330), .B2(new_n326), .ZN(new_n335));
  OAI221_X1 g134(.A(new_n332), .B1(new_n333), .B2(new_n334), .C1(new_n252), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G190gat), .B(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT97), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G134gat), .B(G162gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n336), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n336), .B2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n338), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n334), .A2(new_n333), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OR3_X1    g147(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n343), .B2(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n313), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G230gat), .A2(G233gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n297), .B1(new_n326), .B2(new_n330), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n356));
  INV_X1    g155(.A(new_n315), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n325), .A2(new_n328), .A3(new_n315), .A4(new_n329), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n292), .A3(new_n287), .A4(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n331), .A2(KEYINPUT10), .A3(new_n298), .A4(new_n300), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n354), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n353), .B1(new_n355), .B2(new_n360), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(G120gat), .B(G148gat), .Z(new_n367));
  XNOR2_X1  g166(.A(G176gat), .B(G204gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n366), .B(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n352), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT70), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT70), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G211gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT22), .B1(new_n380), .B2(G218gat), .ZN(new_n381));
  XOR2_X1   g180(.A(G197gat), .B(G204gat), .Z(new_n382));
  OAI21_X1  g181(.A(new_n375), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT70), .B(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n374), .A3(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n373), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n391));
  AND2_X1   g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G141gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT75), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT75), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G141gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(G148gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n395), .A2(G148gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT76), .B(G162gat), .ZN(new_n403));
  INV_X1    g202(.A(G155gat), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT2), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT74), .B(KEYINPUT2), .ZN(new_n407));
  INV_X1    g206(.A(G148gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n408), .A2(G141gat), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n394), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n391), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n406), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT71), .B(KEYINPUT29), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n390), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(G228gat), .A3(G233gat), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n414), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n374), .B1(new_n387), .B2(new_n388), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n421), .B2(KEYINPUT82), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n383), .A2(new_n423), .A3(new_n389), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n402), .A2(new_n405), .B1(new_n410), .B2(new_n394), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n417), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n428));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n419), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n372), .B1(new_n432), .B2(G22gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(KEYINPUT31), .B(G50gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n427), .A2(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n442), .B2(new_n419), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n413), .A2(new_n418), .ZN(new_n444));
  AOI211_X1 g243(.A(G22gat), .B(new_n444), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  OAI22_X1  g244(.A1(new_n433), .A2(new_n437), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n432), .A2(G22gat), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n442), .A2(new_n438), .A3(new_n419), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n372), .A4(new_n436), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT23), .ZN(new_n452));
  INV_X1    g251(.A(G169gat), .ZN(new_n453));
  INV_X1    g252(.A(G176gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT23), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND3_X1   g257(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n460));
  OAI21_X1  g259(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT25), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT25), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n465), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT26), .ZN(new_n468));
  NAND2_X1  g267(.A1(G183gat), .A2(G190gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT26), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(G169gat), .B2(G176gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n451), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n468), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n470), .A3(new_n451), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n476), .A2(KEYINPUT65), .A3(new_n469), .A4(new_n468), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n479));
  INV_X1    g278(.A(G183gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT27), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT27), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G183gat), .ZN(new_n483));
  INV_X1    g282(.A(G190gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(KEYINPUT64), .A2(KEYINPUT28), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G183gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(new_n484), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n479), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI22_X1  g290(.A1(new_n464), .A2(new_n467), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(G127gat), .A2(G134gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(G127gat), .A2(G134gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G113gat), .B(G120gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G120gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G113gat), .ZN(new_n501));
  INV_X1    g300(.A(G113gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(G120gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G127gat), .B(G134gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n499), .A2(new_n506), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n486), .B1(new_n489), .B2(new_n484), .ZN(new_n510));
  AND4_X1   g309(.A1(new_n484), .A2(new_n481), .A3(new_n483), .A4(new_n486), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n475), .B(new_n477), .C1(new_n512), .C2(new_n479), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n458), .A2(new_n463), .A3(KEYINPUT25), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n466), .B1(new_n465), .B2(new_n462), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n509), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT68), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT34), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G43gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n519), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(new_n508), .B2(new_n517), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n527), .B2(KEYINPUT32), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT67), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n492), .A2(new_n507), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n509), .A3(new_n516), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n519), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n532), .B2(KEYINPUT33), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(KEYINPUT67), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n518), .A2(KEYINPUT68), .A3(new_n519), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n527), .B(KEYINPUT32), .C1(new_n534), .C2(new_n525), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n522), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n538), .ZN(new_n542));
  INV_X1    g341(.A(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n545), .A3(new_n521), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT4), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n509), .A2(new_n406), .A3(new_n548), .A4(new_n411), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT79), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT4), .B1(new_n412), .B2(new_n507), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT79), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n426), .A2(new_n552), .A3(new_n548), .A4(new_n509), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G225gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT78), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n509), .B1(new_n426), .B2(new_n414), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n412), .A2(KEYINPUT3), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT5), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n426), .B(new_n509), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n556), .ZN(new_n563));
  AOI211_X1 g362(.A(KEYINPUT5), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT81), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT81), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n426), .A2(new_n566), .A3(new_n548), .A4(new_n509), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n551), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n560), .A2(new_n563), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G1gat), .B(G29gat), .Z(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G85gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT6), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n569), .A2(new_n574), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  INV_X1    g379(.A(new_n390), .ZN(new_n581));
  NAND2_X1  g380(.A1(G226gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT29), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n492), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n513), .A2(KEYINPUT72), .A3(new_n516), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n492), .A2(new_n582), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n581), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n583), .A3(new_n588), .ZN(new_n593));
  INV_X1    g392(.A(new_n416), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n492), .A2(new_n582), .A3(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n390), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G8gat), .B(G36gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(G64gat), .B(G92gat), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n597), .B(new_n598), .Z(new_n599));
  NAND4_X1  g398(.A1(new_n591), .A2(new_n592), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n591), .A2(new_n596), .A3(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT30), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n599), .B(KEYINPUT73), .Z(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n591), .B2(new_n596), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n600), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n580), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n450), .A2(new_n547), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT35), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n449), .A2(new_n446), .B1(new_n541), .B2(new_n546), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(KEYINPUT85), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT85), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n612), .B(new_n600), .C1(new_n602), .C2(new_n604), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT86), .B1(new_n569), .B2(new_n574), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT86), .ZN(new_n616));
  INV_X1    g415(.A(new_n574), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n509), .A2(new_n406), .A3(new_n411), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n406), .A2(new_n411), .B1(new_n499), .B2(new_n506), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n556), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT5), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n554), .B2(new_n559), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n568), .A2(new_n561), .A3(new_n559), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n616), .B(new_n617), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n615), .A2(new_n624), .A3(new_n578), .A4(new_n577), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT35), .B1(new_n625), .B2(new_n576), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n614), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT69), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n547), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT69), .B(KEYINPUT36), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n541), .A2(new_n546), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n615), .A2(new_n624), .ZN(new_n636));
  INV_X1    g435(.A(new_n556), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n557), .A2(new_n558), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n637), .B1(new_n568), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n617), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT39), .B1(new_n562), .B2(new_n556), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT40), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n641), .B(new_n645), .C1(new_n639), .C2(new_n642), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n636), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n611), .A2(new_n647), .A3(new_n613), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n390), .B1(new_n589), .B2(new_n590), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n593), .A2(new_n581), .A3(new_n595), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(KEYINPUT37), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT37), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n591), .A2(new_n652), .A3(new_n596), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n603), .A2(KEYINPUT38), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n655), .A2(new_n601), .ZN(new_n656));
  INV_X1    g455(.A(new_n599), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n652), .B1(new_n591), .B2(new_n596), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT38), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n656), .A2(new_n660), .A3(new_n576), .A4(new_n625), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n648), .A2(new_n450), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n446), .A2(new_n606), .A3(new_n449), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n635), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT87), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n628), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n665), .B1(new_n628), .B2(new_n664), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n276), .B(new_n371), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT98), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT35), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n610), .B2(new_n607), .ZN(new_n672));
  AND4_X1   g471(.A1(new_n450), .A2(new_n547), .A3(new_n614), .A4(new_n626), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n541), .A2(new_n546), .A3(new_n633), .ZN(new_n674));
  INV_X1    g473(.A(new_n630), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n541), .B2(new_n546), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n663), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n648), .A2(new_n450), .A3(new_n661), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n672), .A2(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(KEYINPUT87), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n666), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n276), .A4(new_n371), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n670), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n580), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(G1gat), .ZN(G1324gat));
  INV_X1    g486(.A(new_n614), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT16), .B(G8gat), .Z(new_n689));
  AND4_X1   g488(.A1(KEYINPUT42), .A2(new_n684), .A3(new_n688), .A4(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT99), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n691), .B1(new_n684), .B2(new_n688), .ZN(new_n692));
  AOI211_X1 g491(.A(KEYINPUT99), .B(new_n614), .C1(new_n670), .C2(new_n683), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(G8gat), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT100), .A4(new_n208), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(new_n684), .ZN(new_n702));
  INV_X1    g501(.A(new_n547), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n702), .A2(G15gat), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(G15gat), .B1(new_n702), .B2(new_n635), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n450), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n684), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n351), .ZN(new_n711));
  INV_X1    g510(.A(new_n370), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n711), .A2(new_n312), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT101), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n681), .A2(new_n276), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(new_n214), .A3(new_n685), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT45), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT44), .B(new_n711), .C1(new_n667), .C2(new_n668), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n351), .B1(new_n628), .B2(new_n664), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n722));
  INV_X1    g521(.A(new_n275), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n265), .B1(new_n258), .B2(KEYINPUT18), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n272), .B1(new_n724), .B2(new_n261), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n274), .A2(KEYINPUT102), .A3(new_n275), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(new_n313), .A3(new_n370), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n721), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n580), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n717), .A2(new_n731), .ZN(G1328gat));
  OAI21_X1  g531(.A(G36gat), .B1(new_n730), .B2(new_n614), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n715), .A2(new_n215), .A3(new_n688), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(KEYINPUT103), .A3(KEYINPUT46), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n734), .B2(KEYINPUT46), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n733), .B1(KEYINPUT46), .B2(new_n734), .C1(new_n736), .C2(new_n737), .ZN(G1329gat));
  NOR2_X1   g537(.A1(new_n703), .A2(G43gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n715), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT47), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n715), .B2(new_n739), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT105), .B1(new_n745), .B2(KEYINPUT47), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G43gat), .B1(new_n730), .B2(new_n635), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n740), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n747), .B(new_n749), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n243), .B1(new_n730), .B2(new_n450), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n450), .A2(new_n243), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT106), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n715), .A2(new_n757), .ZN(new_n758));
  AOI211_X1 g557(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n758), .ZN(new_n759));
  AND4_X1   g558(.A1(new_n751), .A2(new_n755), .A3(new_n752), .A4(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1331gat));
  INV_X1    g560(.A(new_n352), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n679), .A2(new_n762), .A3(new_n370), .A4(new_n728), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n580), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n284), .ZN(G1332gat));
  INV_X1    g564(.A(new_n763), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n614), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT108), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n769), .B(new_n770), .Z(G1333gat));
  NOR2_X1   g570(.A1(new_n763), .A2(new_n703), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n774));
  AOI21_X1  g573(.A(G71gat), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n635), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n766), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n775), .B1(G71gat), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n766), .A2(new_n707), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  INV_X1    g580(.A(new_n728), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(new_n313), .A3(new_n712), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n721), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n580), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n782), .A2(new_n313), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n679), .A2(KEYINPUT51), .A3(new_n711), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n719), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n786), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n719), .B2(new_n786), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n685), .A2(new_n321), .A3(new_n370), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n785), .A2(new_n321), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n784), .B2(new_n614), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n794), .B1(new_n789), .B2(new_n791), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n688), .A2(new_n322), .A3(new_n370), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n795), .A2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n803), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n784), .B2(new_n635), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n703), .A2(G99gat), .A3(new_n712), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n795), .B2(new_n808), .ZN(G1338gat));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n791), .ZN(new_n810));
  INV_X1    g609(.A(new_n794), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n450), .A2(G106gat), .A3(new_n712), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(KEYINPUT112), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  INV_X1    g614(.A(new_n813), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n799), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n718), .A2(new_n707), .A3(new_n720), .A4(new_n783), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(new_n819), .C1(new_n795), .C2(new_n816), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT113), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n821), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(G1339gat));
  NAND2_X1  g627(.A1(new_n371), .A2(new_n728), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n362), .A2(new_n363), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n353), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n362), .A2(new_n363), .A3(new_n354), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n369), .B1(new_n364), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n366), .A2(new_n369), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n833), .A2(new_n835), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n836), .B1(new_n842), .B2(KEYINPUT115), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n839), .A2(new_n844), .A3(new_n840), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n248), .A2(new_n264), .A3(new_n263), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n252), .A2(new_n255), .ZN(new_n848));
  INV_X1    g647(.A(new_n248), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n249), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n271), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n349), .A2(new_n275), .A3(new_n350), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n843), .A2(new_n726), .A3(new_n727), .A4(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n275), .A2(new_n370), .A3(new_n852), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n275), .A2(new_n370), .A3(KEYINPUT116), .A4(new_n852), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n854), .B1(new_n861), .B2(new_n351), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n829), .B1(new_n862), .B2(new_n313), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n580), .ZN(new_n865));
  INV_X1    g664(.A(new_n610), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n688), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n276), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n782), .A2(new_n502), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT117), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n871), .B1(new_n869), .B2(new_n873), .ZN(G1340gat));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n370), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g675(.A1(new_n868), .A2(new_n313), .ZN(new_n877));
  XNOR2_X1  g676(.A(KEYINPUT118), .B(G127gat), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n877), .B(new_n878), .ZN(G1342gat));
  NAND2_X1  g678(.A1(new_n868), .A2(new_n711), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n880), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT56), .B1(new_n880), .B2(G134gat), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(G134gat), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n396), .A2(new_n398), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n776), .A2(new_n580), .A3(new_n688), .ZN(new_n886));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n863), .B2(new_n707), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(new_n842), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n836), .B(KEYINPUT119), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n276), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n711), .B1(new_n856), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n312), .B1(new_n892), .B2(new_n854), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n888), .B(new_n450), .C1(new_n893), .C2(new_n829), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n886), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n885), .B1(new_n895), .B2(new_n870), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n776), .A2(new_n450), .A3(new_n688), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n870), .A2(G141gat), .ZN(new_n899));
  AND4_X1   g698(.A1(new_n685), .A2(new_n863), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n782), .B(new_n886), .C1(new_n887), .C2(new_n894), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n885), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n901), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(KEYINPUT58), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n900), .B1(new_n904), .B2(new_n885), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT120), .A3(new_n897), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n902), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n912), .B(new_n902), .C1(new_n907), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  AND2_X1   g713(.A1(new_n865), .A2(new_n898), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n408), .A3(new_n370), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n895), .A2(new_n712), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n917), .A2(KEYINPUT59), .A3(new_n408), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT57), .B1(new_n864), .B2(new_n450), .ZN(new_n920));
  INV_X1    g719(.A(new_n371), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n893), .B1(new_n276), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n888), .A3(new_n707), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n920), .A2(new_n370), .A3(new_n886), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n919), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n916), .B1(new_n918), .B2(new_n925), .ZN(G1345gat));
  NAND3_X1  g725(.A1(new_n915), .A2(new_n404), .A3(new_n313), .ZN(new_n927));
  OAI21_X1  g726(.A(G155gat), .B1(new_n895), .B2(new_n312), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1346gat));
  NOR3_X1   g728(.A1(new_n895), .A2(new_n403), .A3(new_n351), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n711), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n403), .B2(new_n931), .ZN(G1347gat));
  NAND2_X1  g731(.A1(new_n688), .A2(new_n580), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n864), .A2(new_n866), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n453), .A3(new_n782), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT122), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n453), .B1(new_n934), .B2(new_n276), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n936), .A2(new_n937), .ZN(G1348gat));
  NAND2_X1  g737(.A1(new_n934), .A2(new_n370), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g739(.A1(new_n934), .A2(new_n313), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n480), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n942), .B1(new_n489), .B2(new_n941), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1350gat));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n934), .A2(new_n711), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n948), .A3(G190gat), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n947), .B2(G190gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n951), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT61), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n946), .B(new_n956), .C1(new_n950), .C2(new_n951), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n957), .C1(G190gat), .C2(new_n947), .ZN(G1351gat));
  NOR2_X1   g757(.A1(new_n776), .A2(new_n933), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n920), .A2(new_n923), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(G197gat), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n960), .A2(new_n961), .A3(new_n870), .ZN(new_n962));
  INV_X1    g761(.A(new_n959), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n864), .A2(new_n450), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT126), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n782), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n962), .B1(new_n967), .B2(new_n961), .ZN(G1352gat));
  INV_X1    g767(.A(G204gat), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n969), .A3(new_n370), .ZN(new_n970));
  XOR2_X1   g769(.A(new_n970), .B(KEYINPUT62), .Z(new_n971));
  NAND3_X1  g770(.A1(new_n920), .A2(new_n370), .A3(new_n923), .ZN(new_n972));
  OAI21_X1  g771(.A(G204gat), .B1(new_n972), .B2(new_n963), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n973), .ZN(G1353gat));
  NAND3_X1  g773(.A1(new_n966), .A2(new_n385), .A3(new_n313), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n960), .A2(new_n312), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n960), .B2(new_n351), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n711), .A2(new_n386), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n965), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


