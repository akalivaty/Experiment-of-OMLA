//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n209));
  INV_X1    g008(.A(G1gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n209), .B1(KEYINPUT92), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(KEYINPUT92), .B2(new_n210), .ZN(new_n212));
  INV_X1    g011(.A(G15gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(G22gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n215), .A2(G15gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT91), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(G15gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT91), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n212), .A2(new_n217), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(G1gat), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  OAI21_X1  g022(.A(G8gat), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n220), .B1(new_n218), .B2(new_n219), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n210), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n217), .A3(new_n221), .ZN(new_n228));
  INV_X1    g027(.A(G8gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT88), .A2(G29gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G36gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT89), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT88), .B(G29gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(G36gat), .ZN(new_n238));
  INV_X1    g037(.A(G29gat), .ZN(new_n239));
  INV_X1    g038(.A(G36gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT14), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT14), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(G29gat), .B2(G36gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n235), .A2(new_n238), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G43gat), .ZN(new_n247));
  INV_X1    g046(.A(G50gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G43gat), .A2(G50gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT15), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT90), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n241), .A2(new_n243), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT15), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n256), .A3(new_n250), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n253), .A2(new_n252), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n235), .A2(new_n238), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n246), .A2(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT17), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n238), .A3(new_n245), .ZN(new_n262));
  INV_X1    g061(.A(new_n252), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT17), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n264), .B(new_n265), .C1(new_n259), .C2(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n231), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n229), .B1(new_n227), .B2(new_n228), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n258), .ZN(new_n272));
  INV_X1    g071(.A(new_n259), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n272), .A2(new_n273), .B1(new_n262), .B2(new_n263), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n268), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  AOI211_X1 g075(.A(new_n268), .B(new_n231), .C1(new_n261), .C2(new_n266), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT18), .B(new_n208), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n231), .B(new_n260), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n208), .B(KEYINPUT13), .Z(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n267), .A2(KEYINPUT93), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(new_n267), .B2(new_n275), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n284), .B1(new_n286), .B2(new_n208), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n207), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n208), .B1(new_n276), .B2(new_n277), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(new_n283), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n290), .A2(new_n206), .A3(new_n278), .A4(new_n281), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT38), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296));
  NOR2_X1   g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  AND2_X1   g103(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(G190gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n296), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n302), .A2(new_n296), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(KEYINPUT64), .A3(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n303), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT64), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n307), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT26), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n303), .B(new_n319), .C1(new_n321), .C2(new_n297), .ZN(new_n322));
  INV_X1    g121(.A(G183gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT27), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT27), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G183gat), .ZN(new_n326));
  INV_X1    g125(.A(G190gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT28), .A4(new_n327), .ZN(new_n331));
  AOI211_X1 g130(.A(new_n316), .B(new_n322), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  INV_X1    g132(.A(new_n322), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT65), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n315), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT71), .ZN(new_n337));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n339), .A2(KEYINPUT29), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(new_n315), .C1(new_n332), .C2(new_n335), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n333), .A2(new_n334), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n315), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n339), .ZN(new_n346));
  INV_X1    g145(.A(G197gat), .ZN(new_n347));
  INV_X1    g146(.A(G204gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351));
  NAND2_X1  g150(.A1(G211gat), .A2(G218gat), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n349), .A2(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(G211gat), .A2(G218gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT70), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n356), .B1(new_n355), .B2(new_n352), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n354), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n353), .A3(new_n357), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n346), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT37), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n316), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n333), .A2(KEYINPUT65), .A3(new_n334), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n341), .B1(new_n369), .B2(new_n315), .ZN(new_n370));
  INV_X1    g169(.A(new_n342), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n339), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n345), .A2(KEYINPUT29), .A3(new_n339), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n364), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n295), .B1(new_n366), .B2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n343), .A2(new_n346), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n363), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(new_n374), .A3(new_n364), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  NOR3_X1   g184(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT75), .Z(new_n388));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389));
  INV_X1    g188(.A(G113gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT66), .A3(G120gat), .ZN(new_n391));
  INV_X1    g190(.A(G134gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G127gat), .ZN(new_n393));
  INV_X1    g192(.A(G127gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G134gat), .ZN(new_n395));
  AND4_X1   g194(.A1(new_n389), .A2(new_n391), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n390), .A2(G120gat), .ZN(new_n400));
  INV_X1    g199(.A(G120gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(G113gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n389), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(new_n395), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n396), .A2(new_n399), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g204(.A1(G141gat), .A2(G148gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT73), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(G141gat), .ZN(new_n409));
  INV_X1    g208(.A(G148gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT73), .ZN(new_n412));
  NAND2_X1  g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT74), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(G155gat), .ZN(new_n422));
  INV_X1    g221(.A(G162gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT74), .ZN(new_n425));
  NAND2_X1  g224(.A1(G155gat), .A2(G162gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n406), .A2(new_n407), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(KEYINPUT2), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n421), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n405), .A2(new_n420), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n396), .A2(new_n399), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n403), .A2(new_n404), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n420), .A2(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n388), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n436));
  INV_X1    g235(.A(new_n419), .ZN(new_n437));
  XNOR2_X1  g236(.A(G141gat), .B(G148gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT2), .B1(new_n438), .B2(KEYINPUT73), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n437), .B1(new_n439), .B2(new_n414), .ZN(new_n440));
  AND4_X1   g239(.A1(new_n428), .A2(new_n421), .A3(new_n427), .A4(new_n429), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT3), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n443), .A3(new_n430), .ZN(new_n444));
  INV_X1    g243(.A(new_n405), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n388), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n405), .A2(new_n420), .A3(new_n430), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n421), .A2(new_n428), .A3(new_n429), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n451), .A2(new_n427), .B1(new_n416), .B2(new_n419), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n446), .A2(new_n447), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n448), .A2(new_n449), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT4), .B1(new_n452), .B2(new_n405), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(KEYINPUT5), .A3(new_n447), .A4(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g259(.A(G1gat), .B(G29gat), .Z(new_n461));
  XNOR2_X1  g260(.A(G57gat), .B(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n455), .A2(new_n459), .A3(new_n465), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n455), .A2(new_n459), .A3(new_n465), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n455), .B2(new_n459), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(KEYINPUT6), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n338), .B1(new_n337), .B2(new_n342), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n474), .A2(new_n363), .A3(new_n373), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n364), .B1(new_n343), .B2(new_n346), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n385), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n470), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n294), .B1(new_n386), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT6), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n460), .A2(new_n468), .A3(new_n466), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n377), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  INV_X1    g282(.A(new_n385), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n363), .B1(new_n474), .B2(new_n373), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT37), .A3(new_n365), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(new_n295), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n477), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n380), .A2(KEYINPUT37), .A3(new_n381), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n489), .A3(new_n484), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT38), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n488), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G78gat), .B(G106gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(KEYINPUT31), .B(G50gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n496), .B(new_n497), .Z(new_n498));
  OAI21_X1  g297(.A(new_n443), .B1(new_n363), .B2(KEYINPUT29), .ZN(new_n499));
  INV_X1    g298(.A(new_n452), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n364), .B1(new_n502), .B2(new_n444), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n444), .A2(new_n502), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n363), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT77), .ZN(new_n508));
  INV_X1    g307(.A(G228gat), .ZN(new_n509));
  INV_X1    g308(.A(G233gat), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n505), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n509), .A2(new_n510), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n501), .A4(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n511), .A2(new_n515), .A3(new_n215), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n215), .B1(new_n511), .B2(new_n515), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n498), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT79), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n520), .B(new_n498), .C1(new_n516), .C2(new_n517), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n517), .A2(new_n498), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT80), .A4(new_n215), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n511), .A2(new_n515), .A3(new_n215), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(new_n388), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n529), .B2(new_n388), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n431), .A2(new_n434), .A3(new_n388), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT39), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n531), .B2(new_n532), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n537), .A2(KEYINPUT84), .A3(new_n466), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT84), .B1(new_n537), .B2(new_n466), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT40), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n484), .B1(new_n380), .B2(new_n381), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT30), .B1(new_n543), .B2(KEYINPUT72), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n380), .A2(new_n381), .A3(new_n484), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n477), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT40), .B(new_n535), .C1(new_n538), .C2(new_n539), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n542), .A2(new_n469), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n495), .A2(new_n528), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n528), .A2(KEYINPUT81), .ZN(new_n553));
  INV_X1    g352(.A(new_n549), .ZN(new_n554));
  INV_X1    g353(.A(new_n482), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT81), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n519), .A2(new_n527), .A3(new_n557), .A4(new_n521), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n553), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n405), .A2(KEYINPUT67), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n369), .A2(new_n315), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n405), .A2(KEYINPUT67), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n336), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G227gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(new_n510), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n560), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT34), .Z(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n568), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT33), .B1(new_n566), .B2(new_n568), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT68), .B(G71gat), .Z(new_n573));
  INV_X1    g372(.A(G99gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G15gat), .B(G43gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(KEYINPUT32), .B(new_n571), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n572), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n571), .A2(KEYINPUT32), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n570), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n579), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n569), .B(KEYINPUT34), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n583), .A2(KEYINPUT36), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT36), .B1(new_n583), .B2(new_n586), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n552), .A2(new_n559), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n528), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT35), .B1(new_n592), .B2(new_n556), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n549), .A2(new_n482), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n594), .A2(new_n528), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n293), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n422), .ZN(new_n600));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G71gat), .A2(G78gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  AOI22_X1  g406(.A1(KEYINPUT95), .A2(new_n606), .B1(new_n607), .B2(new_n604), .ZN(new_n608));
  INV_X1    g407(.A(G64gat), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(G57gat), .ZN(new_n610));
  INV_X1    g409(.A(G57gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(G64gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n606), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(G64gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(G57gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n606), .B(new_n617), .C1(new_n620), .C2(KEYINPUT95), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n614), .A2(new_n621), .ZN(new_n626));
  OAI211_X1 g425(.A(G231gat), .B(G233gat), .C1(new_n626), .C2(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(G127gat), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n271), .B1(new_n623), .B2(new_n622), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n394), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n629), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n603), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n631), .ZN(new_n635));
  INV_X1    g434(.A(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n602), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT96), .Z(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n261), .A2(new_n266), .ZN(new_n648));
  NAND2_X1  g447(.A1(G85gat), .A2(G92gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT7), .ZN(new_n650));
  NAND2_X1  g449(.A1(G99gat), .A2(G106gat), .ZN(new_n651));
  INV_X1    g450(.A(G85gat), .ZN(new_n652));
  INV_X1    g451(.A(G92gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(KEYINPUT8), .A2(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G99gat), .B(G106gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n650), .A3(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n648), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G190gat), .B(G218gat), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT97), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n642), .B2(new_n641), .ZN(new_n667));
  INV_X1    g466(.A(new_n660), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n260), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n665), .B1(new_n661), .B2(new_n669), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n647), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n661), .A2(new_n669), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n664), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n646), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n640), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT98), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n640), .A2(new_n673), .A3(new_n676), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n656), .A2(KEYINPUT99), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n626), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n660), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n626), .A2(new_n657), .A3(new_n659), .A4(new_n683), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n668), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n685), .A2(new_n687), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n682), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G120gat), .B(G148gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(G176gat), .B(G204gat), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n691), .A2(new_n693), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n678), .A2(new_n680), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n598), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n555), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n210), .ZN(G1324gat));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n554), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G8gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n229), .B2(new_n707), .ZN(new_n711));
  MUX2_X1   g510(.A(new_n710), .B(new_n711), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g511(.A(G15gat), .B1(new_n704), .B2(new_n589), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n591), .A2(new_n213), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n704), .B2(new_n714), .ZN(G1326gat));
  NAND2_X1  g514(.A1(new_n553), .A2(new_n558), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n704), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  NOR2_X1   g518(.A1(new_n701), .A2(new_n640), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n673), .A2(new_n676), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n598), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n236), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n482), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n590), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n552), .A2(KEYINPUT101), .A3(new_n559), .A4(new_n589), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n597), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n722), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI211_X1 g535(.A(new_n735), .B(new_n723), .C1(new_n590), .C2(new_n597), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n293), .A2(new_n721), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n736), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g539(.A1(new_n740), .A2(new_n482), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n729), .B1(new_n741), .B2(new_n727), .ZN(G1328gat));
  NOR3_X1   g541(.A1(new_n725), .A2(G36gat), .A3(new_n554), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT46), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n740), .A2(new_n549), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n240), .ZN(G1329gat));
  INV_X1    g545(.A(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n591), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n583), .A2(new_n586), .A3(KEYINPUT36), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n736), .A2(new_n750), .A3(new_n738), .A4(new_n739), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n726), .A2(new_n247), .A3(new_n591), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT47), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n753), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n757), .B1(new_n751), .B2(G43gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(KEYINPUT102), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n760), .ZN(G1330gat));
  NOR3_X1   g560(.A1(new_n725), .A2(G50gat), .A3(new_n716), .ZN(new_n762));
  INV_X1    g561(.A(new_n716), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n764), .B2(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n528), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n248), .B1(new_n740), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n765), .A2(KEYINPUT48), .B1(new_n767), .B2(new_n769), .ZN(G1331gat));
  NAND4_X1  g569(.A1(new_n293), .A2(new_n678), .A3(new_n680), .A4(new_n701), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n732), .A2(new_n597), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n590), .A2(new_n730), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n482), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n549), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT49), .B(G64gat), .Z(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(new_n779), .ZN(G1333gat));
  NAND2_X1  g579(.A1(new_n774), .A2(new_n750), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G71gat), .ZN(new_n782));
  INV_X1    g581(.A(G71gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n774), .A2(new_n783), .A3(new_n591), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n763), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n597), .A3(new_n732), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n292), .A2(new_n640), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n722), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n789), .A2(KEYINPUT51), .A3(new_n722), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n702), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n652), .A3(new_n482), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n292), .A2(new_n640), .A3(new_n702), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n723), .B1(new_n772), .B2(new_n773), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n738), .B(new_n799), .C1(new_n800), .C2(KEYINPUT44), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT103), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n736), .A2(KEYINPUT103), .A3(new_n738), .A4(new_n799), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n803), .A2(new_n482), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n652), .B2(new_n805), .ZN(G1336gat));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(G92gat), .C1(new_n801), .C2(new_n554), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(KEYINPUT105), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n549), .A2(new_n653), .A3(new_n701), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT104), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n808), .B(new_n809), .C1(new_n796), .C2(new_n811), .ZN(new_n812));
  AOI211_X1 g611(.A(KEYINPUT105), .B(new_n811), .C1(new_n793), .C2(new_n794), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n803), .A2(new_n549), .A3(new_n804), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(G92gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(new_n807), .ZN(G1337gat));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n574), .A3(new_n591), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n803), .A2(new_n750), .A3(new_n804), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n574), .B2(new_n818), .ZN(G1338gat));
  NOR3_X1   g618(.A1(new_n528), .A2(G106gat), .A3(new_n702), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT106), .Z(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n795), .A2(KEYINPUT107), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G106gat), .B1(new_n801), .B2(new_n528), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n803), .A2(new_n763), .A3(new_n804), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(KEYINPUT53), .A3(G106gat), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n795), .A2(new_n822), .B1(KEYINPUT107), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(G1339gat));
  INV_X1    g629(.A(new_n640), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n688), .A2(new_n682), .A3(new_n689), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n691), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n697), .B1(new_n690), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n700), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n292), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g640(.A1(new_n286), .A2(new_n208), .B1(new_n279), .B2(new_n280), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n205), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n291), .A2(new_n701), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n722), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n840), .A2(new_n291), .A3(new_n722), .A4(new_n843), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n831), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n703), .A2(new_n293), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n763), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n482), .A3(new_n554), .A4(new_n591), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n390), .A3(new_n293), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n555), .B1(new_n848), .B2(new_n849), .ZN(new_n853));
  INV_X1    g652(.A(new_n592), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(KEYINPUT108), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(KEYINPUT108), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n554), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n292), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n852), .B1(new_n860), .B2(new_n390), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n851), .A2(new_n401), .A3(new_n702), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n701), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n401), .ZN(G1341gat));
  OAI21_X1  g663(.A(G127gat), .B1(new_n851), .B2(new_n831), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n640), .A2(new_n394), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n858), .B2(new_n866), .ZN(G1342gat));
  NAND3_X1  g666(.A1(new_n859), .A2(new_n392), .A3(new_n722), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n870));
  OAI21_X1  g669(.A(G134gat), .B1(new_n851), .B2(new_n723), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G1343gat));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n874));
  XOR2_X1   g673(.A(new_n874), .B(KEYINPUT116), .Z(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n750), .A2(new_n549), .A3(new_n528), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n853), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n292), .A2(new_n409), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT114), .Z(new_n880));
  NOR2_X1   g679(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n848), .A2(new_n849), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT57), .B1(new_n882), .B2(new_n766), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n763), .A2(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n688), .A2(new_n682), .A3(new_n689), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(new_n690), .A3(new_n834), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n688), .A2(new_n689), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n834), .A3(new_n681), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n698), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n885), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n833), .A2(KEYINPUT110), .A3(new_n835), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n837), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT111), .ZN(new_n894));
  INV_X1    g693(.A(new_n838), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n891), .A2(new_n892), .A3(new_n896), .A4(new_n837), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n292), .A2(new_n894), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n722), .B1(new_n898), .B2(new_n844), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n846), .B1(new_n899), .B2(KEYINPUT112), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT112), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n901), .B(new_n722), .C1(new_n898), .C2(new_n844), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n831), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n884), .B1(new_n903), .B2(new_n849), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n883), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n844), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n894), .A2(new_n897), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n838), .B1(new_n288), .B2(new_n291), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n901), .B1(new_n910), .B2(new_n722), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n899), .A2(KEYINPUT112), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n846), .A3(new_n912), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n913), .A2(new_n831), .B1(new_n293), .B2(new_n703), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT113), .B1(new_n914), .B2(new_n884), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n750), .A2(new_n555), .A3(new_n549), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT109), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n916), .A2(new_n292), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n881), .B1(new_n919), .B2(G141gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n873), .A2(KEYINPUT58), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n876), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n921), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT109), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n917), .B(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n925), .B1(new_n906), .B2(new_n915), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n409), .B1(new_n926), .B2(new_n292), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n923), .B(new_n875), .C1(new_n927), .C2(new_n881), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n922), .A2(new_n928), .ZN(G1344gat));
  INV_X1    g728(.A(new_n878), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n410), .A3(new_n701), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT117), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n701), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n882), .A2(KEYINPUT57), .A3(new_n766), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT57), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n703), .A2(new_n938), .A3(new_n293), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n678), .A2(new_n680), .A3(new_n702), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT119), .B1(new_n940), .B2(new_n292), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n846), .B1(new_n910), .B2(new_n722), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n831), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n937), .B1(new_n944), .B2(new_n716), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n936), .B1(new_n945), .B2(KEYINPUT120), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n947), .B(new_n937), .C1(new_n944), .C2(new_n716), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n934), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n933), .B(KEYINPUT59), .C1(new_n949), .C2(new_n410), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n939), .A2(new_n941), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n831), .B1(new_n899), .B2(new_n847), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n716), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT120), .B1(new_n953), .B2(KEYINPUT57), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n948), .A3(new_n935), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n925), .A2(new_n702), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n410), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT121), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(G148gat), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n960), .B1(new_n926), .B2(new_n701), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n950), .B(new_n959), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n932), .B1(new_n963), .B2(new_n964), .ZN(G1345gat));
  NAND3_X1  g764(.A1(new_n930), .A2(new_n422), .A3(new_n640), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n926), .A2(new_n640), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n422), .ZN(G1346gat));
  AOI21_X1  g767(.A(G162gat), .B1(new_n930), .B2(new_n722), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n723), .A2(new_n423), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n926), .B2(new_n970), .ZN(G1347gat));
  AOI21_X1  g770(.A(new_n482), .B1(new_n848), .B2(new_n849), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n972), .A2(new_n549), .A3(new_n854), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G169gat), .B1(new_n974), .B2(new_n292), .ZN(new_n975));
  NAND4_X1  g774(.A1(new_n850), .A2(new_n555), .A3(new_n549), .A4(new_n591), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n976), .A2(new_n317), .A3(new_n293), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n975), .A2(new_n977), .ZN(G1348gat));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n318), .A3(new_n701), .ZN(new_n979));
  OAI21_X1  g778(.A(G176gat), .B1(new_n976), .B2(new_n702), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1349gat));
  NAND4_X1  g780(.A1(new_n974), .A2(new_n324), .A3(new_n326), .A4(new_n640), .ZN(new_n982));
  OAI21_X1  g781(.A(G183gat), .B1(new_n976), .B2(new_n831), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n985));
  XOR2_X1   g784(.A(new_n984), .B(new_n985), .Z(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n976), .B2(new_n723), .ZN(new_n987));
  XOR2_X1   g786(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n988));
  XNOR2_X1  g787(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n327), .A3(new_n722), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1351gat));
  NOR3_X1   g790(.A1(new_n750), .A2(new_n482), .A3(new_n554), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n955), .A2(new_n292), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n347), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n750), .A2(new_n554), .A3(new_n528), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT124), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n998), .A2(new_n972), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT125), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n292), .A2(new_n347), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(G1352gat));
  NAND3_X1  g801(.A1(new_n999), .A2(new_n348), .A3(new_n701), .ZN(new_n1003));
  XOR2_X1   g802(.A(new_n1003), .B(KEYINPUT62), .Z(new_n1004));
  NAND2_X1  g803(.A1(new_n955), .A2(new_n992), .ZN(new_n1005));
  OAI21_X1  g804(.A(G204gat), .B1(new_n1005), .B2(new_n702), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1353gat));
  NAND3_X1  g806(.A1(new_n955), .A2(new_n640), .A3(new_n992), .ZN(new_n1008));
  AND3_X1   g807(.A1(new_n1008), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1009));
  AOI21_X1  g808(.A(KEYINPUT63), .B1(new_n1008), .B2(G211gat), .ZN(new_n1010));
  OR2_X1    g809(.A1(new_n831), .A2(G211gat), .ZN(new_n1011));
  OAI22_X1  g810(.A1(new_n1009), .A2(new_n1010), .B1(new_n1000), .B2(new_n1011), .ZN(G1354gat));
  OAI21_X1  g811(.A(G218gat), .B1(new_n1005), .B2(new_n723), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n723), .A2(G218gat), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n1000), .B2(new_n1014), .ZN(G1355gat));
endmodule


