//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G97), .A2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n218), .B(new_n223), .C1(G107), .C2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G50), .ZN(new_n225));
  INV_X1    g0025(.A(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(G58), .A2(G232), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n212), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n210), .ZN(new_n234));
  AND2_X1   g0034(.A1(new_n206), .A2(G50), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n215), .B(new_n232), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n217), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n225), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  AND2_X1   g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  OAI21_X1  g0053(.A(KEYINPUT67), .B1(new_n253), .B2(new_n233), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  XOR2_X1   g0062(.A(new_n260), .B(KEYINPUT66), .Z(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(G274), .A3(new_n259), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G222), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G223), .A2(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n253), .A2(new_n233), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(new_n270), .C1(G77), .C2(new_n265), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n262), .A2(new_n264), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n276));
  INV_X1    g0076(.A(G150), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n210), .A2(new_n278), .A3(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(G20), .B2(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT68), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n278), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI221_X1 g0088(.A(new_n276), .B1(new_n277), .B2(new_n283), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n233), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n289), .A2(new_n291), .B1(new_n225), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n209), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n294), .B1(new_n225), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n273), .B(new_n275), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n299), .B2(new_n298), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n272), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n272), .A2(G179), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n298), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(G50), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT74), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n287), .A2(G77), .B1(G20), .B2(new_n202), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT73), .Z(new_n312));
  AOI21_X1  g0112(.A(new_n295), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT11), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n293), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT12), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n292), .B2(G68), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n317), .C1(new_n297), .C2(new_n202), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n318), .B(KEYINPUT75), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(KEYINPUT11), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n226), .A2(new_n266), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n265), .B(new_n323), .C1(G232), .C2(new_n266), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G97), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n278), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n270), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n261), .A2(G238), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(new_n264), .ZN(new_n330));
  XOR2_X1   g0130(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n331));
  OR2_X1    g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT72), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n330), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OR3_X1    g0135(.A1(new_n330), .A2(KEYINPUT72), .A3(new_n331), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G200), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n330), .A2(KEYINPUT13), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n332), .A2(G190), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n322), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(G169), .A3(new_n336), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n332), .A2(G179), .A3(new_n338), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n335), .A2(new_n336), .A3(new_n345), .A4(G169), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n341), .B1(new_n347), .B2(new_n321), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n308), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  AND2_X1   g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(KEYINPUT3), .A2(G33), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT7), .B1(new_n354), .B2(new_n210), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  NOR4_X1   g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .A4(G20), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G58), .A2(G68), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n203), .A2(new_n205), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(new_n282), .B2(G159), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n358), .A2(KEYINPUT76), .A3(KEYINPUT16), .A4(new_n361), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n356), .B1(new_n265), .B2(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n354), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n202), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n360), .A2(G20), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n282), .A2(G159), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n370), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n358), .A2(new_n361), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n366), .A2(KEYINPUT78), .A3(new_n291), .A4(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT78), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT77), .B1(new_n377), .B2(new_n367), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n375), .B(KEYINPUT16), .C1(new_n358), .C2(new_n361), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n364), .A2(new_n291), .A3(new_n365), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n265), .B1(G226), .B2(new_n266), .ZN(new_n387));
  NOR2_X1   g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n387), .A2(new_n388), .B1(new_n278), .B2(new_n221), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n270), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n261), .A2(G232), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(new_n264), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G190), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n284), .B(KEYINPUT68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n296), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT79), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n293), .A2(new_n291), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(new_n293), .B2(new_n286), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n380), .A2(new_n386), .A3(new_n394), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n392), .A2(G200), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n351), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n401), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT17), .A3(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n392), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G169), .B2(new_n392), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n380), .A2(new_n386), .A3(new_n400), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT80), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n380), .A2(new_n386), .A3(new_n412), .A4(new_n400), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n409), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(KEYINPUT81), .A2(KEYINPUT18), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n404), .B(new_n406), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n409), .B(new_n417), .C1(new_n411), .C2(new_n413), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT15), .B(G87), .Z(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n283), .B2(new_n284), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n291), .B1(new_n227), .B2(new_n293), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n227), .B2(new_n297), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT70), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n261), .A2(G244), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n266), .A2(G232), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n265), .B(new_n426), .C1(new_n220), .C2(new_n266), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n270), .C1(G107), .C2(new_n265), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n264), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n424), .B(new_n430), .C1(new_n274), .C2(new_n429), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n304), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n423), .B(new_n432), .C1(G179), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n416), .A2(new_n418), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n350), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G116), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n438), .A2(G20), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n210), .B(G87), .C1(new_n352), .C2(new_n353), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT22), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT22), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n265), .A2(new_n442), .A3(new_n210), .A4(G87), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n210), .A2(G107), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT23), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT24), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n444), .A2(KEYINPUT24), .A3(new_n446), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n291), .A3(new_n449), .ZN(new_n450));
  OR3_X1    g0250(.A1(new_n292), .A2(KEYINPUT25), .A3(G107), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT25), .B1(new_n292), .B2(G107), .ZN(new_n452));
  INV_X1    g0252(.A(G107), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n209), .A2(G33), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n292), .A2(new_n454), .A3(new_n233), .A4(new_n290), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n451), .B(new_n452), .C1(new_n453), .C2(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT89), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n209), .A2(G45), .ZN(new_n460));
  OR2_X1    g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n253), .A2(KEYINPUT67), .A3(new_n233), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n463), .B(G274), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n265), .A2(G257), .A3(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G294), .ZN(new_n468));
  OAI21_X1  g0268(.A(G250), .B1(new_n352), .B2(new_n353), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n467), .B1(new_n278), .B2(new_n468), .C1(G1698), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n270), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  INV_X1    g0273(.A(new_n462), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G264), .B(new_n476), .C1(new_n464), .C2(new_n465), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT5), .B(G41), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n254), .A2(new_n258), .B1(new_n479), .B2(new_n473), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT90), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(G264), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT91), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n478), .B2(new_n482), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n466), .B(new_n471), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(G200), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n477), .A2(KEYINPUT90), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n481), .B1(new_n480), .B2(G264), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n471), .B(new_n466), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n491), .A2(G190), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n459), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n441), .A2(new_n443), .ZN(new_n494));
  INV_X1    g0294(.A(new_n439), .ZN(new_n495));
  AND4_X1   g0295(.A1(KEYINPUT24), .A2(new_n494), .A3(new_n446), .A4(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n447), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n457), .B1(new_n497), .B2(new_n291), .ZN(new_n498));
  OAI21_X1  g0298(.A(KEYINPUT91), .B1(new_n489), .B2(new_n490), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(G179), .A3(new_n466), .A4(new_n471), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n491), .A2(G169), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n493), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n293), .A2(new_n326), .ZN(new_n506));
  INV_X1    g0306(.A(new_n455), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  NOR2_X1   g0309(.A1(KEYINPUT82), .A2(KEYINPUT6), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(G97), .B(G107), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT6), .A2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(KEYINPUT82), .B2(KEYINPUT6), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n518));
  OAI21_X1  g0318(.A(G107), .B1(new_n355), .B2(new_n357), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n509), .B1(new_n520), .B2(new_n291), .ZN(new_n521));
  AOI211_X1 g0321(.A(KEYINPUT83), .B(new_n295), .C1(new_n518), .C2(new_n519), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n506), .B(new_n508), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT4), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G1698), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(G244), .C1(new_n353), .C2(new_n352), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G283), .ZN(new_n527));
  OR2_X1    g0327(.A1(KEYINPUT3), .A2(G33), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT3), .A2(G33), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n228), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n526), .B(new_n527), .C1(new_n530), .C2(KEYINPUT4), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n266), .B1(new_n469), .B2(KEYINPUT4), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n270), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n480), .A2(G257), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n466), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n274), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n523), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(G200), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(G179), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n304), .B2(new_n535), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(new_n538), .B1(new_n523), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n292), .A2(G116), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n455), .A2(new_n216), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n216), .A2(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n291), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT88), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n291), .A2(KEYINPUT88), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n527), .B(new_n210), .C1(G33), .C2(new_n326), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT20), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI221_X4 g0353(.A(new_n548), .B1(new_n216), .B2(G20), .C1(new_n290), .C2(new_n233), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT88), .B1(new_n291), .B2(new_n546), .ZN(new_n555));
  OAI211_X1 g0355(.A(KEYINPUT20), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n543), .B(new_n545), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G264), .B(G1698), .C1(new_n352), .C2(new_n353), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT87), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT87), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n265), .A2(new_n561), .A3(G264), .A4(G1698), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n265), .A2(G257), .A3(new_n266), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n354), .A2(G303), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n560), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n270), .ZN(new_n566));
  OAI211_X1 g0366(.A(G270), .B(new_n476), .C1(new_n464), .C2(new_n465), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n466), .A2(new_n567), .A3(KEYINPUT86), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT86), .B1(new_n466), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n558), .A2(new_n570), .A3(G169), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n542), .B(new_n544), .C1(new_n576), .C2(new_n556), .ZN(new_n577));
  OAI211_X1 g0377(.A(G190), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n466), .A2(new_n567), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT86), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n466), .A2(new_n567), .A3(KEYINPUT86), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n581), .A2(new_n582), .B1(new_n270), .B2(new_n565), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n578), .C1(new_n583), .C2(new_n487), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n558), .A3(G179), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n558), .A2(new_n570), .A3(KEYINPUT21), .A4(G169), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n573), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n265), .A2(new_n210), .A3(G68), .ZN(new_n589));
  XOR2_X1   g0389(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n590));
  NOR2_X1   g0390(.A1(new_n288), .A2(new_n326), .ZN(new_n591));
  AOI21_X1  g0391(.A(G20), .B1(new_n590), .B2(new_n327), .ZN(new_n592));
  NOR3_X1   g0392(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n589), .B1(new_n590), .B2(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n419), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n594), .A2(new_n291), .B1(new_n293), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n507), .A2(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n460), .A2(new_n222), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n460), .A2(G274), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n259), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n259), .A2(KEYINPUT84), .A3(new_n599), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n220), .A2(new_n266), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n265), .B(new_n606), .C1(G244), .C2(new_n266), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n438), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n270), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n598), .B1(G200), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n603), .A2(new_n604), .B1(new_n270), .B2(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n610), .A2(new_n304), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n507), .A2(new_n419), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n596), .A2(new_n615), .B1(new_n612), .B2(new_n407), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n611), .A2(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n505), .A2(new_n541), .A3(new_n588), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n437), .A2(new_n618), .ZN(G372));
  INV_X1    g0419(.A(new_n307), .ZN(new_n620));
  INV_X1    g0420(.A(new_n409), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n410), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(KEYINPUT18), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n347), .A2(new_n321), .ZN(new_n625));
  XOR2_X1   g0425(.A(new_n433), .B(KEYINPUT92), .Z(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n340), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT93), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT93), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n625), .A2(new_n630), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n406), .A2(new_n404), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n624), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n620), .B1(new_n634), .B2(new_n303), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n611), .A2(new_n613), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n488), .A2(new_n492), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n498), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n537), .A2(new_n538), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n573), .A2(new_n585), .A3(new_n586), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n638), .B(new_n639), .C1(new_n504), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n540), .A2(new_n523), .ZN(new_n642));
  AOI211_X1 g0442(.A(KEYINPUT26), .B(new_n636), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n636), .B2(new_n642), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n616), .A2(new_n614), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n635), .B1(new_n437), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n648), .B(KEYINPUT94), .ZN(G369));
  INV_X1    g0449(.A(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(G20), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n209), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n505), .B1(new_n498), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n504), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n640), .A2(new_n658), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n577), .A2(new_n658), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n640), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n587), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n640), .A2(new_n504), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n493), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n658), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT95), .Z(G399));
  INV_X1    g0473(.A(new_n213), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n593), .A2(new_n216), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT96), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n675), .A2(new_n677), .A3(new_n209), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n235), .B2(new_n675), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT28), .Z(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n533), .A2(new_n534), .A3(new_n466), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n583), .A2(G179), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n612), .B(new_n471), .C1(new_n484), .C2(new_n485), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(G179), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n535), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n499), .A2(new_n500), .B1(new_n270), .B2(new_n470), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n688), .A4(new_n612), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n682), .A2(G179), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n486), .A3(new_n570), .A4(new_n610), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n685), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT97), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT97), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n692), .A2(new_n695), .A3(KEYINPUT31), .A4(new_n657), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT31), .B1(new_n618), .B2(new_n657), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n685), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(KEYINPUT98), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n700), .A2(new_n689), .A3(new_n691), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n657), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n697), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G330), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT99), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT99), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n587), .A2(new_n493), .A3(new_n504), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(new_n541), .A3(new_n617), .A4(new_n658), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n709), .A2(KEYINPUT31), .B1(new_n657), .B2(new_n702), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n707), .B(G330), .C1(new_n710), .C2(new_n697), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT29), .B1(new_n647), .B2(new_n657), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n647), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n680), .B1(new_n716), .B2(G1), .ZN(G364));
  OR2_X1    g0517(.A1(new_n666), .A2(G330), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT100), .Z(new_n719));
  NAND2_X1  g0519(.A1(new_n651), .A2(G45), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT101), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(G1), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n675), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n719), .A2(new_n667), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n210), .A2(new_n407), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT104), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT104), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n210), .B2(new_n407), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G190), .A2(G200), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G77), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n274), .A2(G179), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n210), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n274), .A2(G200), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n728), .A2(new_n730), .A3(new_n739), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n265), .B1(new_n326), .B2(new_n738), .C1(new_n740), .C2(new_n201), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n727), .A2(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G190), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(G68), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n210), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n745), .A2(new_n225), .B1(new_n747), .B2(new_n221), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n746), .A2(new_n274), .A3(G200), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n748), .B1(new_n753), .B2(G107), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n746), .A2(new_n731), .ZN(new_n755));
  INV_X1    g0555(.A(G159), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT32), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n736), .A2(new_n744), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G317), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(KEYINPUT33), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n743), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n763), .B1(new_n764), .B2(new_n740), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n735), .A2(G311), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n747), .B(KEYINPUT107), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n738), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n769), .A2(G303), .B1(G294), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n755), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(G329), .ZN(new_n773));
  INV_X1    g0573(.A(new_n745), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n265), .B(new_n773), .C1(G326), .C2(new_n774), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n766), .A2(new_n767), .A3(new_n771), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n752), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n759), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n233), .B1(G20), .B2(new_n304), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n781), .A2(KEYINPUT103), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(KEYINPUT103), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n236), .A2(new_n472), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n674), .A2(new_n265), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(new_n248), .C2(new_n472), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n213), .A2(new_n265), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT102), .Z(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G355), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n788), .B(new_n791), .C1(G116), .C2(new_n213), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n725), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n795), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n785), .B(new_n797), .C1(new_n666), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n726), .A2(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n423), .A2(new_n657), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n626), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n431), .A2(new_n433), .B1(new_n423), .B2(new_n657), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n712), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n706), .B2(new_n711), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n805), .A2(new_n807), .B1(new_n647), .B2(new_n657), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n706), .A2(new_n711), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n806), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n647), .A2(new_n657), .ZN(new_n811));
  INV_X1    g0611(.A(new_n807), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n808), .A2(new_n813), .A3(new_n725), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n735), .A2(G159), .B1(G150), .B2(new_n743), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  INV_X1    g0616(.A(G143), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(new_n745), .C1(new_n817), .C2(new_n740), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n753), .A2(G68), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n354), .B1(new_n772), .B2(G132), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(new_n201), .C2(new_n738), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n769), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  INV_X1    g0625(.A(new_n735), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n354), .B1(new_n825), .B2(new_n745), .C1(new_n826), .C2(new_n216), .ZN(new_n827));
  INV_X1    g0627(.A(G311), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n752), .A2(new_n221), .B1(new_n828), .B2(new_n755), .ZN(new_n829));
  INV_X1    g0629(.A(new_n743), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n830), .A2(new_n777), .B1(new_n326), .B2(new_n738), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n827), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n453), .B2(new_n768), .C1(new_n468), .C2(new_n740), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n824), .A2(new_n833), .B1(new_n782), .B2(new_n783), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n784), .A2(new_n793), .ZN(new_n835));
  AOI211_X1 g0635(.A(new_n725), .B(new_n834), .C1(new_n227), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n794), .B2(new_n804), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n814), .A2(new_n837), .ZN(G384));
  INV_X1    g0638(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n655), .B1(new_n411), .B2(new_n413), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n622), .B1(new_n403), .B2(new_n401), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT37), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT113), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n411), .A2(new_n413), .ZN(new_n845));
  INV_X1    g0645(.A(new_n655), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n845), .B1(new_n621), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT37), .B1(new_n405), .B2(new_n402), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(KEYINPUT113), .B(KEYINPUT37), .C1(new_n840), .C2(new_n841), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n840), .B1(new_n623), .B2(new_n633), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n366), .A2(new_n291), .A3(new_n374), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n400), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT112), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n400), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n846), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n416), .B2(new_n418), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n621), .A3(new_n858), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n403), .B2(new_n401), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT37), .B1(new_n863), .B2(new_n860), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n849), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n861), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n839), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n625), .A2(new_n657), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(new_n865), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n861), .A2(new_n865), .A3(KEYINPUT38), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n867), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n625), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n321), .A2(new_n657), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n875), .A2(new_n657), .B1(new_n348), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n804), .B(new_n658), .C1(new_n643), .C2(new_n646), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n433), .A2(new_n657), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n880), .A2(KEYINPUT111), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(KEYINPUT111), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n861), .B2(new_n865), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n878), .B(new_n885), .C1(new_n866), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n623), .A2(new_n655), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n874), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n436), .B1(new_n714), .B2(new_n715), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n635), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n889), .B(new_n891), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n698), .B2(new_n703), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n877), .A2(new_n894), .A3(new_n806), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n866), .B2(new_n886), .ZN(new_n896));
  NAND2_X1  g0696(.A1(KEYINPUT114), .A2(KEYINPUT40), .ZN(new_n897));
  OR2_X1    g0697(.A1(KEYINPUT114), .A2(KEYINPUT40), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT40), .B(new_n895), .C1(new_n853), .C2(new_n866), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n437), .A2(new_n894), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(G330), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n892), .B(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n209), .B2(new_n651), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n216), .B1(new_n517), .B2(KEYINPUT35), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n907), .B(new_n234), .C1(KEYINPUT35), .C2(new_n517), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT36), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n235), .A2(G77), .A3(new_n359), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n910), .B(KEYINPUT109), .Z(new_n911));
  NOR2_X1   g0711(.A1(new_n202), .A2(G50), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT110), .ZN(new_n913));
  OAI211_X1 g0713(.A(G1), .B(new_n650), .C1(new_n911), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n906), .A2(new_n909), .A3(new_n914), .ZN(G367));
  NAND2_X1  g0715(.A1(new_n523), .A2(new_n657), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n541), .A2(new_n504), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n657), .B1(new_n917), .B2(new_n642), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n639), .A2(new_n642), .A3(new_n916), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n540), .A2(new_n523), .A3(new_n657), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n662), .A2(new_n505), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OR2_X1    g0724(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(KEYINPUT42), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n918), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n658), .B1(new_n596), .B2(new_n597), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n616), .A2(new_n928), .A3(new_n614), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT115), .ZN(new_n930));
  INV_X1    g0730(.A(new_n617), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n928), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n930), .B2(new_n929), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n934), .B2(new_n933), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n927), .A2(KEYINPUT116), .A3(new_n936), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT116), .B1(new_n927), .B2(new_n936), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n668), .A2(new_n922), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n675), .B(KEYINPUT41), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT117), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n647), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n809), .A2(new_n713), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n663), .A2(new_n667), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n668), .A2(new_n923), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n946), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n950), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n716), .A2(KEYINPUT117), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n671), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n919), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT44), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT45), .ZN(new_n958));
  NOR3_X1   g0758(.A1(new_n954), .A2(new_n958), .A3(new_n922), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT45), .B1(new_n671), .B2(new_n921), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n956), .B(new_n957), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n668), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n951), .A2(new_n953), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n945), .B1(new_n963), .B2(new_n716), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n943), .B1(new_n964), .B2(new_n723), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n752), .A2(new_n326), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n735), .B2(G283), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n830), .A2(new_n468), .B1(new_n453), .B2(new_n738), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT46), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n747), .B2(new_n216), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n740), .B2(new_n825), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n969), .A2(new_n265), .A3(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n967), .A2(new_n968), .A3(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n828), .B2(new_n745), .C1(new_n760), .C2(new_n755), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n354), .B1(new_n735), .B2(G50), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n227), .B2(new_n752), .C1(new_n817), .C2(new_n745), .ZN(new_n977));
  INV_X1    g0777(.A(new_n740), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(G150), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n743), .A2(G159), .B1(G137), .B2(new_n772), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n202), .C2(new_n738), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n747), .A2(new_n201), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n784), .ZN(new_n985));
  INV_X1    g0785(.A(new_n787), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n796), .B1(new_n213), .B2(new_n595), .C1(new_n244), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n724), .A3(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT118), .Z(new_n989));
  NAND2_X1  g0789(.A1(new_n933), .A2(new_n795), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n965), .A2(new_n991), .ZN(G387));
  NAND2_X1  g0792(.A1(new_n951), .A2(new_n953), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n675), .C1(new_n716), .C2(new_n952), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n354), .B1(new_n978), .B2(G50), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n227), .B2(new_n747), .C1(new_n756), .C2(new_n745), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n395), .B2(new_n743), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n770), .A2(new_n419), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n772), .A2(G150), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n966), .B1(new_n735), .B2(G68), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n735), .A2(G303), .B1(G311), .B2(new_n743), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n760), .B2(new_n740), .C1(new_n764), .C2(new_n745), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT48), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n777), .B2(new_n738), .C1(new_n468), .C2(new_n747), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT49), .Z(new_n1006));
  AOI21_X1  g0806(.A(new_n265), .B1(new_n772), .B2(G326), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n752), .B2(new_n216), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n784), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n284), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n225), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n202), .A2(new_n227), .ZN(new_n1014));
  NOR4_X1   g0814(.A1(new_n1013), .A2(G45), .A3(new_n1014), .A4(new_n677), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n787), .B1(new_n241), .B2(new_n472), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n790), .A2(new_n677), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n213), .A2(G107), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n796), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n659), .A2(new_n660), .A3(new_n795), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1010), .A2(new_n724), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n723), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n994), .B(new_n1022), .C1(new_n1023), .C2(new_n950), .ZN(G393));
  AND3_X1   g0824(.A1(new_n951), .A2(new_n953), .A3(new_n962), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n962), .B1(new_n951), .B2(new_n953), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n675), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n962), .A2(new_n723), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n796), .B1(new_n251), .B2(new_n986), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G97), .B2(new_n674), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n752), .A2(new_n221), .B1(new_n202), .B2(new_n747), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n354), .B(new_n1032), .C1(G143), .C2(new_n772), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n770), .A2(G77), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n735), .A2(new_n1011), .B1(G50), .B2(new_n743), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n740), .A2(new_n756), .B1(new_n277), .B2(new_n745), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT51), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n740), .A2(new_n828), .B1(new_n760), .B2(new_n745), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1039), .B(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n265), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n772), .A2(G322), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n747), .A2(new_n777), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n735), .B2(G294), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n753), .A2(G107), .B1(G116), .B2(new_n770), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1042), .A2(new_n1043), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n830), .A2(new_n825), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1038), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n725), .B(new_n1031), .C1(new_n1049), .C2(new_n784), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n921), .B2(new_n798), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1029), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(KEYINPUT120), .B1(new_n1028), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1026), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n675), .A3(new_n963), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT120), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1055), .A2(new_n1056), .A3(new_n1029), .A4(new_n1051), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1053), .A2(new_n1057), .ZN(G390));
  NAND2_X1  g0858(.A1(new_n867), .A2(new_n873), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n820), .B1(new_n453), .B2(new_n830), .C1(new_n777), .C2(new_n745), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1034), .B1(new_n768), .B2(new_n221), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n354), .B1(new_n755), .B2(new_n468), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(new_n326), .B2(new_n826), .C1(new_n216), .C2(new_n740), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n826), .A2(new_n1065), .B1(new_n816), .B2(new_n830), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT122), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n747), .A2(new_n277), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT53), .ZN(new_n1070));
  INV_X1    g0870(.A(G132), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(new_n225), .B2(new_n752), .C1(new_n1071), .C2(new_n740), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n265), .B1(new_n738), .B2(new_n756), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G125), .B2(new_n772), .ZN(new_n1075));
  INV_X1    g0875(.A(G128), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1073), .B(new_n1075), .C1(new_n1076), .C2(new_n745), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1064), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1059), .A2(new_n793), .B1(new_n784), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n725), .B1(new_n835), .B2(new_n286), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT121), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n879), .A2(new_n882), .A3(new_n884), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1083), .A2(new_n877), .B1(new_n625), .B2(new_n657), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1059), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n807), .A2(new_n878), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n868), .B1(new_n885), .B2(new_n878), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n866), .B2(new_n853), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n895), .A2(G330), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1087), .B1(new_n867), .B2(new_n873), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n853), .A2(new_n866), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n1023), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n894), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n350), .A2(new_n1098), .A3(G330), .A4(new_n435), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n890), .A2(new_n635), .A3(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1090), .B1(new_n807), .B2(new_n878), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n885), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1098), .A2(G330), .A3(new_n804), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n877), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1086), .A2(new_n1083), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1100), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1027), .B1(new_n1096), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1089), .A2(new_n1106), .A3(new_n1095), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1082), .B(new_n1097), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(G378));
  NAND3_X1  g0911(.A1(new_n899), .A2(G330), .A3(new_n900), .ZN(new_n1112));
  XOR2_X1   g0912(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1113));
  XNOR2_X1  g0913(.A(new_n308), .B(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n298), .A2(new_n846), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1116), .A2(new_n899), .A3(G330), .A4(new_n900), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1118), .A2(new_n889), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n889), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n738), .A2(new_n202), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n735), .A2(new_n419), .B1(G283), .B2(new_n772), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n201), .B2(new_n752), .C1(new_n326), .C2(new_n830), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(G107), .C2(new_n978), .ZN(new_n1126));
  AOI211_X1 g0926(.A(G41), .B(new_n265), .C1(new_n774), .C2(G116), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1126), .B(new_n1127), .C1(new_n227), .C2(new_n747), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT58), .Z(new_n1129));
  NOR2_X1   g0929(.A1(new_n738), .A2(new_n277), .ZN(new_n1130));
  INV_X1    g0930(.A(G125), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n740), .A2(new_n1076), .B1(new_n1131), .B2(new_n745), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1130), .B(new_n1132), .C1(new_n735), .C2(G137), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n1071), .B2(new_n830), .C1(new_n747), .C2(new_n1065), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n1135));
  XNOR2_X1  g0935(.A(new_n1134), .B(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n772), .A2(G124), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G33), .B(G41), .C1(new_n753), .C2(G159), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n225), .B1(new_n352), .B2(G41), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n784), .B1(new_n1129), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT124), .Z(new_n1143));
  INV_X1    g0943(.A(new_n835), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n724), .B1(new_n1144), .B2(G50), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1116), .A2(new_n793), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT125), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT125), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1122), .A2(new_n723), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1100), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1109), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n889), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1118), .A2(new_n889), .A3(new_n1119), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1153), .A2(KEYINPUT57), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n675), .ZN(new_n1159));
  AOI21_X1  g0959(.A(KEYINPUT57), .B1(new_n1122), .B2(new_n1153), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1151), .B1(new_n1159), .B2(new_n1160), .ZN(G375));
  AOI21_X1  g0961(.A(new_n265), .B1(new_n735), .B2(G107), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n753), .A2(G77), .B1(G294), .B2(new_n774), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n216), .C2(new_n830), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n768), .A2(new_n326), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n740), .A2(new_n777), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n998), .B1(new_n825), .B2(new_n755), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n354), .B1(new_n735), .B2(G150), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n753), .A2(G58), .B1(G132), .B2(new_n774), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(new_n225), .C2(new_n738), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n768), .A2(new_n756), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n830), .A2(new_n1065), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n740), .A2(new_n816), .B1(new_n1076), .B2(new_n755), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n784), .B1(new_n1168), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1176), .B(new_n724), .C1(G68), .C2(new_n1144), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n877), .B2(new_n793), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n723), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1102), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n944), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1182), .B2(new_n1106), .ZN(G381));
  OR2_X1    g0983(.A1(G375), .A2(G378), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1184), .A2(G384), .A3(G381), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1053), .A2(new_n1057), .A3(new_n965), .A4(new_n991), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n1186), .A2(G396), .A3(G393), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(G407));
  OAI211_X1 g0988(.A(G407), .B(G213), .C1(G343), .C2(new_n1184), .ZN(G409));
  NAND2_X1  g0989(.A1(G375), .A2(G378), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n656), .A2(G213), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1122), .A2(new_n944), .A3(new_n1153), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1110), .A2(new_n1151), .A3(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(G384), .B(KEYINPUT126), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1027), .B1(new_n1181), .B2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1107), .C1(new_n1196), .C2(new_n1181), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1180), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1195), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G384), .A2(KEYINPUT126), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1180), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(KEYINPUT62), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n656), .A2(G213), .A3(G2897), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1207), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT61), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G375), .A2(G378), .B1(G213), .B2(new_n656), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT62), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1193), .A4(new_n1203), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1205), .A2(new_n1212), .A3(new_n1213), .A4(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(G396), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(G390), .A2(G387), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1053), .A2(new_n1057), .B1(new_n965), .B2(new_n991), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  XOR2_X1   g1021(.A(G393), .B(G396), .Z(new_n1222));
  NAND2_X1  g1022(.A1(G390), .A2(G387), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(new_n1223), .A3(new_n1186), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1217), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1225), .A2(KEYINPUT61), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1214), .A2(KEYINPUT63), .A3(new_n1193), .A4(new_n1203), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1206), .B2(new_n1211), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1204), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1227), .B(new_n1228), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1232), .ZN(G405));
  NAND2_X1  g1033(.A1(new_n1184), .A2(new_n1190), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1225), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1203), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1237), .A2(new_n1184), .A3(new_n1190), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(G402));
endmodule


