

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U546 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U547 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  NOR2_X2 U548 ( .A1(G164), .A2(G1384), .ZN(n603) );
  AND2_X1 U549 ( .A1(n712), .A2(n513), .ZN(n511) );
  AND2_X1 U550 ( .A1(n681), .A2(n701), .ZN(n512) );
  OR2_X1 U551 ( .A1(n711), .A2(n710), .ZN(n513) );
  INV_X1 U552 ( .A(KEYINPUT29), .ZN(n649) );
  XNOR2_X1 U553 ( .A(n650), .B(n649), .ZN(n656) );
  AND2_X1 U554 ( .A1(n512), .A2(n686), .ZN(n685) );
  AND2_X1 U555 ( .A1(n713), .A2(n511), .ZN(n714) );
  NOR2_X1 U556 ( .A1(G651), .A2(n570), .ZN(n797) );
  AND2_X1 U557 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X2 U558 ( .A(n514), .B(KEYINPUT17), .ZN(n882) );
  NAND2_X1 U559 ( .A1(n882), .A2(G138), .ZN(n515) );
  XNOR2_X1 U560 ( .A(n515), .B(KEYINPUT92), .ZN(n522) );
  INV_X1 U561 ( .A(G2105), .ZN(n518) );
  AND2_X1 U562 ( .A1(n518), .A2(G2104), .ZN(n881) );
  NAND2_X1 U563 ( .A1(G102), .A2(n881), .ZN(n517) );
  AND2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U565 ( .A1(G114), .A2(n885), .ZN(n516) );
  AND2_X1 U566 ( .A1(n517), .A2(n516), .ZN(n520) );
  NOR2_X1 U567 ( .A1(G2104), .A2(n518), .ZN(n887) );
  NAND2_X1 U568 ( .A1(G126), .A2(n887), .ZN(n519) );
  AND2_X1 U569 ( .A1(n520), .A2(n519), .ZN(n521) );
  INV_X1 U570 ( .A(KEYINPUT93), .ZN(n523) );
  XNOR2_X1 U571 ( .A(n524), .B(n523), .ZN(G164) );
  NAND2_X1 U572 ( .A1(n882), .A2(G137), .ZN(n527) );
  NAND2_X1 U573 ( .A1(G101), .A2(n881), .ZN(n525) );
  XOR2_X1 U574 ( .A(KEYINPUT23), .B(n525), .Z(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G113), .A2(n885), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G125), .A2(n887), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(G160) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n570) );
  INV_X1 U581 ( .A(G651), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n570), .A2(n532), .ZN(n794) );
  NAND2_X1 U583 ( .A1(G75), .A2(n794), .ZN(n536) );
  NOR2_X1 U584 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n533), .Z(n534) );
  XNOR2_X1 U586 ( .A(KEYINPUT66), .B(n534), .ZN(n798) );
  NAND2_X1 U587 ( .A1(G62), .A2(n798), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n539) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U590 ( .A1(n793), .A2(G88), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT86), .B(n537), .Z(n538) );
  NOR2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n797), .A2(G50), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(G303) );
  NAND2_X1 U595 ( .A1(n797), .A2(G51), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G63), .A2(n798), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U598 ( .A(KEYINPUT6), .B(n544), .ZN(n551) );
  NAND2_X1 U599 ( .A1(G89), .A2(n793), .ZN(n545) );
  XNOR2_X1 U600 ( .A(n545), .B(KEYINPUT4), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n546), .B(KEYINPUT76), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G76), .A2(n794), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U604 ( .A(n549), .B(KEYINPUT5), .Z(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U606 ( .A(KEYINPUT77), .B(n552), .Z(n553) );
  XOR2_X1 U607 ( .A(KEYINPUT7), .B(n553), .Z(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(n797), .A2(G53), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G65), .A2(n798), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U612 ( .A(KEYINPUT70), .B(n556), .Z(n560) );
  NAND2_X1 U613 ( .A1(G91), .A2(n793), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G78), .A2(n794), .ZN(n557) );
  AND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(G299) );
  NAND2_X1 U617 ( .A1(n797), .A2(G52), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G64), .A2(n798), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n569) );
  NAND2_X1 U620 ( .A1(n794), .A2(G77), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT69), .B(n563), .ZN(n566) );
  NAND2_X1 U622 ( .A1(n793), .A2(G90), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT68), .B(n564), .Z(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U625 ( .A(n567), .B(KEYINPUT9), .ZN(n568) );
  NOR2_X1 U626 ( .A1(n569), .A2(n568), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G87), .A2(n570), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n798), .A2(n573), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n797), .A2(G49), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n575), .A2(n574), .ZN(G288) );
  NAND2_X1 U633 ( .A1(G86), .A2(n793), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G61), .A2(n798), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U636 ( .A(KEYINPUT84), .B(n578), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G73), .A2(n794), .ZN(n579) );
  XNOR2_X1 U638 ( .A(n579), .B(KEYINPUT85), .ZN(n580) );
  XNOR2_X1 U639 ( .A(n580), .B(KEYINPUT2), .ZN(n581) );
  NOR2_X1 U640 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n797), .A2(G48), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n584), .A2(n583), .ZN(G305) );
  INV_X1 U643 ( .A(G303), .ZN(G166) );
  NAND2_X1 U644 ( .A1(n798), .A2(G60), .ZN(n585) );
  XNOR2_X1 U645 ( .A(n585), .B(KEYINPUT67), .ZN(n590) );
  NAND2_X1 U646 ( .A1(G85), .A2(n793), .ZN(n587) );
  NAND2_X1 U647 ( .A1(G72), .A2(n794), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT65), .B(n588), .Z(n589) );
  NOR2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n797), .A2(G47), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n592), .A2(n591), .ZN(G290) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n602) );
  NOR2_X1 U654 ( .A1(n603), .A2(n602), .ZN(n749) );
  XOR2_X1 U655 ( .A(G2067), .B(KEYINPUT37), .Z(n746) );
  NAND2_X1 U656 ( .A1(G104), .A2(n881), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G140), .A2(n882), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U659 ( .A(KEYINPUT34), .B(n595), .ZN(n600) );
  NAND2_X1 U660 ( .A1(G116), .A2(n885), .ZN(n597) );
  NAND2_X1 U661 ( .A1(G128), .A2(n887), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(KEYINPUT35), .B(n598), .Z(n599) );
  NOR2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U665 ( .A(KEYINPUT36), .B(n601), .Z(n895) );
  AND2_X1 U666 ( .A1(n746), .A2(n895), .ZN(n918) );
  NAND2_X1 U667 ( .A1(n749), .A2(n918), .ZN(n743) );
  INV_X1 U668 ( .A(n743), .ZN(n715) );
  INV_X1 U669 ( .A(KEYINPUT64), .ZN(n606) );
  INV_X1 U670 ( .A(n602), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X2 U672 ( .A(n606), .B(n605), .ZN(n651) );
  INV_X1 U673 ( .A(n651), .ZN(n657) );
  NOR2_X1 U674 ( .A1(n657), .A2(G2090), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n657), .A2(G8), .ZN(n711) );
  NOR2_X1 U676 ( .A1(G1971), .A2(n711), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n609), .A2(G303), .ZN(n669) );
  NAND2_X1 U679 ( .A1(G2072), .A2(n651), .ZN(n610) );
  XNOR2_X1 U680 ( .A(KEYINPUT27), .B(n610), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n657), .A2(G1956), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT97), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U684 ( .A(n614), .B(KEYINPUT98), .ZN(n617) );
  INV_X1 U685 ( .A(G299), .ZN(n966) );
  NOR2_X1 U686 ( .A1(n617), .A2(n966), .ZN(n616) );
  XNOR2_X1 U687 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n648) );
  NAND2_X1 U689 ( .A1(n966), .A2(n617), .ZN(n646) );
  NAND2_X1 U690 ( .A1(n798), .A2(G56), .ZN(n618) );
  XOR2_X1 U691 ( .A(KEYINPUT14), .B(n618), .Z(n624) );
  NAND2_X1 U692 ( .A1(n793), .A2(G81), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G68), .A2(n794), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U696 ( .A(KEYINPUT13), .B(n622), .Z(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n797), .A2(G43), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n975) );
  NAND2_X1 U700 ( .A1(n651), .A2(G1996), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT26), .ZN(n629) );
  NAND2_X1 U702 ( .A1(n657), .A2(G1341), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U704 ( .A1(n975), .A2(n630), .ZN(n641) );
  NAND2_X1 U705 ( .A1(G79), .A2(n794), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G54), .A2(n797), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G92), .A2(n793), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G66), .A2(n798), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT15), .ZN(n965) );
  NAND2_X1 U713 ( .A1(G2067), .A2(n651), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n657), .A2(G1348), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n965), .A2(n642), .ZN(n640) );
  OR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n965), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n650) );
  XOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .Z(n943) );
  NAND2_X1 U723 ( .A1(n943), .A2(n651), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n657), .A2(G1961), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U726 ( .A(KEYINPUT96), .B(n654), .Z(n661) );
  NAND2_X1 U727 ( .A1(G171), .A2(n661), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n667) );
  INV_X1 U729 ( .A(KEYINPUT31), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n657), .A2(G2084), .ZN(n699) );
  NOR2_X1 U731 ( .A1(G1966), .A2(n711), .ZN(n673) );
  NOR2_X1 U732 ( .A1(n699), .A2(n673), .ZN(n658) );
  NAND2_X1 U733 ( .A1(G8), .A2(n658), .ZN(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT30), .B(n659), .ZN(n660) );
  NOR2_X1 U735 ( .A1(G168), .A2(n660), .ZN(n663) );
  NOR2_X1 U736 ( .A1(G171), .A2(n661), .ZN(n662) );
  NOR2_X1 U737 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n677) );
  NAND2_X1 U740 ( .A1(G286), .A2(n677), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U742 ( .A1(G8), .A2(n670), .ZN(n672) );
  XOR2_X1 U743 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n671) );
  XNOR2_X1 U744 ( .A(n672), .B(n671), .ZN(n704) );
  INV_X1 U745 ( .A(n673), .ZN(n678) );
  AND2_X1 U746 ( .A1(n678), .A2(KEYINPUT100), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n677), .A2(n674), .ZN(n700) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n974) );
  INV_X1 U749 ( .A(n974), .ZN(n675) );
  OR2_X1 U750 ( .A1(n711), .A2(n675), .ZN(n689) );
  INV_X1 U751 ( .A(n689), .ZN(n676) );
  AND2_X1 U752 ( .A1(n700), .A2(n676), .ZN(n681) );
  INV_X1 U753 ( .A(KEYINPUT100), .ZN(n680) );
  NAND2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U755 ( .A1(n680), .A2(n679), .ZN(n701) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n688), .A2(KEYINPUT33), .ZN(n682) );
  NOR2_X1 U758 ( .A1(n682), .A2(n711), .ZN(n684) );
  XOR2_X1 U759 ( .A(G1981), .B(G305), .Z(n962) );
  INV_X1 U760 ( .A(n962), .ZN(n683) );
  NOR2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n704), .A2(n685), .ZN(n695) );
  INV_X1 U763 ( .A(n686), .ZN(n693) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U765 ( .A1(n688), .A2(n687), .ZN(n980) );
  OR2_X1 U766 ( .A1(n689), .A2(n980), .ZN(n691) );
  INV_X1 U767 ( .A(KEYINPUT33), .ZN(n690) );
  AND2_X1 U768 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U769 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U770 ( .A(n696), .B(KEYINPUT102), .ZN(n713) );
  NAND2_X1 U771 ( .A1(G8), .A2(G166), .ZN(n697) );
  NOR2_X1 U772 ( .A1(G2090), .A2(n697), .ZN(n698) );
  XNOR2_X1 U773 ( .A(n698), .B(KEYINPUT103), .ZN(n707) );
  NAND2_X1 U774 ( .A1(G8), .A2(n699), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n700), .A2(n701), .ZN(n702) );
  NAND2_X1 U776 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U779 ( .A1(n708), .A2(n711), .ZN(n712) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n709) );
  XOR2_X1 U781 ( .A(n709), .B(KEYINPUT24), .Z(n710) );
  NOR2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n881), .A2(G95), .ZN(n716) );
  XNOR2_X1 U784 ( .A(n716), .B(KEYINPUT94), .ZN(n718) );
  NAND2_X1 U785 ( .A1(G119), .A2(n887), .ZN(n717) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U787 ( .A1(G131), .A2(n882), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G107), .A2(n885), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U790 ( .A1(n722), .A2(n721), .ZN(n877) );
  INV_X1 U791 ( .A(G1991), .ZN(n940) );
  NOR2_X1 U792 ( .A1(n877), .A2(n940), .ZN(n732) );
  NAND2_X1 U793 ( .A1(G117), .A2(n885), .ZN(n724) );
  NAND2_X1 U794 ( .A1(G129), .A2(n887), .ZN(n723) );
  NAND2_X1 U795 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U796 ( .A(n725), .B(KEYINPUT95), .ZN(n727) );
  NAND2_X1 U797 ( .A1(G141), .A2(n882), .ZN(n726) );
  NAND2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U799 ( .A1(n881), .A2(G105), .ZN(n728) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(n728), .Z(n729) );
  OR2_X1 U801 ( .A1(n730), .A2(n729), .ZN(n864) );
  AND2_X1 U802 ( .A1(n864), .A2(G1996), .ZN(n731) );
  NOR2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n739) );
  XOR2_X1 U804 ( .A(G1986), .B(G290), .Z(n977) );
  NAND2_X1 U805 ( .A1(n739), .A2(n977), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n733), .A2(n749), .ZN(n734) );
  NAND2_X1 U807 ( .A1(n735), .A2(n734), .ZN(n752) );
  NOR2_X1 U808 ( .A1(G1996), .A2(n864), .ZN(n736) );
  XNOR2_X1 U809 ( .A(KEYINPUT104), .B(n736), .ZN(n920) );
  AND2_X1 U810 ( .A1(n940), .A2(n877), .ZN(n923) );
  NOR2_X1 U811 ( .A1(G1986), .A2(G290), .ZN(n737) );
  XOR2_X1 U812 ( .A(n737), .B(KEYINPUT105), .Z(n738) );
  NOR2_X1 U813 ( .A1(n923), .A2(n738), .ZN(n740) );
  INV_X1 U814 ( .A(n739), .ZN(n917) );
  NOR2_X1 U815 ( .A1(n740), .A2(n917), .ZN(n741) );
  NOR2_X1 U816 ( .A1(n920), .A2(n741), .ZN(n742) );
  XNOR2_X1 U817 ( .A(n742), .B(KEYINPUT39), .ZN(n744) );
  NAND2_X1 U818 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U819 ( .A(n745), .B(KEYINPUT106), .ZN(n748) );
  NOR2_X1 U820 ( .A1(n895), .A2(n746), .ZN(n747) );
  XNOR2_X1 U821 ( .A(n747), .B(KEYINPUT107), .ZN(n933) );
  NAND2_X1 U822 ( .A1(n748), .A2(n933), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n754) );
  XNOR2_X1 U825 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n753) );
  XNOR2_X1 U826 ( .A(n754), .B(n753), .ZN(G329) );
  INV_X1 U827 ( .A(G171), .ZN(G301) );
  XOR2_X1 U828 ( .A(G2443), .B(G2446), .Z(n756) );
  XNOR2_X1 U829 ( .A(G2427), .B(G2451), .ZN(n755) );
  XNOR2_X1 U830 ( .A(n756), .B(n755), .ZN(n762) );
  XOR2_X1 U831 ( .A(G2430), .B(G2454), .Z(n758) );
  XNOR2_X1 U832 ( .A(G1341), .B(G1348), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n758), .B(n757), .ZN(n760) );
  XOR2_X1 U834 ( .A(G2435), .B(G2438), .Z(n759) );
  XNOR2_X1 U835 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U836 ( .A(n762), .B(n761), .Z(n763) );
  AND2_X1 U837 ( .A1(G14), .A2(n763), .ZN(G401) );
  AND2_X1 U838 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U839 ( .A1(G111), .A2(n885), .ZN(n772) );
  NAND2_X1 U840 ( .A1(G123), .A2(n887), .ZN(n764) );
  XNOR2_X1 U841 ( .A(n764), .B(KEYINPUT18), .ZN(n767) );
  NAND2_X1 U842 ( .A1(G135), .A2(n882), .ZN(n765) );
  XNOR2_X1 U843 ( .A(n765), .B(KEYINPUT80), .ZN(n766) );
  NAND2_X1 U844 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U845 ( .A1(G99), .A2(n881), .ZN(n768) );
  XNOR2_X1 U846 ( .A(KEYINPUT81), .B(n768), .ZN(n769) );
  NOR2_X1 U847 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U848 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U849 ( .A(n773), .B(KEYINPUT82), .ZN(n924) );
  XNOR2_X1 U850 ( .A(n924), .B(G2096), .ZN(n774) );
  OR2_X1 U851 ( .A1(G2100), .A2(n774), .ZN(G156) );
  INV_X1 U852 ( .A(G132), .ZN(G219) );
  NAND2_X1 U853 ( .A1(G7), .A2(G661), .ZN(n775) );
  XNOR2_X1 U854 ( .A(n775), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U855 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n777) );
  XNOR2_X1 U856 ( .A(G223), .B(KEYINPUT73), .ZN(n834) );
  NAND2_X1 U857 ( .A1(G567), .A2(n834), .ZN(n776) );
  XNOR2_X1 U858 ( .A(n777), .B(n776), .ZN(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n784) );
  OR2_X1 U860 ( .A1(n975), .A2(n784), .ZN(G153) );
  INV_X1 U861 ( .A(n965), .ZN(n791) );
  NOR2_X1 U862 ( .A1(n791), .A2(G868), .ZN(n778) );
  XNOR2_X1 U863 ( .A(n778), .B(KEYINPUT75), .ZN(n780) );
  NAND2_X1 U864 ( .A1(G868), .A2(G301), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(G284) );
  INV_X1 U866 ( .A(G868), .ZN(n814) );
  NOR2_X1 U867 ( .A1(G286), .A2(n814), .ZN(n782) );
  NOR2_X1 U868 ( .A1(G868), .A2(G299), .ZN(n781) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U870 ( .A(KEYINPUT78), .B(n783), .ZN(G297) );
  NAND2_X1 U871 ( .A1(n784), .A2(G559), .ZN(n785) );
  NAND2_X1 U872 ( .A1(n785), .A2(n791), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U874 ( .A1(G868), .A2(n975), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G868), .A2(n791), .ZN(n787) );
  NOR2_X1 U876 ( .A1(G559), .A2(n787), .ZN(n788) );
  NOR2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U878 ( .A(KEYINPUT79), .B(n790), .Z(G282) );
  NAND2_X1 U879 ( .A1(n791), .A2(G559), .ZN(n812) );
  XNOR2_X1 U880 ( .A(n975), .B(n812), .ZN(n792) );
  NOR2_X1 U881 ( .A1(n792), .A2(G860), .ZN(n804) );
  NAND2_X1 U882 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n803) );
  NAND2_X1 U885 ( .A1(n797), .A2(G55), .ZN(n800) );
  NAND2_X1 U886 ( .A1(G67), .A2(n798), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT83), .B(n801), .Z(n802) );
  OR2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n815) );
  XOR2_X1 U890 ( .A(n804), .B(n815), .Z(G145) );
  XOR2_X1 U891 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n805) );
  XNOR2_X1 U892 ( .A(G288), .B(n805), .ZN(n806) );
  XNOR2_X1 U893 ( .A(G305), .B(n806), .ZN(n808) );
  XNOR2_X1 U894 ( .A(n966), .B(G166), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U896 ( .A(n809), .B(n975), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(G290), .ZN(n811) );
  XOR2_X1 U898 ( .A(n815), .B(n811), .Z(n898) );
  XNOR2_X1 U899 ( .A(n812), .B(n898), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U903 ( .A1(G2084), .A2(G2078), .ZN(n819) );
  XOR2_X1 U904 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n818) );
  XNOR2_X1 U905 ( .A(n819), .B(n818), .ZN(n820) );
  NAND2_X1 U906 ( .A1(n820), .A2(G2090), .ZN(n821) );
  XOR2_X1 U907 ( .A(KEYINPUT89), .B(n821), .Z(n822) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U909 ( .A1(n823), .A2(G2072), .ZN(n824) );
  XNOR2_X1 U910 ( .A(KEYINPUT90), .B(n824), .ZN(G158) );
  XNOR2_X1 U911 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U912 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U913 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NAND2_X1 U914 ( .A1(G108), .A2(G120), .ZN(n825) );
  NOR2_X1 U915 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G69), .A2(n826), .ZN(n910) );
  NAND2_X1 U917 ( .A1(n910), .A2(G567), .ZN(n831) );
  NOR2_X1 U918 ( .A1(G220), .A2(G219), .ZN(n827) );
  XOR2_X1 U919 ( .A(KEYINPUT22), .B(n827), .Z(n828) );
  NOR2_X1 U920 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U921 ( .A1(G96), .A2(n829), .ZN(n909) );
  NAND2_X1 U922 ( .A1(n909), .A2(G2106), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n838) );
  NAND2_X1 U924 ( .A1(G661), .A2(G483), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT91), .B(n832), .Z(n833) );
  NOR2_X1 U926 ( .A1(n838), .A2(n833), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U933 ( .A(n838), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n840) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n842) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U941 ( .A(G2084), .B(G2078), .ZN(n845) );
  XNOR2_X1 U942 ( .A(n846), .B(n845), .ZN(G227) );
  XNOR2_X1 U943 ( .A(G1956), .B(KEYINPUT110), .ZN(n856) );
  XOR2_X1 U944 ( .A(G1976), .B(G1981), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1966), .B(G1961), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1986), .B(G1991), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1971), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2474), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G124), .A2(n887), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U956 ( .A1(n885), .A2(G112), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G100), .A2(n881), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G136), .A2(n882), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U961 ( .A1(n863), .A2(n862), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n866) );
  XOR2_X1 U963 ( .A(n864), .B(n924), .Z(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n876) );
  NAND2_X1 U965 ( .A1(G118), .A2(n885), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G130), .A2(n887), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U968 ( .A1(n881), .A2(G106), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT111), .B(n869), .Z(n871) );
  NAND2_X1 U970 ( .A1(n882), .A2(G142), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT45), .B(n872), .Z(n873) );
  NOR2_X1 U973 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(n876), .B(n875), .Z(n879) );
  XNOR2_X1 U975 ( .A(G164), .B(n877), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U977 ( .A(n880), .B(G162), .Z(n894) );
  NAND2_X1 U978 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n892) );
  NAND2_X1 U981 ( .A1(n885), .A2(G115), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n886), .B(KEYINPUT112), .ZN(n889) );
  NAND2_X1 U983 ( .A1(G127), .A2(n887), .ZN(n888) );
  NAND2_X1 U984 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n890), .Z(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n912) );
  XNOR2_X1 U987 ( .A(G160), .B(n912), .ZN(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U989 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U990 ( .A1(G37), .A2(n897), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n965), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U993 ( .A(G301), .B(n900), .Z(n901) );
  NOR2_X1 U994 ( .A1(G37), .A2(n901), .ZN(n902) );
  XOR2_X1 U995 ( .A(KEYINPUT113), .B(n902), .Z(G397) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n903) );
  XOR2_X1 U997 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U998 ( .A1(G319), .A2(n904), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G401), .A2(n905), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT114), .B(n906), .ZN(n908) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n908), .A2(n907), .ZN(G225) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(G120), .ZN(G236) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  INV_X1 U1007 ( .A(G96), .ZN(G221) );
  INV_X1 U1008 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n911), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U1011 ( .A(G261), .ZN(G325) );
  XOR2_X1 U1012 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n936) );
  XNOR2_X1 U1013 ( .A(G2072), .B(n912), .ZN(n915) );
  XOR2_X1 U1014 ( .A(G164), .B(G2078), .Z(n913) );
  XNOR2_X1 U1015 ( .A(KEYINPUT117), .B(n913), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT50), .ZN(n932) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n930) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT51), .B(n921), .ZN(n928) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(n926), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1031 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n959) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n959), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n938), .A2(G29), .ZN(n1018) );
  XNOR2_X1 U1034 ( .A(G2084), .B(G34), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT54), .ZN(n958) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n955) );
  XNOR2_X1 U1037 ( .A(n940), .B(G25), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(n941), .A2(G28), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(n942), .B(KEYINPUT120), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(n943), .B(G27), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G32), .B(G1996), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1043 ( .A(KEYINPUT121), .B(n946), .Z(n950) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n953), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT122), .B(n956), .Z(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(n959), .ZN(n961) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n961), .ZN(n1014) );
  XOR2_X1 U1055 ( .A(G16), .B(KEYINPUT56), .Z(n985) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(n964), .B(KEYINPUT57), .ZN(n972) );
  XOR2_X1 U1059 ( .A(n965), .B(G1348), .Z(n968) );
  XNOR2_X1 U1060 ( .A(n966), .B(G1956), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G1961), .B(G301), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n983) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n979) );
  XOR2_X1 U1067 ( .A(G1341), .B(n975), .Z(n976) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1072 ( .A1(n985), .A2(n984), .ZN(n1011) );
  XOR2_X1 U1073 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n1008) );
  XNOR2_X1 U1074 ( .A(KEYINPUT59), .B(G1348), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(n986), .B(G4), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G1956), .B(G20), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G6), .B(G1981), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(KEYINPUT123), .B(n989), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT60), .B(n994), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(G1976), .B(G23), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1986), .B(G24), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1087 ( .A(G1971), .B(KEYINPUT124), .Z(n997) );
  XNOR2_X1 U1088 ( .A(G22), .B(n997), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT58), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(G16), .A2(n1009), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1099 ( .A(KEYINPUT126), .B(n1012), .Z(n1013) );
  NOR2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(G11), .A2(n1015), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1019), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

