//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1311, new_n1312, new_n1313, new_n1314, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n201), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n207), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n212), .B1(KEYINPUT1), .B2(new_n223), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G68), .B(G77), .Z(new_n238));
  XOR2_X1   g0038(.A(G50), .B(G58), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n245), .B1(new_n202), .B2(KEYINPUT8), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT8), .B(G58), .ZN(new_n247));
  OAI21_X1  g0047(.A(new_n246), .B1(new_n247), .B2(new_n245), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT65), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n250), .B(new_n246), .C1(new_n247), .C2(new_n245), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n257), .B1(G150), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n255), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n224), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n206), .B2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G50), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n253), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n273), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n277), .A2(G223), .B1(new_n280), .B2(G77), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G222), .A3(new_n273), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n214), .ZN(new_n291));
  INV_X1    g0091(.A(G41), .ZN(new_n292));
  INV_X1    g0092(.A(G45), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n294), .A2(new_n286), .A3(G274), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT68), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n297), .A2(G200), .B1(new_n298), .B2(KEYINPUT10), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n288), .A2(G190), .A3(new_n296), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n271), .A2(new_n272), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n303), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n271), .A2(new_n305), .A3(new_n301), .A4(new_n272), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n297), .A2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n297), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n269), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT14), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n219), .A2(G1698), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(G226), .B2(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n319), .B2(new_n280), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n295), .B1(new_n320), .B2(new_n287), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n290), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n289), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(G238), .A3(new_n325), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n322), .B1(new_n321), .B2(new_n326), .ZN(new_n328));
  OAI211_X1 g0128(.A(G169), .B(new_n316), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n294), .A2(new_n286), .A3(G274), .ZN(new_n330));
  NOR2_X1   g0130(.A1(G226), .A2(G1698), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n219), .B2(G1698), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n282), .B1(G33), .B2(G97), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n330), .B1(new_n333), .B2(new_n286), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n324), .A2(G238), .A3(new_n325), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT13), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n321), .A2(new_n322), .A3(new_n326), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G179), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(new_n337), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n316), .B1(new_n340), .B2(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT71), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n315), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT71), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(new_n338), .A4(new_n329), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n254), .A2(G77), .B1(G20), .B2(new_n215), .ZN(new_n348));
  INV_X1    g0148(.A(new_n259), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n201), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n263), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n351), .B(KEYINPUT11), .Z(new_n352));
  INV_X1    g0152(.A(KEYINPUT67), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n265), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n206), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n267), .A2(G68), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n265), .A2(G68), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n357), .B(new_n359), .C1(KEYINPUT12), .C2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n347), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n336), .A2(G190), .A3(new_n337), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n340), .A2(G200), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G244), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n330), .B1(new_n368), .B2(new_n290), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n216), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G232), .B2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n282), .ZN(new_n372));
  INV_X1    g0172(.A(G107), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n286), .B1(new_n280), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n369), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G190), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n375), .ZN(new_n378));
  XOR2_X1   g0178(.A(KEYINPUT15), .B(G87), .Z(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n349), .B2(new_n247), .ZN(new_n381));
  INV_X1    g0181(.A(G77), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n381), .A2(new_n263), .B1(new_n382), .B2(new_n358), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n267), .A2(G77), .A3(new_n356), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n385), .B(new_n388), .C1(G169), .C2(new_n375), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n313), .A2(new_n364), .A3(new_n367), .A4(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n267), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n252), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n265), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n393), .B1(new_n394), .B2(new_n252), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT72), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n275), .A2(new_n207), .A3(new_n276), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n276), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT72), .B1(new_n397), .B2(new_n398), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n202), .A2(new_n215), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G58), .A2(G68), .ZN(new_n405));
  OAI21_X1  g0205(.A(G20), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n259), .A2(G159), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT16), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n280), .B2(new_n207), .ZN(new_n411));
  INV_X1    g0211(.A(new_n400), .ZN(new_n412));
  OAI21_X1  g0212(.A(G68), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n263), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n395), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT75), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT73), .ZN(new_n418));
  NOR2_X1   g0218(.A1(G223), .A2(G1698), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n214), .B2(G1698), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n282), .B1(G33), .B2(G87), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n421), .B2(new_n286), .ZN(new_n422));
  OR2_X1    g0222(.A1(G223), .A2(G1698), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n214), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n423), .B(new_n424), .C1(new_n278), .C2(new_n279), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n286), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT73), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n286), .A2(G232), .A3(new_n289), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n330), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT74), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n330), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n432), .A2(new_n387), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n330), .A2(new_n430), .A3(new_n433), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n433), .B1(new_n330), .B2(new_n430), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n427), .ZN(new_n440));
  AOI21_X1  g0240(.A(G169), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n417), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n432), .A3(new_n434), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n309), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(KEYINPUT75), .C1(new_n429), .C2(new_n435), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n416), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT18), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n416), .A2(new_n442), .A3(new_n448), .A4(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(new_n429), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n437), .A2(new_n438), .A3(G190), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n453), .B1(new_n443), .B2(new_n377), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT76), .B1(new_n416), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n415), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT16), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT72), .B1(new_n411), .B2(new_n412), .ZN(new_n458));
  INV_X1    g0258(.A(new_n402), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n215), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n460), .B2(new_n408), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT76), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n443), .A2(new_n377), .ZN(new_n464));
  INV_X1    g0264(.A(G190), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n439), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n466), .B2(new_n429), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(new_n463), .A3(new_n395), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n451), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n416), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT17), .B1(new_n470), .B2(new_n467), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n450), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n391), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n356), .A2(new_n379), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT19), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(KEYINPUT81), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(G20), .B1(new_n275), .B2(new_n276), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n207), .B1(new_n317), .B2(new_n479), .ZN(new_n486));
  INV_X1    g0286(.A(G87), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(new_n220), .A3(new_n373), .ZN(new_n488));
  AOI22_X1  g0288(.A1(new_n485), .A2(G68), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n263), .ZN(new_n491));
  OAI211_X1 g0291(.A(KEYINPUT82), .B(new_n477), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n484), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n476), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n206), .A2(G33), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n491), .A2(new_n265), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n379), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT80), .B(G250), .C1(new_n293), .C2(G1), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT80), .ZN(new_n503));
  AOI21_X1  g0303(.A(G274), .B1(new_n503), .B2(G250), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n206), .A2(G45), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n286), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n253), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(G238), .A2(G1698), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n368), .B2(G1698), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n509), .B1(new_n511), .B2(new_n282), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n512), .B2(new_n286), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G169), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n507), .B(G179), .C1(new_n512), .C2(new_n286), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n492), .A2(new_n495), .B1(G87), .B2(new_n499), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT83), .B1(new_n513), .B2(new_n465), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n216), .A2(new_n273), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n368), .A2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(new_n278), .C2(new_n279), .ZN(new_n521));
  INV_X1    g0321(.A(new_n509), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n286), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n293), .A2(G1), .ZN(new_n524));
  INV_X1    g0324(.A(G250), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(KEYINPUT80), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n524), .B1(new_n526), .B2(G274), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n287), .B1(new_n527), .B2(new_n502), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(G190), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n518), .A2(new_n531), .B1(G200), .B2(new_n513), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n501), .A2(new_n516), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n349), .B2(new_n382), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n259), .A2(KEYINPUT77), .A3(G77), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n538), .A2(new_n220), .A3(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n537), .B1(new_n541), .B2(new_n207), .ZN(new_n542));
  OAI21_X1  g0342(.A(G107), .B1(new_n401), .B2(new_n402), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(KEYINPUT78), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT78), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(G107), .C1(new_n401), .C2(new_n402), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n263), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n265), .A2(G97), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n499), .B2(G97), .ZN(new_n550));
  OAI211_X1 g0350(.A(G250), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT79), .ZN(new_n552));
  OAI211_X1 g0352(.A(G244), .B(new_n273), .C1(new_n278), .C2(new_n279), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT4), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n287), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g0359(.A(KEYINPUT5), .B(G41), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(G274), .A3(new_n286), .A4(new_n524), .ZN(new_n561));
  AND2_X1   g0361(.A1(KEYINPUT5), .A2(G41), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT5), .A2(G41), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n524), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n286), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n221), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(new_n465), .A3(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n553), .A2(new_n554), .B1(G33), .B2(G283), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT79), .B1(new_n277), .B2(G250), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT79), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n551), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(new_n556), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n566), .B1(new_n573), .B2(new_n287), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n568), .B1(G200), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n548), .A2(new_n550), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n387), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n559), .A2(new_n567), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n309), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n491), .B1(new_n544), .B2(new_n546), .ZN(new_n580));
  INV_X1    g0380(.A(new_n550), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n577), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n533), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n358), .A2(new_n508), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n356), .A2(new_n491), .A3(G116), .A4(new_n497), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n262), .A2(new_n224), .B1(G20), .B2(new_n508), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(G33), .B2(G283), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n253), .A2(G97), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT85), .ZN(new_n590));
  AOI21_X1  g0390(.A(KEYINPUT85), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT20), .B(new_n587), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(G257), .B(new_n273), .C1(new_n278), .C2(new_n279), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(KEYINPUT84), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n277), .A2(G264), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT84), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n282), .A2(new_n600), .A3(G257), .A4(new_n273), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n280), .A2(G303), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n598), .A2(new_n599), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n287), .ZN(new_n604));
  INV_X1    g0404(.A(G270), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n561), .B1(new_n565), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  OR3_X1    g0408(.A1(new_n596), .A2(new_n608), .A3(new_n387), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n606), .B1(new_n603), .B2(new_n287), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G190), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n596), .C1(new_n377), .C2(new_n610), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n584), .A2(new_n585), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n594), .A2(new_n595), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n309), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT21), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n608), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n615), .B2(new_n608), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n609), .B(new_n612), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n564), .A2(G264), .A3(new_n286), .ZN(new_n621));
  NOR2_X1   g0421(.A1(G250), .A2(G1698), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n221), .B2(G1698), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n623), .A2(new_n282), .B1(G33), .B2(G294), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n561), .B(new_n621), .C1(new_n624), .C2(new_n286), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n309), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n221), .A2(G1698), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(G250), .B2(G1698), .ZN(new_n628));
  INV_X1    g0428(.A(G294), .ZN(new_n629));
  OAI22_X1  g0429(.A1(new_n628), .A2(new_n280), .B1(new_n253), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n287), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n387), .A3(new_n561), .A4(new_n621), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT23), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n207), .B2(G107), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n373), .A2(KEYINPUT23), .A3(G20), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n509), .B2(new_n207), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT22), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n485), .B2(G87), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n207), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT22), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT24), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n485), .A2(new_n638), .A3(G87), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(KEYINPUT22), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT24), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n637), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n491), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT25), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n265), .B2(G107), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n265), .A2(new_n650), .A3(G107), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n499), .A2(G107), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n633), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n649), .A2(new_n655), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n625), .A2(new_n465), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n625), .A2(G200), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n633), .B(KEYINPUT86), .C1(new_n649), .C2(new_n655), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NOR4_X1   g0464(.A1(new_n475), .A2(new_n583), .A3(new_n620), .A4(new_n664), .ZN(G372));
  NAND2_X1  g0465(.A1(new_n455), .A2(new_n468), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n471), .B1(new_n666), .B2(KEYINPUT17), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n362), .B1(new_n342), .B2(new_n346), .ZN(new_n668));
  INV_X1    g0468(.A(new_n367), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n389), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n667), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n447), .A2(new_n449), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT90), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n307), .B1(new_n673), .B2(KEYINPUT90), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n312), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n501), .A2(new_n516), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n529), .B2(new_n377), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n513), .A2(KEYINPUT87), .A3(G200), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n680), .A2(new_n681), .B1(new_n518), .B2(new_n531), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n517), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n677), .B1(new_n684), .B2(new_n582), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT88), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n517), .A2(new_n532), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g0489(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n690));
  OR3_X1    g0490(.A1(new_n689), .A2(new_n582), .A3(new_n690), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT88), .B(new_n677), .C1(new_n684), .C2(new_n582), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n678), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n501), .A2(new_n516), .B1(new_n517), .B2(new_n682), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n662), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n576), .A2(new_n582), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n615), .A2(new_n608), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT21), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n617), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(new_n609), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n656), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n694), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n676), .B1(new_n475), .B2(new_n706), .ZN(G369));
  NAND2_X1  g0507(.A1(new_n701), .A2(new_n609), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G213), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G343), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n596), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n620), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G330), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n659), .B2(new_n715), .ZN(new_n722));
  INV_X1    g0522(.A(new_n656), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n714), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n708), .A2(new_n715), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n664), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n656), .A2(new_n714), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(new_n210), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n488), .A2(G116), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n227), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n714), .B1(new_n693), .B2(new_n704), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n697), .A2(KEYINPUT93), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT93), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n576), .A2(new_n582), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n658), .A2(new_n663), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n696), .B1(new_n702), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n694), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n690), .B1(new_n689), .B2(new_n582), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(KEYINPUT92), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT92), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n751), .B(new_n690), .C1(new_n689), .C2(new_n582), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n579), .A2(new_n577), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n548), .B2(new_n550), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(new_n695), .A3(KEYINPUT26), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n750), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n714), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n740), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n741), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n621), .B1(new_n624), .B2(new_n286), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n515), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n761), .A2(new_n610), .A3(new_n559), .A4(new_n567), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT30), .ZN(new_n763));
  AND3_X1   g0563(.A1(new_n762), .A2(KEYINPUT91), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n763), .B1(new_n762), .B2(KEYINPUT91), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n625), .A2(new_n387), .A3(new_n513), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n574), .A2(new_n766), .A3(new_n610), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT31), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n768), .A2(new_n769), .A3(new_n715), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n762), .A2(KEYINPUT91), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n762), .A2(KEYINPUT91), .A3(new_n763), .ZN(new_n773));
  INV_X1    g0573(.A(new_n767), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(KEYINPUT31), .B1(new_n775), .B2(new_n714), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n664), .A2(new_n620), .ZN(new_n778));
  INV_X1    g0578(.A(new_n583), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n778), .A2(new_n779), .A3(new_n715), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G330), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n759), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n738), .B1(new_n784), .B2(G1), .ZN(G364));
  INV_X1    g0585(.A(G13), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n787), .B(KEYINPUT94), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G45), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G1), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n733), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n720), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G330), .B2(new_n718), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n732), .A2(new_n280), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G355), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G116), .B2(new_n210), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n732), .A2(new_n282), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n227), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(new_n293), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n240), .A2(G45), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n796), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n224), .B1(G20), .B2(new_n309), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n791), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G179), .A2(G200), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(G20), .B1(new_n811), .B2(new_n465), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT97), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT97), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n220), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n207), .A2(new_n465), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n377), .A2(G179), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n487), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n387), .A2(G200), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n821), .B1(G58), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n207), .A2(G190), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n819), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n825), .B1(new_n373), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n822), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n207), .A2(new_n387), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(new_n465), .A3(G200), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n282), .B1(new_n829), .B2(new_n382), .C1(new_n831), .C2(new_n215), .ZN(new_n832));
  NOR3_X1   g0632(.A1(new_n817), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n830), .A2(G190), .A3(G200), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(KEYINPUT95), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT95), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n201), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT96), .ZN(new_n839));
  INV_X1    g0639(.A(new_n826), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n811), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n826), .A2(KEYINPUT96), .A3(new_n810), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(G159), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT32), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n847), .A2(new_n827), .B1(new_n829), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G303), .ZN(new_n850));
  XOR2_X1   g0650(.A(KEYINPUT33), .B(G317), .Z(new_n851));
  OAI221_X1 g0651(.A(new_n280), .B1(new_n820), .B2(new_n850), .C1(new_n831), .C2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n849), .B(new_n852), .C1(G322), .C2(new_n824), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n844), .A2(G329), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n853), .B(new_n854), .C1(new_n629), .C2(new_n816), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n837), .B(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G326), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n838), .A2(new_n846), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT99), .ZN(new_n862));
  INV_X1    g0662(.A(new_n806), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n861), .B2(KEYINPUT99), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n809), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n805), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n718), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n793), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(G396));
  NOR2_X1   g0669(.A1(new_n389), .A2(new_n715), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(KEYINPUT101), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n385), .A2(new_n714), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n871), .A2(new_n872), .B1(new_n390), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n706), .B2(new_n714), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n390), .A2(new_n873), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n705), .A2(new_n715), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n791), .B1(new_n880), .B2(new_n782), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n782), .B2(new_n880), .ZN(new_n882));
  INV_X1    g0682(.A(new_n791), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n806), .A2(new_n803), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n382), .B2(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n823), .A2(new_n629), .B1(new_n829), .B2(new_n508), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n280), .B1(new_n827), .B2(new_n487), .C1(new_n831), .C2(new_n847), .ZN(new_n887));
  INV_X1    g0687(.A(new_n820), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n886), .B(new_n887), .C1(G107), .C2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n848), .B2(new_n843), .ZN(new_n890));
  INV_X1    g0690(.A(new_n837), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n817), .B(new_n890), .C1(G303), .C2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n829), .ZN(new_n893));
  AOI22_X1  g0693(.A1(G143), .A2(new_n824), .B1(new_n893), .B2(G159), .ZN(new_n894));
  INV_X1    g0694(.A(G150), .ZN(new_n895));
  INV_X1    g0695(.A(G137), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n894), .B1(new_n895), .B2(new_n831), .C1(new_n837), .C2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT34), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n280), .B1(new_n844), .B2(G132), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n900), .A2(KEYINPUT100), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(KEYINPUT100), .ZN(new_n902));
  INV_X1    g0702(.A(new_n827), .ZN(new_n903));
  AOI22_X1  g0703(.A1(G50), .A2(new_n888), .B1(new_n903), .B2(G68), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n816), .B2(new_n202), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n892), .B1(new_n898), .B2(new_n906), .ZN(new_n907));
  OAI221_X1 g0707(.A(new_n885), .B1(new_n907), .B2(new_n863), .C1(new_n878), .C2(new_n804), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n882), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(G384));
  NOR2_X1   g0710(.A1(new_n788), .A2(new_n206), .ZN(new_n911));
  INV_X1    g0711(.A(G330), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT38), .ZN(new_n913));
  INV_X1    g0713(.A(new_n712), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n416), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n667), .B2(new_n672), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT37), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n446), .A2(new_n917), .A3(new_n915), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n455), .A2(new_n468), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n446), .B(new_n915), .C1(new_n416), .C2(new_n454), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n918), .A2(new_n919), .B1(new_n920), .B2(KEYINPUT37), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n913), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n413), .A2(new_n409), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT16), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n413), .A2(KEYINPUT103), .A3(new_n409), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n415), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n249), .A2(new_n265), .A3(new_n251), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n393), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n442), .B(new_n445), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n914), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n931), .A2(new_n455), .A3(new_n468), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n923), .A2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(KEYINPUT38), .C1(new_n472), .C2(new_n932), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n922), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n874), .B1(new_n777), .B2(new_n780), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n362), .A2(new_n715), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n364), .A2(new_n367), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n939), .B1(new_n668), .B2(new_n669), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(KEYINPUT40), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT104), .B1(new_n937), .B2(new_n944), .ZN(new_n945));
  NOR4_X1   g0745(.A1(new_n583), .A2(new_n664), .A3(new_n620), .A4(new_n714), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n769), .B1(new_n768), .B2(new_n715), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n775), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n878), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n940), .B1(new_n364), .B2(new_n367), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n668), .A2(new_n669), .A3(new_n939), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n922), .A2(new_n936), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT104), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(KEYINPUT40), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n945), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n932), .B1(new_n667), .B2(new_n672), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n919), .A2(new_n918), .B1(new_n933), .B2(KEYINPUT37), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n913), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n936), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT40), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n958), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT105), .Z(new_n967));
  AND2_X1   g0767(.A1(new_n474), .A2(new_n781), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n912), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n389), .A2(new_n714), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n953), .B1(new_n879), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n962), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT39), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n955), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n364), .A2(new_n714), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n975), .C2(new_n962), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n450), .A2(new_n712), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n474), .B1(new_n741), .B2(new_n758), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n981), .A2(new_n676), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n980), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n911), .B1(new_n970), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n970), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT35), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n541), .A2(new_n986), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n508), .B(new_n226), .C1(new_n541), .C2(new_n986), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n987), .B1(new_n989), .B2(KEYINPUT102), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT102), .B2(new_n989), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT36), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n404), .A2(new_n227), .A3(new_n382), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n215), .A2(G50), .ZN(new_n994));
  OAI211_X1 g0794(.A(G1), .B(new_n786), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n985), .A2(new_n992), .A3(new_n995), .ZN(G367));
  INV_X1    g0796(.A(new_n379), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n807), .B1(new_n210), .B2(new_n997), .C1(new_n798), .C2(new_n236), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n791), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n282), .B1(new_n829), .B2(new_n201), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n903), .A2(G77), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n202), .B2(new_n820), .C1(new_n895), .C2(new_n823), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n831), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1000), .B(new_n1002), .C1(G159), .C2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n215), .B2(new_n816), .C1(new_n896), .C2(new_n843), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n857), .A2(G143), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n858), .A2(new_n848), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n280), .B1(new_n827), .B2(new_n220), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n823), .A2(new_n850), .B1(new_n829), .B2(new_n847), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n844), .C2(G317), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n888), .A2(G116), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT46), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1011), .A2(new_n1012), .B1(new_n831), .B2(new_n629), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1010), .B(new_n1014), .C1(new_n373), .C2(new_n816), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n999), .B1(new_n1017), .B2(new_n806), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n517), .A2(new_n715), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n678), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n695), .B2(new_n1019), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT106), .Z(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n805), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT108), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n727), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n725), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n728), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n722), .A2(KEYINPUT108), .A3(new_n724), .A4(new_n727), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(new_n720), .ZN(new_n1031));
  AND3_X1   g0831(.A1(new_n1031), .A2(new_n782), .A3(new_n759), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n714), .B1(new_n580), .B2(new_n581), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n745), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n754), .A2(new_n714), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n730), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT45), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1034), .B(new_n1035), .C1(new_n729), .C2(new_n728), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT44), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n726), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n726), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1032), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT109), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT109), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n1039), .A2(new_n726), .A3(new_n1042), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n726), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1052), .B2(new_n1032), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n784), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n733), .B(KEYINPUT41), .Z(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n790), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1036), .A2(new_n728), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1058), .A2(KEYINPUT42), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT107), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT43), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n582), .B1(new_n1034), .B2(new_n746), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1058), .A2(KEYINPUT42), .B1(new_n1065), .B2(new_n715), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1063), .A2(new_n1064), .A3(new_n1022), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n726), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1066), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1022), .A2(new_n1064), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1022), .A2(new_n1064), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1068), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1024), .B1(new_n1057), .B2(new_n1075), .ZN(G387));
  XOR2_X1   g0876(.A(new_n733), .B(KEYINPUT115), .Z(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1032), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n784), .B2(new_n1031), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1031), .A2(new_n790), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n735), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n794), .A2(new_n1082), .B1(new_n373), .B2(new_n732), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n233), .A2(new_n293), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n247), .A2(G50), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT50), .Z(new_n1086));
  OAI211_X1 g0886(.A(new_n735), .B(new_n293), .C1(new_n215), .C2(new_n382), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n797), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n883), .B1(new_n1089), .B2(new_n807), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n816), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n379), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n201), .A2(new_n823), .B1(new_n820), .B2(new_n382), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n280), .B(new_n1093), .C1(G97), .C2(new_n903), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(new_n895), .C2(new_n843), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n252), .A2(new_n1003), .B1(G68), .B2(new_n893), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT110), .Z(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G159), .C2(new_n891), .ZN(new_n1098));
  XOR2_X1   g0898(.A(KEYINPUT111), .B(G322), .Z(new_n1099));
  NAND2_X1  g0899(.A1(new_n857), .A2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n824), .B1(new_n893), .B2(G303), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n848), .C2(new_n831), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT112), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1103), .A2(KEYINPUT48), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(KEYINPUT48), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1091), .A2(G283), .B1(G294), .B2(new_n888), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT113), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(KEYINPUT113), .A3(new_n1106), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1104), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT49), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n280), .B1(new_n508), .B2(new_n827), .C1(new_n843), .C2(new_n859), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1111), .B2(KEYINPUT49), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1098), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1090), .B1(new_n1115), .B2(new_n863), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n725), .B2(new_n866), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1116), .A2(KEYINPUT114), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1080), .B(new_n1081), .C1(new_n1118), .C2(new_n1119), .ZN(G393));
  INV_X1    g0920(.A(new_n1032), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1046), .A2(new_n1043), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1078), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1034), .A2(new_n805), .A3(new_n1035), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n807), .B1(new_n220), .B2(new_n210), .C1(new_n798), .C2(new_n243), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n891), .A2(G317), .B1(G311), .B2(new_n824), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT52), .Z(new_n1128));
  NAND2_X1  g0928(.A1(new_n844), .A2(new_n1099), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1003), .A2(G303), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n282), .B1(new_n903), .B2(G107), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G283), .A2(new_n888), .B1(new_n893), .B2(G294), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n1091), .ZN(new_n1134));
  INV_X1    g0934(.A(G159), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n837), .A2(new_n895), .B1(new_n1135), .B2(new_n823), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n1137));
  XNOR2_X1  g0937(.A(new_n1136), .B(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n844), .A2(G143), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1003), .A2(G50), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n280), .B1(new_n903), .B2(G87), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n829), .A2(new_n247), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G68), .B2(new_n888), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G77), .B2(new_n1091), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1128), .A2(new_n1134), .B1(new_n1138), .B2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n791), .B(new_n1126), .C1(new_n1146), .C2(new_n863), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT117), .Z(new_n1148));
  AOI22_X1  g0948(.A1(new_n1052), .A2(new_n790), .B1(new_n1125), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(G390));
  NOR2_X1   g0950(.A1(new_n962), .A2(new_n975), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT39), .B1(new_n922), .B2(new_n936), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n973), .A2(new_n977), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n714), .B(new_n874), .C1(new_n748), .C2(new_n756), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n943), .B1(new_n1154), .B2(new_n971), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n937), .A2(new_n977), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT118), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n938), .A2(G330), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1158), .B1(new_n1159), .B2(new_n953), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n938), .A2(KEYINPUT118), .A3(G330), .A4(new_n943), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1153), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n971), .B1(new_n739), .B2(new_n878), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1164), .A2(new_n953), .B1(new_n364), .B2(new_n714), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n976), .B1(new_n975), .B2(new_n962), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1165), .A2(new_n1166), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1159), .A2(new_n953), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1163), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n474), .A2(G330), .A3(new_n781), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n981), .A2(new_n676), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1164), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n943), .B1(new_n938), .B2(G330), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1168), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1159), .A2(new_n953), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n757), .A2(new_n878), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1178), .A3(new_n972), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1170), .A2(new_n1181), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n1077), .A3(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1163), .B(new_n790), .C1(new_n1169), .C2(new_n1167), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT119), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1166), .A2(new_n803), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n884), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n791), .B1(new_n252), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n888), .A2(G150), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1191), .A2(KEYINPUT53), .B1(new_n831), .B2(new_n896), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(KEYINPUT53), .B2(new_n1191), .ZN(new_n1193));
  INV_X1    g0993(.A(G132), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(KEYINPUT54), .B(G143), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n823), .A2(new_n1194), .B1(new_n829), .B2(new_n1195), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n280), .B(new_n1196), .C1(G50), .C2(new_n903), .ZN(new_n1197));
  INV_X1    g0997(.A(G125), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1193), .B(new_n1197), .C1(new_n1198), .C2(new_n843), .ZN(new_n1199));
  INV_X1    g0999(.A(G128), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n816), .A2(new_n1135), .B1(new_n1200), .B2(new_n837), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n282), .B(new_n821), .C1(G107), .C2(new_n1003), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n844), .A2(G294), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n893), .A2(G97), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G116), .A2(new_n824), .B1(new_n903), .B2(G68), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n816), .A2(new_n382), .B1(new_n847), .B2(new_n837), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n1199), .A2(new_n1201), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1190), .B1(new_n1208), .B2(new_n806), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1188), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1184), .A2(new_n1187), .A3(new_n1210), .ZN(G378));
  NAND3_X1  g1011(.A1(new_n974), .A2(new_n978), .A3(new_n979), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n912), .B1(new_n963), .B2(new_n964), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT121), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n269), .B(new_n914), .C1(new_n307), .C2(new_n310), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n269), .A2(new_n914), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n304), .A2(new_n311), .A3(new_n306), .A4(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1218), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1225), .A2(KEYINPUT121), .A3(new_n1219), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n958), .A2(new_n1213), .A3(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n958), .B2(new_n1213), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1212), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n957), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n950), .A2(new_n953), .A3(new_n964), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n956), .B1(new_n1234), .B2(new_n955), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1213), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n1229), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n958), .A2(new_n1227), .A3(new_n1213), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n980), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1232), .A2(new_n1239), .A3(KEYINPUT122), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1172), .B1(new_n1170), .B2(new_n1181), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT122), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1212), .C1(new_n1228), .C2(new_n1231), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT57), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1078), .B1(new_n1247), .B2(new_n1241), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1240), .A2(new_n790), .A3(new_n1243), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n883), .B1(new_n201), .B2(new_n884), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n837), .A2(new_n1198), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1195), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n888), .A2(new_n1253), .B1(new_n893), .B2(G137), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1254), .B1(new_n1200), .B2(new_n823), .C1(new_n1194), .C2(new_n831), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n1252), .B(new_n1255), .C1(G150), .C2(new_n1091), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT120), .Z(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n844), .A2(G124), .ZN(new_n1261));
  AOI211_X1 g1061(.A(G33), .B(G41), .C1(new_n903), .C2(G159), .ZN(new_n1262));
  AND4_X1   g1062(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n816), .A2(new_n215), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n282), .A2(G41), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n382), .B2(new_n820), .C1(new_n220), .C2(new_n831), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n827), .A2(new_n202), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n997), .A2(new_n829), .B1(new_n373), .B2(new_n823), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n847), .B2(new_n843), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1264), .B(new_n1270), .C1(G116), .C2(new_n891), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT58), .ZN(new_n1272));
  AOI211_X1 g1072(.A(G50), .B(new_n1265), .C1(new_n253), .C2(new_n292), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(KEYINPUT58), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1263), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1251), .B1(new_n1275), .B2(new_n863), .C1(new_n1227), .C2(new_n804), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1250), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1249), .A2(new_n1277), .ZN(G375));
  INV_X1    g1078(.A(new_n1172), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1180), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n1056), .A3(new_n1181), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n953), .A2(new_n803), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n791), .B1(G68), .B2(new_n1189), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1001), .A2(new_n280), .ZN(new_n1285));
  XOR2_X1   g1085(.A(new_n1285), .B(KEYINPUT123), .Z(new_n1286));
  OAI211_X1 g1086(.A(new_n1286), .B(new_n1092), .C1(new_n629), .C2(new_n837), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n220), .A2(new_n820), .B1(new_n823), .B2(new_n847), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G107), .B2(new_n893), .ZN(new_n1289));
  OAI221_X1 g1089(.A(new_n1289), .B1(new_n508), .B2(new_n831), .C1(new_n850), .C2(new_n843), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n280), .B(new_n1267), .C1(new_n1003), .C2(new_n1253), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n896), .A2(new_n823), .B1(new_n820), .B2(new_n1135), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(G150), .B2(new_n893), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1291), .B(new_n1293), .C1(new_n1200), .C2(new_n843), .ZN(new_n1294));
  OAI22_X1  g1094(.A1(new_n816), .A2(new_n201), .B1(new_n1194), .B2(new_n837), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n1287), .A2(new_n1290), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1284), .B1(new_n1296), .B2(new_n806), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n1180), .A2(new_n790), .B1(new_n1283), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1282), .A2(new_n1298), .ZN(G381));
  OR4_X1    g1099(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n790), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1047), .A2(KEYINPUT109), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1052), .A2(new_n1049), .A3(new_n1032), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n783), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1301), .B1(new_n1304), .B2(new_n1055), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(G390), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1024), .A3(new_n1308), .ZN(new_n1309));
  OR4_X1    g1109(.A1(G378), .A2(new_n1300), .A3(new_n1309), .A4(G375), .ZN(G407));
  AND3_X1   g1110(.A1(new_n1184), .A2(new_n1187), .A3(new_n1210), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n713), .A2(G213), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(KEYINPUT124), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G407), .B(G213), .C1(G375), .C2(new_n1314), .ZN(G409));
  XNOR2_X1  g1115(.A(G393), .B(new_n868), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1024), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1317), .B(G390), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1308), .B1(new_n1307), .B2(new_n1024), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1316), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(G387), .A2(G390), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1316), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(new_n1322), .A3(new_n1309), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1320), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1249), .A2(G378), .A3(new_n1277), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1232), .A2(new_n1239), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT125), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1232), .A2(new_n1239), .A3(KEYINPUT125), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1328), .A2(new_n790), .A3(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1240), .A2(new_n1241), .A3(new_n1056), .A4(new_n1243), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1330), .A2(new_n1276), .A3(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1311), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1325), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1313), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1181), .A2(new_n1077), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT60), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1279), .A2(new_n1280), .A3(new_n1338), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1337), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1298), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n909), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1341), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1345), .A2(new_n1339), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G384), .B(new_n1298), .C1(new_n1346), .C2(new_n1337), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1313), .A2(G2897), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1344), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1344), .B2(new_n1347), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(KEYINPUT61), .B1(new_n1336), .B2(new_n1351), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1344), .A2(new_n1347), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1334), .A2(new_n1335), .A3(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT63), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1313), .B1(new_n1325), .B2(new_n1333), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1357), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1324), .A2(new_n1352), .A3(new_n1356), .A4(new_n1358), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1357), .A2(KEYINPUT62), .A3(new_n1353), .ZN(new_n1360));
  AOI21_X1  g1160(.A(KEYINPUT62), .B1(new_n1357), .B2(new_n1353), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n1352), .B(KEYINPUT126), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1362));
  AND3_X1   g1162(.A1(new_n1320), .A2(new_n1323), .A3(KEYINPUT127), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT127), .B1(new_n1320), .B2(new_n1323), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1362), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT62), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1354), .A2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1357), .A2(KEYINPUT62), .A3(new_n1353), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(KEYINPUT126), .B1(new_n1370), .B2(new_n1352), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1359), .B1(new_n1366), .B2(new_n1371), .ZN(G405));
  XNOR2_X1  g1172(.A(G375), .B(G378), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1373), .B(new_n1353), .ZN(new_n1374));
  XNOR2_X1  g1174(.A(new_n1374), .B(new_n1324), .ZN(G402));
endmodule


