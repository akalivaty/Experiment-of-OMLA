//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  AND2_X1   g000(.A1(G116), .A2(G119), .ZN(new_n187));
  NOR2_X1   g001(.A1(G116), .A2(G119), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n191), .A2(KEYINPUT5), .A3(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(G113), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT2), .A2(G113), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n196), .B(new_n197), .C1(new_n187), .C2(new_n188), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n193), .A2(new_n198), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G101), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n198), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n198), .B2(KEYINPUT68), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n196), .A2(new_n197), .ZN(new_n220));
  OAI22_X1  g034(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n189), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n198), .A2(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT69), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n220), .A2(new_n189), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n198), .A2(KEYINPUT68), .A3(new_n217), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n216), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n213), .A2(G101), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n228), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n206), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n212), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT86), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT6), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  AOI211_X1 g052(.A(new_n236), .B(new_n212), .C1(new_n227), .C2(new_n233), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT87), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n221), .A2(new_n226), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n233), .A3(new_n215), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n211), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n236), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n211), .A3(new_n237), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT6), .A4(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT64), .A3(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n253), .A2(new_n261), .B1(new_n264), .B2(new_n250), .ZN(new_n265));
  INV_X1    g079(.A(G125), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n248), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n256), .A2(new_n258), .B1(G143), .B2(new_n255), .ZN(new_n268));
  OAI22_X1  g082(.A1(new_n268), .A2(new_n252), .B1(new_n263), .B2(new_n249), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT88), .A3(G125), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n260), .B(KEYINPUT66), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G128), .ZN(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT66), .B1(new_n275), .B2(new_n260), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n261), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n260), .A2(new_n262), .A3(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n275), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n267), .B(new_n270), .C1(G125), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G224), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n282), .A2(new_n285), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OR3_X1    g102(.A1(new_n234), .A2(KEYINPUT6), .A3(new_n237), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n240), .A2(new_n247), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n282), .A2(new_n291), .A3(new_n284), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n236), .B(KEYINPUT8), .Z(new_n293));
  AOI21_X1  g107(.A(new_n210), .B1(new_n193), .B2(new_n198), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n212), .B2(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n246), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  OAI22_X1  g110(.A1(new_n286), .A2(new_n287), .B1(KEYINPUT7), .B2(new_n285), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G210), .B1(G237), .B2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n290), .A2(new_n298), .A3(new_n300), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(KEYINPUT89), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  XOR2_X1   g119(.A(new_n305), .B(KEYINPUT85), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n303), .A2(KEYINPUT89), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n304), .A2(new_n308), .A3(KEYINPUT90), .A4(new_n307), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G217), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(G234), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT78), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n266), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n318), .A4(G125), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n320), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n255), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n320), .A2(new_n322), .A3(G146), .A4(new_n325), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  XNOR2_X1  g144(.A(G119), .B(G128), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G110), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(KEYINPUT23), .C1(new_n335), .C2(G119), .ZN(new_n336));
  INV_X1    g150(.A(G119), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G128), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n336), .B(new_n338), .C1(new_n334), .C2(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n329), .B(new_n332), .C1(new_n333), .C2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G125), .B(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n255), .ZN(new_n344));
  AOI21_X1  g158(.A(G110), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n330), .A2(new_n331), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n328), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT22), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n342), .A2(new_n347), .A3(new_n351), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n315), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n317), .B1(new_n355), .B2(KEYINPUT25), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n353), .A2(new_n357), .A3(new_n315), .A4(new_n354), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n356), .A2(new_n361), .A3(new_n358), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n354), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n316), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NOR2_X1   g182(.A1(G472), .A2(G902), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT11), .ZN(new_n372));
  INV_X1    g186(.A(G134), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(G137), .ZN(new_n374));
  INV_X1    g188(.A(G137), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT11), .A3(G134), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(G137), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n374), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n373), .A2(G137), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n375), .A2(G134), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n277), .B2(new_n280), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n374), .A2(new_n378), .A3(new_n376), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G131), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n269), .B1(new_n386), .B2(new_n379), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n371), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT67), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT67), .B(new_n371), .C1(new_n384), .C2(new_n387), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT70), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n379), .A2(new_n382), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n379), .B2(new_n382), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n281), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n386), .A2(new_n379), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n265), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n390), .A2(new_n241), .A3(new_n391), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT31), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n260), .B1(new_n271), .B2(new_n272), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G128), .A3(new_n273), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n279), .B1(new_n405), .B2(new_n261), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n379), .A2(new_n382), .A3(new_n392), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n398), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n241), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT26), .B(G101), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(G237), .A2(G953), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G210), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT72), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n414), .B(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n411), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n400), .A2(new_n401), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n401), .B1(new_n400), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n396), .A2(new_n226), .A3(new_n221), .A4(new_n398), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n241), .B1(new_n387), .B2(new_n384), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT28), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT73), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n411), .B2(KEYINPUT28), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(KEYINPUT73), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n418), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n370), .B1(new_n422), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT74), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n368), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n400), .A2(new_n419), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT31), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n400), .A2(new_n401), .A3(new_n419), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n369), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n426), .A2(new_n428), .A3(new_n443), .A4(new_n430), .ZN(new_n444));
  INV_X1    g258(.A(new_n418), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n428), .A2(new_n430), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n410), .A2(new_n241), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n423), .A3(KEYINPUT75), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n410), .A2(new_n450), .A3(new_n241), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(KEYINPUT28), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT76), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n454), .A3(KEYINPUT28), .A4(new_n451), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n447), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n446), .B1(new_n456), .B2(new_n443), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n400), .A2(new_n423), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n445), .ZN(new_n459));
  AOI21_X1  g273(.A(G902), .B1(new_n459), .B2(new_n443), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G472), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n367), .B1(new_n442), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n279), .B1(new_n206), .B2(new_n209), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n277), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n335), .B1(new_n260), .B2(KEYINPUT1), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n264), .A2(new_n468), .B1(new_n278), .B2(new_n275), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n210), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n471), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n397), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n466), .A2(new_n277), .B1(new_n210), .B2(new_n469), .ZN(new_n474));
  INV_X1    g288(.A(new_n397), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n474), .A2(new_n475), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT81), .B1(new_n478), .B2(KEYINPUT12), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n465), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G140), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n283), .A2(G227), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT10), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n470), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n210), .A2(KEYINPUT10), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n485), .B1(new_n406), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n264), .A2(new_n250), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n215), .B(new_n488), .C1(new_n268), .C2(new_n252), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n231), .B2(new_n232), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n483), .B1(new_n491), .B2(new_n475), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n471), .A2(KEYINPUT12), .A3(new_n397), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT84), .A3(new_n476), .A4(new_n472), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n480), .A2(new_n492), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n490), .ZN(new_n498));
  INV_X1    g312(.A(new_n486), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n499), .A2(new_n281), .B1(new_n484), .B2(new_n470), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n475), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n397), .B1(new_n487), .B2(new_n490), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n483), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G469), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n464), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n483), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n476), .A3(new_n472), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n501), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n492), .A2(new_n502), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT82), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n501), .B1(new_n477), .B2(new_n479), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n483), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n492), .A2(new_n502), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(G902), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n507), .B1(new_n518), .B2(new_n506), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT82), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n315), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n464), .A3(G469), .ZN(new_n523));
  XNOR2_X1  g337(.A(KEYINPUT9), .B(G234), .ZN(new_n524));
  OAI21_X1  g338(.A(G221), .B1(new_n524), .B2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G475), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n415), .A2(G143), .A3(G214), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(G143), .B1(new_n415), .B2(G214), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(KEYINPUT18), .A2(G131), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n343), .B(new_n255), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT91), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n343), .A2(new_n255), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(new_n538), .A3(new_n344), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n533), .A2(new_n534), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G237), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n283), .A3(G214), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n257), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n377), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT92), .ZN(new_n545));
  OAI21_X1  g359(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n547), .A3(new_n377), .A4(new_n528), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT17), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT17), .B(G131), .C1(new_n529), .C2(new_n530), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n327), .A2(new_n328), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n549), .A2(new_n550), .B1(new_n552), .B2(KEYINPUT94), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n327), .A2(new_n554), .A3(new_n328), .A4(new_n551), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n540), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(G113), .B(G122), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(new_n199), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT95), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n540), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n552), .A2(KEYINPUT94), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n545), .A2(new_n550), .A3(new_n546), .A4(new_n548), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n565));
  INV_X1    g379(.A(new_n558), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n556), .A2(new_n558), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n527), .B1(new_n570), .B2(KEYINPUT96), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT96), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n564), .A2(new_n566), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n559), .B2(new_n567), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n574), .B2(G902), .ZN(new_n575));
  AND2_X1   g389(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n576));
  NOR2_X1   g390(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n343), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n343), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n328), .B1(new_n579), .B2(G146), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n549), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n566), .B1(new_n581), .B2(new_n540), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n569), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n527), .A2(new_n315), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT20), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT20), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n583), .A2(new_n587), .A3(new_n527), .A4(new_n315), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n571), .A2(new_n575), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n257), .A2(G128), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n335), .A2(G143), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n257), .A2(KEYINPUT98), .A3(KEYINPUT13), .A4(G128), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n593), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G134), .ZN(new_n598));
  INV_X1    g412(.A(G122), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G116), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n191), .A2(G122), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n202), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n202), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT97), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  INV_X1    g420(.A(new_n604), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(new_n602), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n591), .A2(new_n595), .A3(new_n373), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n598), .A2(new_n605), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n591), .A2(new_n595), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G134), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n607), .B1(new_n612), .B2(new_n609), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n599), .A2(G116), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n202), .B1(new_n614), .B2(KEYINPUT14), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT14), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n600), .A2(new_n601), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(KEYINPUT99), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n524), .A2(new_n314), .A3(G953), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n610), .A2(new_n620), .A3(new_n622), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n621), .A2(KEYINPUT100), .A3(new_n623), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n315), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT101), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(KEYINPUT101), .A3(new_n315), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT15), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G478), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT102), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n632), .A2(new_n634), .A3(G478), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n631), .A2(new_n632), .B1(new_n634), .B2(G478), .ZN(new_n640));
  INV_X1    g454(.A(new_n638), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT102), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n283), .A2(G952), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(G234), .B2(G237), .ZN(new_n645));
  NAND2_X1  g459(.A1(G234), .A2(G237), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(G902), .A3(G953), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT103), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT21), .B(G898), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n645), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n589), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n526), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n313), .A2(new_n463), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT104), .B(G101), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G3));
  NAND2_X1  g470(.A1(new_n439), .A2(new_n315), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n433), .B1(G472), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n367), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n526), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n565), .B1(new_n564), .B2(new_n566), .ZN(new_n662));
  AOI211_X1 g476(.A(KEYINPUT95), .B(new_n558), .C1(new_n560), .C2(new_n563), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n569), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(KEYINPUT96), .A3(new_n315), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n575), .A2(new_n665), .A3(G475), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n586), .A2(new_n588), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n627), .A2(new_n669), .A3(new_n628), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n624), .A2(KEYINPUT33), .A3(new_n626), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(G478), .A3(new_n315), .ZN(new_n673));
  INV_X1    g487(.A(G478), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n629), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n290), .A2(new_n298), .A3(new_n300), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n300), .B1(new_n290), .B2(new_n298), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n307), .B(new_n651), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n661), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT34), .B(G104), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  NAND4_X1  g498(.A1(new_n666), .A2(new_n639), .A3(new_n642), .A4(new_n667), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n661), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NAND2_X1  g503(.A1(new_n348), .A2(KEYINPUT105), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n342), .A2(new_n691), .A3(new_n347), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n365), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n360), .A2(new_n696), .A3(new_n362), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT106), .B1(new_n658), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n657), .A2(G472), .ZN(new_n699));
  AND4_X1   g513(.A1(KEYINPUT106), .A2(new_n699), .A3(new_n440), .A4(new_n697), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n313), .A2(new_n653), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  OAI211_X1 g519(.A(new_n697), .B(new_n307), .C1(new_n678), .C2(new_n679), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n442), .B2(new_n462), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n519), .A2(new_n523), .A3(new_n525), .ZN(new_n708));
  INV_X1    g522(.A(new_n685), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT108), .B(G900), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n645), .B1(new_n648), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n709), .A2(new_n710), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT109), .B1(new_n685), .B2(new_n712), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n707), .A2(new_n708), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XOR2_X1   g531(.A(new_n712), .B(KEYINPUT39), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n708), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT40), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n304), .A2(new_n308), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT38), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n643), .ZN(new_n725));
  INV_X1    g539(.A(new_n697), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n725), .A2(new_n668), .A3(new_n307), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n458), .A2(new_n445), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n449), .A2(new_n451), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n315), .B1(new_n732), .B2(new_n445), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n433), .A2(new_n434), .A3(new_n368), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT32), .B1(new_n440), .B2(KEYINPUT74), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n728), .B2(new_n727), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n721), .A2(new_n724), .A3(new_n729), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G143), .ZN(G45));
  NAND3_X1  g555(.A1(new_n668), .A2(new_n676), .A3(new_n713), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n707), .A2(new_n708), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  NAND2_X1  g559(.A1(new_n442), .A2(new_n462), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n505), .A2(new_n506), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n505), .A2(new_n506), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n525), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n746), .A2(new_n681), .A3(new_n659), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n659), .A3(new_n686), .A4(new_n750), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G116), .ZN(G18));
  AND4_X1   g569(.A1(new_n589), .A2(new_n643), .A3(new_n651), .A4(new_n697), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n307), .B1(new_n678), .B2(new_n679), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n749), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n746), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NOR3_X1   g574(.A1(new_n757), .A2(new_n589), .A3(new_n643), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n422), .B1(new_n456), .B2(new_n445), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n369), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n699), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n367), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n749), .A2(new_n650), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  NOR2_X1   g582(.A1(new_n764), .A2(new_n726), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n758), .A3(new_n743), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n306), .B1(new_n304), .B2(new_n308), .ZN(new_n773));
  INV_X1    g587(.A(new_n525), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n775));
  AOI211_X1 g589(.A(G469), .B(G902), .C1(new_n497), .C2(new_n504), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n514), .A2(new_n516), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n506), .B1(new_n777), .B2(new_n315), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n775), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n510), .A2(new_n511), .ZN(new_n780));
  OAI21_X1  g594(.A(G469), .B1(new_n780), .B2(G902), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n748), .A2(new_n781), .A3(KEYINPUT111), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n774), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n746), .A2(new_n659), .A3(new_n773), .A4(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n772), .B1(new_n784), .B2(new_n742), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n440), .B(KEYINPUT32), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n367), .B1(new_n786), .B2(new_n462), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n742), .A2(new_n772), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n783), .A3(new_n773), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  NAND2_X1  g605(.A1(new_n714), .A2(new_n715), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n373), .ZN(G36));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n512), .B2(new_n517), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n795), .A2(KEYINPUT112), .A3(new_n506), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n780), .A2(KEYINPUT45), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT112), .B1(new_n795), .B2(new_n506), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(G469), .A2(G902), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n776), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n525), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n589), .A2(new_n676), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT43), .ZN(new_n808));
  INV_X1    g622(.A(new_n676), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n668), .A2(KEYINPUT43), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n658), .A2(new_n726), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT44), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n722), .A2(new_n307), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n806), .A2(new_n718), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  NAND2_X1  g633(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n804), .A2(new_n821), .A3(new_n525), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n814), .A2(new_n746), .A3(new_n659), .A4(new_n742), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  INV_X1    g639(.A(new_n747), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n776), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT49), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n807), .A2(new_n367), .A3(new_n306), .A4(new_n774), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n723), .A3(new_n738), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n814), .A2(new_n749), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n738), .A3(new_n659), .A4(new_n645), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n677), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n808), .A2(new_n810), .A3(new_n645), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n758), .A3(new_n765), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n833), .A2(new_n835), .A3(new_n644), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n787), .A3(new_n831), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT48), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n836), .B2(new_n838), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n765), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n773), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n820), .A2(new_n822), .ZN(new_n846));
  INV_X1    g660(.A(new_n827), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n774), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n832), .A2(new_n668), .A3(new_n676), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n834), .A2(new_n769), .A3(new_n831), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n723), .A2(new_n306), .A3(new_n750), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n843), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n856), .A2(KEYINPUT120), .A3(KEYINPUT50), .ZN(new_n857));
  NOR2_X1   g671(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n855), .A2(new_n843), .A3(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT51), .B(new_n854), .C1(new_n857), .C2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n842), .B1(new_n851), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n822), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n821), .B1(new_n804), .B2(new_n525), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n850), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(KEYINPUT119), .A3(new_n773), .A4(new_n844), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT119), .ZN(new_n866));
  INV_X1    g680(.A(new_n850), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n820), .B2(new_n822), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n868), .B2(new_n845), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n857), .A2(new_n859), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n853), .A3(new_n852), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n865), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT51), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n861), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n726), .A2(new_n875), .A3(new_n713), .ZN(new_n876));
  OAI21_X1  g690(.A(KEYINPUT115), .B1(new_n697), .B2(new_n712), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n761), .A2(new_n878), .A3(new_n737), .A4(new_n783), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n716), .A2(new_n744), .A3(new_n770), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n880), .A2(KEYINPUT116), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n881), .B1(new_n880), .B2(KEYINPUT116), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n589), .A2(KEYINPUT113), .A3(new_n809), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n668), .B2(new_n676), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n885), .A2(new_n887), .A3(new_n650), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n313), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n313), .A2(new_n888), .A3(KEYINPUT114), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n661), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n636), .A2(new_n638), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n589), .A2(new_n894), .A3(new_n651), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n526), .A2(new_n660), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n313), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n654), .A2(new_n702), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n793), .B1(new_n785), .B2(new_n789), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n751), .A2(new_n754), .A3(new_n759), .A4(new_n767), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n773), .A2(new_n697), .A3(new_n713), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n668), .A2(new_n894), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n708), .A2(new_n746), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n764), .A2(new_n677), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n783), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n893), .A2(new_n898), .A3(new_n899), .A4(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n884), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(KEYINPUT53), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n880), .B(KEYINPUT52), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT54), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT117), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n908), .B2(new_n911), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(new_n909), .B2(KEYINPUT53), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n918));
  OAI211_X1 g732(.A(KEYINPUT117), .B(new_n912), .C1(new_n908), .C2(new_n911), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n874), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(G952), .A2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n830), .B1(new_n921), .B2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n283), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n916), .A2(new_n915), .ZN(new_n926));
  AND4_X1   g740(.A1(new_n893), .A2(new_n898), .A3(new_n899), .A4(new_n907), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n927), .B(KEYINPUT53), .C1(new_n883), .C2(new_n882), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n240), .A2(new_n247), .A3(new_n289), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n288), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(KEYINPUT56), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n929), .A2(new_n939), .A3(G210), .A4(G902), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(new_n933), .ZN(G51));
  XOR2_X1   g756(.A(new_n800), .B(KEYINPUT57), .Z(new_n943));
  AOI21_X1  g757(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n918), .A2(new_n926), .A3(new_n919), .A4(new_n928), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n497), .A2(new_n504), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n929), .A2(G902), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(new_n799), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n924), .B1(new_n948), .B2(new_n950), .ZN(G54));
  AOI21_X1  g765(.A(new_n315), .B1(new_n917), .B2(new_n919), .ZN(new_n952));
  NAND2_X1  g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n583), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n584), .A2(new_n953), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n929), .A2(G902), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n925), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT123), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n584), .B1(new_n949), .B2(new_n953), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT123), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n925), .A4(new_n957), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(new_n920), .A2(new_n914), .ZN(new_n964));
  NAND2_X1  g778(.A1(G478), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT59), .Z(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n672), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n672), .A2(new_n967), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n929), .A2(KEYINPUT54), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n920), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n968), .A2(new_n924), .A3(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n695), .B(KEYINPUT124), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n929), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n974), .B1(new_n917), .B2(new_n919), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n925), .B(new_n977), .C1(new_n978), .C2(new_n364), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n929), .A2(new_n975), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n924), .B1(new_n982), .B2(new_n363), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(KEYINPUT61), .A3(new_n977), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(G66));
  INV_X1    g799(.A(new_n900), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n893), .A2(new_n898), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G224), .A2(G953), .ZN(new_n988));
  OAI22_X1  g802(.A1(new_n987), .A2(G953), .B1(new_n649), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n931), .B1(G898), .B2(new_n283), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(G69));
  NAND4_X1  g805(.A1(new_n806), .A2(new_n718), .A3(new_n761), .A4(new_n787), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n716), .A2(new_n744), .A3(new_n770), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n899), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n824), .A2(new_n818), .A3(new_n992), .A4(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n995), .A2(G953), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n390), .A2(new_n391), .A3(new_n399), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(new_n579), .Z(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n740), .A2(new_n993), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n1000), .A2(KEYINPUT62), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n885), .A2(new_n887), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n589), .B2(new_n894), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n463), .A2(new_n773), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1003), .A2(new_n719), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n1000), .B2(KEYINPUT62), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1001), .A2(new_n1006), .A3(new_n818), .A4(new_n824), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n283), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n996), .A2(new_n999), .B1(new_n1008), .B2(new_n998), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT126), .Z(new_n1011));
  OAI21_X1  g825(.A(new_n999), .B1(new_n995), .B2(G953), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT125), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1009), .B(new_n1013), .ZN(G72));
  XNOR2_X1  g828(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n1007), .B2(new_n987), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n924), .B1(new_n1018), .B2(new_n731), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1017), .B1(new_n995), .B2(new_n987), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n459), .ZN(new_n1021));
  INV_X1    g835(.A(new_n459), .ZN(new_n1022));
  AND3_X1   g836(.A1(new_n1022), .A2(new_n730), .A3(new_n1017), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n910), .B2(new_n913), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(G57));
endmodule


