

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591;

  XOR2_X1 U321 ( .A(G162GAT), .B(G50GAT), .Z(n405) );
  XNOR2_X1 U322 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U323 ( .A(n467), .B(n466), .ZN(n572) );
  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n466) );
  XNOR2_X1 U325 ( .A(n407), .B(n406), .ZN(n408) );
  INV_X1 U326 ( .A(KEYINPUT11), .ZN(n411) );
  XNOR2_X1 U327 ( .A(n465), .B(KEYINPUT48), .ZN(n549) );
  OR2_X1 U328 ( .A1(n291), .A2(n572), .ZN(n469) );
  XOR2_X1 U329 ( .A(n367), .B(n366), .Z(n527) );
  XOR2_X1 U330 ( .A(n464), .B(KEYINPUT47), .Z(n289) );
  OR2_X1 U331 ( .A1(n456), .A2(n459), .ZN(n290) );
  NAND2_X1 U332 ( .A1(n527), .A2(n455), .ZN(n291) );
  AND2_X1 U333 ( .A1(n552), .A2(n558), .ZN(n461) );
  XOR2_X1 U334 ( .A(G155GAT), .B(G22GAT), .Z(n376) );
  INV_X1 U335 ( .A(KEYINPUT24), .ZN(n298) );
  XNOR2_X1 U336 ( .A(n299), .B(n298), .ZN(n300) );
  INV_X1 U337 ( .A(KEYINPUT31), .ZN(n425) );
  XNOR2_X1 U338 ( .A(n301), .B(n300), .ZN(n305) );
  XNOR2_X1 U339 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U340 ( .A(n428), .B(n427), .ZN(n430) );
  NAND2_X1 U341 ( .A1(n290), .A2(n289), .ZN(n465) );
  XNOR2_X1 U342 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U343 ( .A(n327), .B(KEYINPUT26), .Z(n574) );
  XNOR2_X1 U344 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U345 ( .A(n435), .B(KEYINPUT41), .Z(n558) );
  INV_X1 U346 ( .A(G106GAT), .ZN(n452) );
  XNOR2_X1 U347 ( .A(n475), .B(KEYINPUT58), .ZN(n476) );
  XNOR2_X1 U348 ( .A(n452), .B(KEYINPUT44), .ZN(n453) );
  XNOR2_X1 U349 ( .A(n477), .B(n476), .ZN(G1351GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n293) );
  XNOR2_X1 U351 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n292) );
  XNOR2_X1 U352 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U353 ( .A(KEYINPUT88), .B(n376), .Z(n295) );
  XNOR2_X1 U354 ( .A(G218GAT), .B(n405), .ZN(n294) );
  XNOR2_X1 U355 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U356 ( .A(n297), .B(n296), .Z(n301) );
  NAND2_X1 U357 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT87), .Z(n303) );
  XNOR2_X1 U359 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n353) );
  XNOR2_X1 U361 ( .A(n353), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n311) );
  XOR2_X1 U363 ( .A(G197GAT), .B(KEYINPUT21), .Z(n307) );
  XNOR2_X1 U364 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n307), .B(n306), .ZN(n330) );
  XOR2_X1 U366 ( .A(G78GAT), .B(KEYINPUT71), .Z(n309) );
  XNOR2_X1 U367 ( .A(G148GAT), .B(G106GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n421) );
  XOR2_X1 U369 ( .A(n330), .B(n421), .Z(n310) );
  XOR2_X1 U370 ( .A(n311), .B(n310), .Z(n455) );
  INV_X1 U371 ( .A(n455), .ZN(n341) );
  XOR2_X1 U372 ( .A(n341), .B(KEYINPUT67), .Z(n312) );
  XOR2_X1 U373 ( .A(n312), .B(KEYINPUT28), .Z(n521) );
  XOR2_X1 U374 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n420) );
  XOR2_X1 U375 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n314) );
  XNOR2_X1 U376 ( .A(G183GAT), .B(G169GAT), .ZN(n313) );
  XNOR2_X1 U377 ( .A(n314), .B(n313), .ZN(n316) );
  XOR2_X1 U378 ( .A(G190GAT), .B(KEYINPUT17), .Z(n315) );
  XOR2_X1 U379 ( .A(n316), .B(n315), .Z(n336) );
  XNOR2_X1 U380 ( .A(G120GAT), .B(G99GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n317), .B(G71GAT), .ZN(n429) );
  XOR2_X1 U382 ( .A(G134GAT), .B(G43GAT), .Z(n401) );
  XOR2_X1 U383 ( .A(n429), .B(n401), .Z(n319) );
  NAND2_X1 U384 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U385 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U386 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n321) );
  XNOR2_X1 U387 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n320) );
  XNOR2_X1 U388 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U389 ( .A(n323), .B(n322), .Z(n325) );
  XOR2_X1 U390 ( .A(KEYINPUT0), .B(G127GAT), .Z(n359) );
  XOR2_X1 U391 ( .A(G113GAT), .B(G15GAT), .Z(n443) );
  XNOR2_X1 U392 ( .A(n359), .B(n443), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U394 ( .A(n336), .B(n326), .Z(n505) );
  INV_X1 U395 ( .A(n505), .ZN(n537) );
  NAND2_X1 U396 ( .A1(n537), .A2(n341), .ZN(n327) );
  INV_X1 U397 ( .A(n574), .ZN(n338) );
  XOR2_X1 U398 ( .A(G8GAT), .B(G92GAT), .Z(n329) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U400 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U401 ( .A(n331), .B(n330), .Z(n335) );
  XNOR2_X1 U402 ( .A(G218GAT), .B(G36GAT), .ZN(n332) );
  XNOR2_X1 U403 ( .A(n332), .B(KEYINPUT74), .ZN(n410) );
  XNOR2_X1 U404 ( .A(G64GAT), .B(G204GAT), .ZN(n333) );
  XNOR2_X1 U405 ( .A(n333), .B(G176GAT), .ZN(n431) );
  XNOR2_X1 U406 ( .A(n410), .B(n431), .ZN(n334) );
  XNOR2_X1 U407 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U408 ( .A(n337), .B(n336), .Z(n529) );
  INV_X1 U409 ( .A(n529), .ZN(n503) );
  XOR2_X1 U410 ( .A(n503), .B(KEYINPUT27), .Z(n369) );
  NOR2_X1 U411 ( .A1(n338), .A2(n369), .ZN(n339) );
  XNOR2_X1 U412 ( .A(KEYINPUT95), .B(n339), .ZN(n344) );
  NOR2_X1 U413 ( .A1(n529), .A2(n537), .ZN(n340) );
  NOR2_X1 U414 ( .A1(n341), .A2(n340), .ZN(n342) );
  XNOR2_X1 U415 ( .A(KEYINPUT25), .B(n342), .ZN(n343) );
  NAND2_X1 U416 ( .A1(n344), .A2(n343), .ZN(n368) );
  XOR2_X1 U417 ( .A(KEYINPUT92), .B(G57GAT), .Z(n346) );
  XNOR2_X1 U418 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n345) );
  XNOR2_X1 U419 ( .A(n346), .B(n345), .ZN(n367) );
  XOR2_X1 U420 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n348) );
  XNOR2_X1 U421 ( .A(G113GAT), .B(G120GAT), .ZN(n347) );
  XNOR2_X1 U422 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U423 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n350) );
  XNOR2_X1 U424 ( .A(KEYINPUT94), .B(G1GAT), .ZN(n349) );
  XNOR2_X1 U425 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U426 ( .A(n352), .B(n351), .Z(n365) );
  XOR2_X1 U427 ( .A(n353), .B(KEYINPUT91), .Z(n355) );
  NAND2_X1 U428 ( .A1(G225GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U429 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U430 ( .A(G148GAT), .B(G155GAT), .Z(n357) );
  XNOR2_X1 U431 ( .A(G162GAT), .B(G134GAT), .ZN(n356) );
  XNOR2_X1 U432 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U433 ( .A(n358), .B(G85GAT), .Z(n361) );
  XNOR2_X1 U434 ( .A(G29GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U435 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U436 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U437 ( .A(n365), .B(n364), .ZN(n366) );
  NAND2_X1 U438 ( .A1(n368), .A2(n527), .ZN(n372) );
  XOR2_X1 U439 ( .A(KEYINPUT84), .B(n505), .Z(n370) );
  INV_X1 U440 ( .A(n521), .ZN(n510) );
  OR2_X1 U441 ( .A1(n369), .A2(n527), .ZN(n551) );
  NOR2_X1 U442 ( .A1(n510), .A2(n551), .ZN(n535) );
  NAND2_X1 U443 ( .A1(n370), .A2(n535), .ZN(n371) );
  NAND2_X1 U444 ( .A1(n372), .A2(n371), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n373), .B(KEYINPUT96), .ZN(n484) );
  XOR2_X1 U446 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n375) );
  XNOR2_X1 U447 ( .A(KEYINPUT77), .B(KEYINPUT79), .ZN(n374) );
  XNOR2_X1 U448 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U449 ( .A(G78GAT), .B(G211GAT), .Z(n378) );
  XOR2_X1 U450 ( .A(G1GAT), .B(G8GAT), .Z(n446) );
  XNOR2_X1 U451 ( .A(n376), .B(n446), .ZN(n377) );
  XNOR2_X1 U452 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U453 ( .A(n380), .B(n379), .Z(n382) );
  NAND2_X1 U454 ( .A1(G231GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U456 ( .A(n383), .B(KEYINPUT80), .Z(n387) );
  XOR2_X1 U457 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n385) );
  XNOR2_X1 U458 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n384) );
  XNOR2_X1 U459 ( .A(n385), .B(n384), .ZN(n432) );
  XNOR2_X1 U460 ( .A(n432), .B(KEYINPUT15), .ZN(n386) );
  XNOR2_X1 U461 ( .A(n387), .B(n386), .ZN(n395) );
  XOR2_X1 U462 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n389) );
  XNOR2_X1 U463 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U464 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U465 ( .A(G71GAT), .B(G15GAT), .Z(n391) );
  XNOR2_X1 U466 ( .A(G127GAT), .B(G183GAT), .ZN(n390) );
  XNOR2_X1 U467 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U468 ( .A(n393), .B(n392), .Z(n394) );
  XOR2_X1 U469 ( .A(n395), .B(n394), .Z(n584) );
  INV_X1 U470 ( .A(n584), .ZN(n471) );
  AND2_X1 U471 ( .A1(n484), .A2(n471), .ZN(n396) );
  XNOR2_X1 U472 ( .A(n396), .B(KEYINPUT102), .ZN(n418) );
  INV_X1 U473 ( .A(KEYINPUT36), .ZN(n417) );
  XOR2_X1 U474 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n398) );
  XNOR2_X1 U475 ( .A(G190GAT), .B(KEYINPUT65), .ZN(n397) );
  XNOR2_X1 U476 ( .A(n398), .B(n397), .ZN(n416) );
  XOR2_X1 U477 ( .A(KEYINPUT66), .B(G106GAT), .Z(n400) );
  XNOR2_X1 U478 ( .A(G99GAT), .B(KEYINPUT72), .ZN(n399) );
  XNOR2_X1 U479 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U480 ( .A(n402), .B(n401), .Z(n409) );
  XNOR2_X1 U481 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n403), .B(KEYINPUT7), .ZN(n442) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G92GAT), .Z(n424) );
  XOR2_X1 U484 ( .A(n442), .B(n424), .Z(n407) );
  NAND2_X1 U485 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U486 ( .A(n409), .B(n408), .ZN(n414) );
  XNOR2_X1 U487 ( .A(n410), .B(KEYINPUT10), .ZN(n412) );
  XOR2_X1 U488 ( .A(n416), .B(n415), .Z(n481) );
  XNOR2_X1 U489 ( .A(n417), .B(n481), .ZN(n586) );
  NAND2_X1 U490 ( .A1(n418), .A2(n586), .ZN(n419) );
  XNOR2_X1 U491 ( .A(n420), .B(n419), .ZN(n497) );
  XOR2_X1 U492 ( .A(KEYINPUT32), .B(n421), .Z(n423) );
  NAND2_X1 U493 ( .A1(G230GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n424), .B(KEYINPUT33), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U497 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n456) );
  XNOR2_X1 U499 ( .A(n456), .B(KEYINPUT64), .ZN(n435) );
  INV_X1 U500 ( .A(n558), .ZN(n566) );
  XOR2_X1 U501 ( .A(G197GAT), .B(G22GAT), .Z(n437) );
  XNOR2_X1 U502 ( .A(G141GAT), .B(G43GAT), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U504 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n439) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(KEYINPUT68), .ZN(n438) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n451) );
  XOR2_X1 U508 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U509 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(n447) );
  XOR2_X1 U511 ( .A(n447), .B(n446), .Z(n449) );
  XNOR2_X1 U512 ( .A(G36GAT), .B(G50GAT), .ZN(n448) );
  XNOR2_X1 U513 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U514 ( .A(n451), .B(n450), .Z(n552) );
  NOR2_X1 U515 ( .A1(n566), .A2(n552), .ZN(n516) );
  NAND2_X1 U516 ( .A1(n497), .A2(n516), .ZN(n531) );
  NOR2_X1 U517 ( .A1(n521), .A2(n531), .ZN(n454) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(G1339GAT) );
  NAND2_X1 U519 ( .A1(n586), .A2(n584), .ZN(n457) );
  XOR2_X1 U520 ( .A(KEYINPUT45), .B(n457), .Z(n458) );
  INV_X1 U521 ( .A(n552), .ZN(n576) );
  NAND2_X1 U522 ( .A1(n458), .A2(n576), .ZN(n459) );
  XNOR2_X1 U523 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n460) );
  XNOR2_X1 U524 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U525 ( .A(n481), .ZN(n564) );
  NOR2_X1 U526 ( .A1(n462), .A2(n564), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n463), .A2(n471), .ZN(n464) );
  NAND2_X1 U528 ( .A1(n503), .A2(n549), .ZN(n467) );
  XOR2_X1 U529 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U531 ( .A1(n470), .A2(n505), .ZN(n567) );
  NOR2_X1 U532 ( .A1(n471), .A2(n567), .ZN(n474) );
  INV_X1 U533 ( .A(KEYINPUT124), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(G183GAT), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(G1350GAT) );
  NOR2_X1 U536 ( .A1(n481), .A2(n567), .ZN(n477) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n475) );
  NOR2_X1 U538 ( .A1(n576), .A2(n567), .ZN(n480) );
  INV_X1 U539 ( .A(G169GAT), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n478), .B(KEYINPUT122), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1348GAT) );
  NOR2_X1 U542 ( .A1(n576), .A2(n456), .ZN(n498) );
  NAND2_X1 U543 ( .A1(n584), .A2(n481), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(KEYINPUT81), .ZN(n483) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n483), .ZN(n485) );
  AND2_X1 U546 ( .A1(n485), .A2(n484), .ZN(n515) );
  NAND2_X1 U547 ( .A1(n498), .A2(n515), .ZN(n494) );
  NOR2_X1 U548 ( .A1(n527), .A2(n494), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT97), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NOR2_X1 U552 ( .A1(n529), .A2(n494), .ZN(n489) );
  XOR2_X1 U553 ( .A(KEYINPUT98), .B(n489), .Z(n490) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n537), .A2(n494), .ZN(n492) );
  XNOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n493), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n521), .A2(n494), .ZN(n495) );
  XOR2_X1 U560 ( .A(KEYINPUT100), .B(n495), .Z(n496) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n496), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n498), .A2(n497), .ZN(n499) );
  XOR2_X1 U563 ( .A(KEYINPUT38), .B(n499), .Z(n511) );
  INV_X1 U564 ( .A(n527), .ZN(n573) );
  NAND2_X1 U565 ( .A1(n511), .A2(n573), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT101), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U569 ( .A1(n511), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n511), .A2(n505), .ZN(n509) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n507) );
  XNOR2_X1 U573 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n514) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n518) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n522) );
  NOR2_X1 U582 ( .A1(n527), .A2(n522), .ZN(n517) );
  XOR2_X1 U583 ( .A(n518), .B(n517), .Z(G1332GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n519) );
  XOR2_X1 U585 ( .A(G64GAT), .B(n519), .Z(G1333GAT) );
  NOR2_X1 U586 ( .A1(n537), .A2(n522), .ZN(n520) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n526) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n524) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT109), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NOR2_X1 U593 ( .A1(n527), .A2(n531), .ZN(n528) );
  XOR2_X1 U594 ( .A(G85GAT), .B(n528), .Z(G1336GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n531), .ZN(n530) );
  XOR2_X1 U596 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U597 ( .A1(n537), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G99GAT), .B(n534), .ZN(G1338GAT) );
  NAND2_X1 U601 ( .A1(n535), .A2(n549), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n552), .A2(n545), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U606 ( .A1(n545), .A2(n558), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n542) );
  NAND2_X1 U610 ( .A1(n545), .A2(n584), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U612 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n564), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n574), .ZN(n550) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n552), .A2(n563), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT117), .B(n557), .Z(n560) );
  NAND2_X1 U626 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  XOR2_X1 U628 ( .A(G155GAT), .B(KEYINPUT119), .Z(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n584), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n571) );
  XOR2_X1 U634 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n569) );
  XNOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n581) );
  NOR2_X1 U640 ( .A1(n576), .A2(n581), .ZN(n578) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U646 ( .A(n581), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n587), .A2(n456), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n591) );
  XOR2_X1 U652 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(G1355GAT) );
endmodule

