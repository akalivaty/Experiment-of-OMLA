//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n460), .A2(G137), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  XNOR2_X1  g052(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n478), .B1(G136), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n466), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT68), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n479), .C2(new_n480), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n466), .A2(G114), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n466), .C1(new_n479), .C2(new_n480), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n460), .A2(new_n497), .A3(G138), .A4(new_n466), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G88), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n508));
  OAI211_X1 g083(.A(G50), .B(G543), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(G75), .A2(G543), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n505), .B2(G62), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n506), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G166));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n502), .B2(new_n503), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G51), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n502), .A2(new_n503), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n521), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n512), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n524), .A2(G90), .B1(new_n516), .B2(G52), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT5), .B(G543), .Z(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G651), .B1(new_n516), .B2(G43), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n524), .A2(G81), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n535), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(G91), .B2(new_n524), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n504), .A2(G53), .A3(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n516), .A2(new_n554), .A3(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(G299));
  OR2_X1    g132(.A1(new_n521), .A2(new_n525), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT72), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n521), .A2(new_n525), .A3(KEYINPUT72), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(G286));
  NAND2_X1  g137(.A1(new_n513), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g138(.A(G62), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n522), .B2(new_n523), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n565), .B2(new_n510), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n566), .A2(new_n567), .A3(new_n509), .A4(new_n506), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n563), .A2(new_n568), .ZN(G303));
  NAND2_X1  g144(.A1(new_n504), .A2(new_n505), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n570), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT74), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT75), .B(G651), .C1(new_n505), .C2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n577), .A2(new_n578), .B1(G49), .B2(new_n516), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n574), .A2(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n516), .A2(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n516), .A2(new_n583), .A3(G48), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n535), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G86), .B2(new_n524), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n524), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G47), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(new_n591), .B(new_n592), .C1(new_n512), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n570), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n535), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n516), .B2(G54), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n600), .A2(new_n604), .A3(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n595), .B1(G868), .B2(new_n609), .ZN(G284));
  OAI21_X1  g185(.A(new_n595), .B1(G868), .B2(new_n609), .ZN(G321));
  NOR2_X1   g186(.A1(G299), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n561), .B2(G868), .ZN(G297));
  AOI21_X1  g188(.A(new_n612), .B1(new_n561), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n615), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n618), .A2(KEYINPUT78), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT78), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G868), .C2(new_n541), .ZN(G323));
  XOR2_X1   g197(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n482), .A2(G2104), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n487), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n482), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n466), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n641), .B(new_n647), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n651), .B2(new_n649), .ZN(G401));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT81), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT17), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT82), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n660), .B(new_n662), .C1(new_n659), .C2(new_n655), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n655), .A2(new_n657), .A3(new_n661), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT18), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n661), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n665), .C1(new_n656), .C2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  INV_X1    g252(.A(new_n672), .ZN(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n677), .B(new_n681), .C1(new_n678), .C2(new_n680), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G20), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT23), .Z(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G299), .B2(G16), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1956), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G21), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G168), .B2(new_n690), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT94), .Z(new_n697));
  OAI21_X1  g272(.A(new_n694), .B1(new_n697), .B2(G1966), .ZN(new_n698));
  NOR2_X1   g273(.A1(G29), .A2(G33), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT92), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n482), .A2(G139), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n703), .B(new_n704), .C1(new_n466), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2072), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT93), .Z(new_n711));
  AOI211_X1 g286(.A(new_n698), .B(new_n711), .C1(G1966), .C2(new_n697), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n707), .B1(new_n713), .B2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G160), .B2(G29), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G2084), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT95), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n707), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n482), .A2(G141), .ZN(new_n720));
  NAND3_X1  g295(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT26), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n469), .A2(G105), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G129), .B2(new_n487), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n719), .B1(new_n725), .B2(new_n707), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT27), .B(G1996), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n707), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n487), .A2(G128), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G116), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n482), .B2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G2067), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n690), .A2(G5), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G171), .B2(new_n690), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G1961), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n718), .A2(new_n728), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n690), .A2(G4), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n609), .B2(new_n690), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G1348), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(G1348), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n707), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n707), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2090), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n690), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n541), .B2(new_n690), .ZN(new_n753));
  AOI22_X1  g328(.A1(new_n708), .A2(new_n709), .B1(G1341), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  NAND2_X1  g330(.A1(G164), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G27), .B2(G29), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n754), .B1(G1341), .B2(new_n753), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n759), .A2(new_n707), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n635), .B2(new_n707), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G2084), .B2(new_n716), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n757), .A2(new_n755), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n764), .B(new_n765), .C1(G1961), .C2(new_n740), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n751), .A2(new_n758), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n712), .A2(new_n747), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT96), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n690), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n690), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT87), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n774), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n690), .A2(G22), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT88), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n513), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT89), .B(G1971), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(G6), .A2(G16), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G305), .B2(new_n690), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G1981), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(G1981), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n777), .B(new_n782), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT90), .ZN(new_n791));
  MUX2_X1   g366(.A(G24), .B(G290), .S(G16), .Z(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT85), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1986), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n707), .A2(G25), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n487), .A2(G119), .ZN(new_n796));
  OAI21_X1  g371(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n797));
  INV_X1    g372(.A(G107), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G2105), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n482), .B2(G131), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n795), .B1(new_n802), .B2(new_n707), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  XOR2_X1   g379(.A(new_n803), .B(new_n804), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n794), .A2(new_n805), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n790), .A2(new_n791), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n791), .B1(new_n790), .B2(new_n806), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n788), .A2(new_n789), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n771), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n771), .A3(new_n810), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n770), .B1(new_n812), .B2(new_n813), .ZN(G311));
  INV_X1    g389(.A(new_n770), .ZN(new_n815));
  INV_X1    g390(.A(new_n813), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n811), .B2(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(new_n524), .A2(G93), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n516), .A2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n818), .B(new_n819), .C1(new_n512), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n609), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n540), .B(new_n821), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT97), .Z(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n829), .B2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n824), .B1(new_n831), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n801), .B(new_n627), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n496), .A2(new_n498), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n492), .A2(new_n493), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n486), .B2(G126), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n736), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(new_n725), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n725), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n706), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n487), .A2(G130), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  INV_X1    g424(.A(G118), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(G2105), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n482), .B2(G142), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n706), .B(new_n845), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n842), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n847), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n853), .B1(new_n847), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n836), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(new_n835), .A3(new_n856), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n859), .A2(new_n861), .A3(KEYINPUT102), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n489), .B(new_n635), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n473), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G37), .ZN(new_n868));
  INV_X1    g443(.A(new_n866), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n869), .A2(new_n859), .A3(new_n861), .A4(KEYINPUT102), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n617), .B(new_n827), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n600), .A2(new_n604), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(G299), .ZN(new_n877));
  INV_X1    g452(.A(G299), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT103), .A3(new_n605), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n879), .C1(new_n878), .C2(new_n605), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(KEYINPUT104), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n880), .B(KEYINPUT41), .Z(new_n883));
  INV_X1    g458(.A(new_n874), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n881), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G290), .B(KEYINPUT105), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n890), .A2(G288), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(G288), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G305), .B(new_n513), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n891), .B2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT42), .B1(new_n895), .B2(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n873), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n889), .A2(new_n903), .A3(KEYINPUT106), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n887), .B1(new_n882), .B2(new_n885), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n902), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n904), .A2(new_n905), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(G868), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT108), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n821), .A2(new_n619), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(KEYINPUT108), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n914), .B1(new_n910), .B2(G868), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n912), .A2(new_n915), .ZN(G295));
  NOR2_X1   g491(.A1(new_n912), .A2(new_n915), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g493(.A1(G301), .A2(new_n558), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(G286), .B2(G301), .ZN(new_n920));
  INV_X1    g495(.A(new_n827), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n880), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT110), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n883), .ZN(new_n927));
  INV_X1    g502(.A(new_n898), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(new_n880), .C1(new_n922), .C2(new_n923), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n927), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n927), .A2(new_n924), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n931), .B(new_n868), .C1(new_n932), .C2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n898), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n937));
  NAND4_X1  g512(.A1(new_n936), .A2(new_n868), .A3(new_n931), .A4(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n918), .B1(new_n934), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n937), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n868), .A3(new_n931), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n940), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n943), .B2(new_n918), .ZN(G397));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G164), .B2(G1384), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n465), .A2(new_n472), .A3(G40), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g525(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(KEYINPUT46), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n736), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n725), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n951), .A2(new_n952), .B1(new_n955), .B2(new_n948), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n949), .B2(new_n725), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n948), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n948), .A2(KEYINPUT111), .A3(new_n949), .A4(new_n725), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  INV_X1    g536(.A(new_n725), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n950), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n964), .B(KEYINPUT112), .Z(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n802), .A2(new_n804), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n966), .A2(new_n967), .B1(G2067), .B2(new_n736), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n957), .B1(new_n968), .B2(new_n948), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n801), .B(new_n804), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n948), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n965), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n948), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n969), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n585), .A2(new_n589), .A3(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT114), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n773), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT115), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  INV_X1    g564(.A(new_n984), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n585), .B2(new_n589), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n466), .B1(new_n461), .B2(new_n463), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n993), .A2(new_n471), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1384), .B1(new_n837), .B2(new_n839), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT49), .A3(new_n984), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n992), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n985), .B1(new_n988), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1000), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n563), .A2(G8), .A3(new_n568), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n563), .A2(KEYINPUT55), .A3(G8), .A4(new_n568), .ZN(new_n1009));
  INV_X1    g584(.A(G1971), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n995), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1011));
  NOR3_X1   g586(.A1(G164), .A2(new_n945), .A3(G1384), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n996), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G2090), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n995), .ZN(new_n1018));
  AOI221_X4 g593(.A(new_n999), .B1(new_n1008), .B2(new_n1009), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n574), .A2(G1976), .A3(new_n579), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1000), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(G8), .A3(new_n997), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1003), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n1004), .A2(new_n1005), .B1(new_n1020), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n999), .A2(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1031), .B2(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1019), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g608(.A(KEYINPUT116), .B(new_n999), .C1(new_n1013), .C2(new_n1018), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1026), .A2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1014), .A2(new_n1016), .A3(new_n995), .ZN(new_n1036));
  INV_X1    g611(.A(G2084), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n840), .A2(KEYINPUT45), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n946), .A2(new_n1039), .A3(new_n995), .ZN(new_n1040));
  INV_X1    g615(.A(G1966), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1036), .A2(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n561), .A2(G8), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT117), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1014), .A2(new_n1016), .A3(new_n1037), .A4(new_n995), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(G8), .A4(new_n561), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1033), .A2(new_n1035), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1033), .A2(new_n1050), .A3(new_n1035), .A4(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1026), .A2(new_n1053), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1019), .A2(new_n1032), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1050), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1027), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT57), .ZN(new_n1062));
  AOI211_X1 g637(.A(new_n1061), .B(new_n1062), .C1(new_n551), .C2(new_n556), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n556), .A2(new_n551), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n1038), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n947), .B1(new_n1068), .B2(new_n945), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT56), .B(G2072), .Z(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1039), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT119), .B(G1956), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1016), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n995), .B1(new_n996), .B2(new_n1015), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1067), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1067), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1078));
  INV_X1    g653(.A(G1348), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n998), .A2(new_n953), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1080), .A2(new_n1081), .B1(new_n607), .B2(new_n608), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1072), .A2(new_n1067), .A3(new_n1076), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1078), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1067), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1077), .A3(KEYINPUT61), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n607), .A2(new_n1091), .A3(new_n608), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1092), .A3(new_n1081), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n609), .A2(KEYINPUT60), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n1081), .A4(new_n609), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1086), .A2(new_n1090), .A3(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n946), .A2(new_n949), .A3(new_n1039), .A4(new_n995), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT58), .B(G1341), .Z(new_n1101));
  AOI22_X1  g676(.A1(new_n1099), .A2(new_n1100), .B1(new_n997), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1069), .A2(KEYINPUT121), .A3(new_n949), .A4(new_n1039), .ZN(new_n1103));
  AOI211_X1 g678(.A(KEYINPUT59), .B(new_n540), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n997), .A2(new_n1101), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1105), .B1(new_n1108), .B2(new_n541), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1083), .B1(new_n1098), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1083), .C1(new_n1098), .C2(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1069), .A2(KEYINPUT53), .A3(new_n755), .A4(new_n1039), .ZN(new_n1116));
  INV_X1    g691(.A(G1961), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1116), .A2(KEYINPUT123), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT123), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1040), .B2(G2078), .ZN(new_n1123));
  AOI21_X1  g698(.A(G301), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(new_n1118), .A3(new_n1116), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1115), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(G301), .B(new_n1123), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1115), .B1(new_n1125), .B2(G171), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1045), .A2(G168), .A3(new_n1046), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G8), .ZN(new_n1132));
  AOI21_X1  g707(.A(G168), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT51), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1131), .A2(new_n1135), .A3(G8), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AND4_X1   g712(.A1(new_n1130), .A2(new_n1033), .A3(new_n1137), .A4(new_n1035), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1112), .A2(new_n1114), .A3(new_n1127), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1060), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1060), .B2(new_n1139), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1124), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1137), .A2(KEYINPUT62), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1141), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(G290), .A2(G1986), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n948), .B1(new_n978), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n965), .A2(new_n1149), .A3(new_n973), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n982), .B1(new_n1147), .B2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(G319), .ZN(new_n1153));
  NOR4_X1   g727(.A1(G229), .A2(G227), .A3(G401), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n871), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1155), .A2(new_n943), .ZN(G308));
  OR2_X1    g730(.A1(new_n1155), .A2(new_n943), .ZN(G225));
endmodule


