//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G20), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT64), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(new_n203), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n213), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT1), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(new_n210), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n221), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n222), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n229), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n214), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n208), .A2(new_n256), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n255), .A2(new_n257), .B1(G150), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n204), .A2(G20), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n253), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n252), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n207), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G50), .B2(new_n263), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n215), .B1(new_n256), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G274), .ZN(new_n273));
  INV_X1    g0073(.A(G45), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(new_n275), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(G226), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G222), .ZN(new_n286));
  INV_X1    g0086(.A(new_n284), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G223), .A3(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n287), .ZN(new_n290));
  AOI211_X1 g0090(.A(new_n277), .B(new_n280), .C1(new_n290), .C2(new_n278), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(G190), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n270), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT68), .B(G179), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n269), .B1(new_n291), .B2(G169), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT17), .ZN(new_n303));
  MUX2_X1   g0103(.A(G223), .B(G226), .S(G1698), .Z(new_n304));
  NAND2_X1  g0104(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n307), .A3(G33), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n308), .A3(new_n281), .ZN(new_n309));
  INV_X1    g0109(.A(G87), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n256), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT73), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n309), .A2(new_n315), .A3(new_n312), .ZN(new_n316));
  AND3_X1   g0116(.A1(new_n314), .A2(new_n278), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G274), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n278), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n275), .ZN(new_n320));
  INV_X1    g0120(.A(new_n279), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n234), .ZN(new_n322));
  OAI21_X1  g0122(.A(G200), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n208), .B1(new_n218), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G159), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n258), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT72), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT72), .B1(new_n325), .B2(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n308), .A2(new_n281), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n208), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G68), .ZN(new_n336));
  AOI21_X1  g0136(.A(G20), .B1(new_n308), .B2(new_n281), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n334), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n332), .B(KEYINPUT16), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT16), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n334), .B1(new_n287), .B2(G20), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n334), .A2(G20), .ZN(new_n342));
  AOI21_X1  g0142(.A(G33), .B1(new_n305), .B2(new_n307), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n203), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n328), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n339), .A2(new_n348), .A3(new_n252), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n272), .B1(new_n313), .B2(KEYINPUT73), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n322), .B1(new_n350), .B2(new_n316), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G190), .ZN(new_n352));
  INV_X1    g0152(.A(new_n265), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n255), .A2(new_n266), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n353), .A2(new_n354), .B1(new_n263), .B2(new_n255), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n323), .A2(new_n349), .A3(new_n352), .A4(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n303), .B1(new_n357), .B2(KEYINPUT74), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n351), .A2(new_n292), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  AOI211_X1 g0160(.A(new_n360), .B(new_n322), .C1(new_n350), .C2(new_n316), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n203), .B1(new_n337), .B2(new_n334), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n282), .A2(G33), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT71), .B(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(G33), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT7), .B1(new_n366), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n363), .A2(new_n367), .B1(new_n330), .B2(new_n331), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n253), .B1(new_n368), .B2(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n355), .B1(new_n369), .B2(new_n348), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n362), .A2(new_n370), .A3(new_n371), .A4(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n349), .A2(new_n356), .ZN(new_n373));
  INV_X1    g0173(.A(new_n322), .ZN(new_n374));
  INV_X1    g0174(.A(new_n297), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n311), .B1(new_n366), .B2(new_n304), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n278), .B1(new_n376), .B2(new_n315), .ZN(new_n377));
  INV_X1    g0177(.A(new_n316), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n374), .B(new_n375), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G169), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n351), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n373), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT18), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT18), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n358), .A2(new_n372), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n285), .A2(G232), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n284), .A2(G107), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT69), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n272), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT69), .A4(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G244), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n320), .B1(new_n321), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(G190), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n266), .A2(G77), .ZN(new_n399));
  OAI22_X1  g0199(.A1(new_n353), .A2(new_n399), .B1(G77), .B2(new_n263), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n255), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n401));
  INV_X1    g0201(.A(new_n257), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT15), .B(G87), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n404), .B2(new_n252), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n396), .B1(new_n392), .B2(new_n393), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n398), .B(new_n405), .C1(new_n292), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n297), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n405), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n406), .B2(G169), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NOR4_X1   g0213(.A1(new_n302), .A2(new_n386), .A3(new_n408), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n264), .A2(new_n203), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n289), .B2(new_n402), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .A3(new_n252), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n418), .B2(new_n252), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT70), .ZN(new_n424));
  AOI22_X1  g0224(.A1(G238), .A2(new_n279), .B1(new_n319), .B2(new_n275), .ZN(new_n425));
  INV_X1    g0225(.A(G1698), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n281), .A2(new_n283), .A3(G226), .A4(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n281), .A2(new_n283), .A3(G232), .A4(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n425), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(G179), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n425), .A2(new_n431), .A3(new_n434), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n434), .B1(new_n425), .B2(new_n431), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n439), .B2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n433), .A2(new_n435), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n424), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n441), .A3(G169), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT70), .A4(new_n436), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n423), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n442), .A2(G200), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n433), .A2(G190), .A3(new_n435), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n449), .A2(new_n423), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n414), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT19), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n257), .A2(new_n456), .A3(G97), .ZN(new_n457));
  NOR2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n310), .B1(new_n429), .B2(new_n208), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n459), .B2(new_n456), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n308), .A2(new_n208), .A3(G68), .A4(new_n281), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n252), .ZN(new_n463));
  INV_X1    g0263(.A(new_n403), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(new_n263), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(KEYINPUT76), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT76), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n253), .B1(new_n460), .B2(new_n461), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n253), .B(new_n263), .C1(G1), .C2(new_n256), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(new_n310), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n207), .A2(G45), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n474), .A2(G250), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n319), .A2(new_n475), .B1(new_n272), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n256), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G238), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n395), .B2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n366), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(new_n272), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n473), .B1(new_n483), .B2(G200), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n471), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT77), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(new_n308), .A3(new_n281), .ZN(new_n488));
  INV_X1    g0288(.A(new_n479), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n272), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n476), .A2(new_n272), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n273), .B2(new_n474), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n471), .A2(KEYINPUT77), .A3(new_n484), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n487), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n472), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n464), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n471), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT75), .ZN(new_n500));
  INV_X1    g0300(.A(new_n490), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n380), .B1(new_n501), .B2(new_n477), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n490), .A2(new_n492), .A3(new_n297), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n483), .A2(G169), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT75), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n499), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g0309(.A1(KEYINPUT5), .A2(G41), .ZN(new_n510));
  NAND2_X1  g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n474), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n278), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n513), .A2(G264), .B1(new_n319), .B2(new_n512), .ZN(new_n514));
  MUX2_X1   g0314(.A(G250), .B(G257), .S(G1698), .Z(new_n515));
  AOI22_X1  g0315(.A1(new_n366), .A2(new_n515), .B1(G33), .B2(G294), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(G190), .C1(new_n272), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n319), .A2(new_n512), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n511), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n475), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n272), .ZN(new_n521));
  INV_X1    g0321(.A(G264), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n515), .A2(new_n308), .A3(new_n281), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G294), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n272), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT25), .B1(new_n264), .B2(new_n529), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n472), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT79), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT22), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(new_n310), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n308), .A2(new_n208), .A3(new_n281), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n208), .A2(G87), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n284), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT23), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n208), .B2(G107), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n529), .A2(KEYINPUT23), .A3(G20), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n542), .A2(new_n543), .B1(new_n479), .B2(new_n208), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n538), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT24), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n538), .A2(new_n540), .A3(new_n547), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n535), .B1(new_n549), .B2(new_n252), .ZN(new_n550));
  AOI211_X1 g0350(.A(KEYINPUT79), .B(new_n253), .C1(new_n546), .C2(new_n548), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n528), .B(new_n534), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n252), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT79), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n549), .A2(new_n535), .A3(new_n252), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n533), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n523), .A2(new_n526), .ZN(new_n557));
  INV_X1    g0357(.A(G179), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(G169), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n552), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G283), .ZN(new_n563));
  INV_X1    g0363(.A(G97), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n563), .B(new_n208), .C1(G33), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n478), .A2(G20), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n252), .A3(new_n566), .ZN(new_n567));
  OR3_X1    g0367(.A1(new_n567), .A2(KEYINPUT78), .A3(KEYINPUT20), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n265), .B(G116), .C1(G1), .C2(new_n256), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n264), .A2(new_n478), .ZN(new_n570));
  XOR2_X1   g0370(.A(KEYINPUT78), .B(KEYINPUT20), .Z(new_n571));
  NAND2_X1  g0371(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n520), .A2(G270), .A3(new_n272), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G257), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n522), .B2(G1698), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n366), .A2(new_n576), .B1(G303), .B2(new_n284), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n518), .B(new_n574), .C1(new_n577), .C2(new_n272), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n573), .B1(new_n578), .B2(G200), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n360), .B2(new_n578), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n366), .A2(new_n576), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n284), .A2(G303), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n272), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n574), .A2(new_n518), .ZN(new_n585));
  OAI21_X1  g0385(.A(G169), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n570), .B1(new_n472), .B2(new_n478), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n567), .A2(KEYINPUT78), .A3(KEYINPUT20), .ZN(new_n588));
  INV_X1    g0388(.A(new_n572), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n581), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n584), .A2(new_n585), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G179), .A3(new_n573), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n573), .A2(new_n578), .A3(KEYINPUT21), .A4(G169), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n580), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n529), .B1(new_n341), .B2(new_n345), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n597), .A2(new_n564), .A3(G107), .ZN(new_n598));
  XNOR2_X1  g0398(.A(G97), .B(G107), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n600), .A2(new_n208), .B1(new_n289), .B2(new_n258), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n252), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n264), .A2(new_n564), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n497), .A2(G97), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n395), .A2(G1698), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT4), .B1(new_n366), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(KEYINPUT4), .A2(G244), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n281), .A2(new_n283), .A3(new_n608), .A4(new_n426), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n281), .A2(new_n283), .A3(G250), .A4(G1698), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n563), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n278), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n513), .A2(G257), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n518), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(G190), .A3(new_n518), .A4(new_n613), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n605), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n380), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(new_n297), .A3(new_n518), .A4(new_n613), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n595), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n455), .A2(new_n509), .A3(new_n562), .A4(new_n623), .ZN(G372));
  AOI22_X1  g0424(.A1(new_n471), .A2(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT80), .ZN(new_n626));
  INV_X1    g0426(.A(new_n473), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n471), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g0428(.A(KEYINPUT80), .B(new_n473), .C1(new_n467), .C2(new_n470), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n483), .A2(G200), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n494), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n552), .A2(new_n617), .A3(new_n621), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n556), .B2(new_n560), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n495), .A2(new_n494), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT77), .B1(new_n471), .B2(new_n484), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n638), .B(new_n508), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n625), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT76), .B1(new_n463), .B2(new_n466), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n469), .A2(new_n468), .A3(new_n465), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n627), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT80), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n471), .A2(new_n626), .A3(new_n627), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n632), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n638), .A4(new_n643), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n637), .A2(new_n642), .A3(new_n643), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n455), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT81), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n373), .A2(new_n381), .A3(new_n384), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n384), .B1(new_n373), .B2(new_n381), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n383), .A2(KEYINPUT81), .A3(new_n385), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n448), .B1(new_n451), .B2(new_n413), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n358), .B(new_n372), .C1(new_n660), .C2(KEYINPUT82), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n660), .A2(KEYINPUT82), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n300), .B1(new_n663), .B2(new_n296), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n653), .A2(new_n664), .ZN(G369));
  INV_X1    g0465(.A(new_n635), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT83), .Z(new_n669));
  INV_X1    g0469(.A(G213), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n670), .B1(new_n667), .B2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n590), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n666), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n595), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n679), .A2(KEYINPUT84), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(KEYINPUT84), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n556), .A2(new_n560), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n556), .A2(new_n675), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n683), .A2(new_n675), .B1(new_n561), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n683), .A2(new_n674), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n635), .A2(new_n674), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n562), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(G399));
  NAND2_X1  g0490(.A1(new_n211), .A2(new_n271), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n207), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n458), .A2(new_n310), .A3(new_n478), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n693), .A2(new_n695), .B1(new_n220), .B2(new_n692), .ZN(new_n696));
  XNOR2_X1  g0496(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n652), .A2(new_n675), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n650), .B1(new_n633), .B2(new_n638), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n643), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT87), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n649), .A2(new_n638), .A3(new_n643), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT87), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n496), .A2(new_n650), .A3(new_n508), .A4(new_n638), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n643), .A4(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n703), .A2(new_n637), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n675), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n700), .B1(new_n710), .B2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n557), .A2(new_n493), .A3(new_n612), .A4(new_n613), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n592), .A2(G179), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n483), .A2(new_n526), .A3(new_n523), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n578), .A2(new_n558), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n612), .A2(new_n613), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n716), .A2(new_n717), .A3(new_n718), .A4(KEYINPUT30), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n557), .A2(new_n375), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n483), .A3(new_n614), .A4(new_n578), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT86), .A3(new_n674), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT86), .B1(new_n722), .B2(new_n674), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n725), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT31), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(new_n723), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n509), .A2(new_n562), .A3(new_n623), .A4(new_n675), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n711), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n698), .B1(new_n733), .B2(G1), .ZN(G364));
  INV_X1    g0534(.A(G13), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G45), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT88), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n693), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n678), .B2(G330), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n682), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT89), .Z(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n678), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n215), .B1(new_n208), .B2(G169), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n749), .A2(KEYINPUT90), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(KEYINPUT90), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n297), .A2(new_n208), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT93), .Z(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n208), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n757), .A2(G326), .B1(G294), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n208), .A2(G179), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n287), .B1(new_n766), .B2(G329), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n754), .A2(new_n764), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n360), .A3(G200), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(KEYINPUT92), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n360), .A2(G200), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n754), .A2(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n774), .A2(G283), .B1(G322), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT95), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n754), .A2(new_n360), .A3(G200), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n770), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n761), .A2(KEYINPUT94), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n762), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n776), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n789), .A2(new_n202), .B1(new_n289), .B2(new_n768), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G107), .B2(new_n774), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n759), .A2(new_n564), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n765), .A2(new_n326), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT91), .B(KEYINPUT32), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n287), .B1(new_n779), .B2(new_n310), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n792), .B(new_n796), .C1(new_n793), .C2(new_n795), .ZN(new_n797));
  INV_X1    g0597(.A(new_n755), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G50), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n784), .A2(G68), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n791), .A2(new_n797), .A3(new_n799), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n753), .B1(new_n788), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n739), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n211), .A2(new_n287), .ZN(new_n804));
  INV_X1    g0604(.A(G355), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(G116), .B2(new_n211), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n249), .A2(new_n274), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n211), .A2(new_n333), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n274), .B2(new_n220), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n752), .A2(new_n745), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n803), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n748), .A2(new_n802), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n742), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n753), .A2(new_n744), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n803), .B1(new_n817), .B2(G77), .ZN(new_n818));
  INV_X1    g0618(.A(new_n768), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  XNOR2_X1  g0621(.A(KEYINPUT97), .B(G143), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n783), .C1(new_n789), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G137), .B2(new_n798), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT34), .Z(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n366), .B1(new_n826), .B2(new_n765), .C1(new_n202), .C2(new_n759), .ZN(new_n827));
  INV_X1    g0627(.A(new_n774), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n203), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n827), .B(new_n829), .C1(G50), .C2(new_n780), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n798), .A2(G303), .B1(new_n819), .B2(G116), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n783), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT96), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n776), .A2(G294), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n287), .B(new_n792), .C1(G311), .C2(new_n766), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G87), .A2(new_n774), .B1(new_n780), .B2(G107), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n835), .A2(new_n836), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n818), .B1(new_n840), .B2(new_n752), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n675), .A2(new_n405), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n394), .A2(new_n397), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n405), .B1(new_n844), .B2(new_n380), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n407), .A2(new_n843), .B1(new_n845), .B2(new_n409), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n410), .A2(new_n412), .A3(new_n674), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT98), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT98), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n845), .A2(new_n409), .A3(new_n675), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n411), .B1(new_n406), .B2(G190), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n844), .A2(G200), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n842), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n849), .B(new_n850), .C1(new_n853), .C2(new_n413), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n841), .B1(new_n855), .B2(new_n744), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT99), .Z(new_n857));
  XNOR2_X1  g0657(.A(new_n699), .B(new_n855), .ZN(new_n858));
  INV_X1    g0658(.A(new_n732), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n803), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n860), .A2(KEYINPUT100), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(new_n860), .B2(KEYINPUT100), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n857), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n736), .A2(new_n207), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n722), .A2(new_n674), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n728), .A2(KEYINPUT101), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n730), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n455), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT102), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n332), .B1(new_n336), .B2(new_n338), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n340), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n355), .B1(new_n369), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n672), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n386), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n357), .B1(new_n672), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g0678(.A(G169), .B1(new_n317), .B2(new_n322), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n875), .B1(new_n379), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT37), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n672), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n373), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n382), .A2(new_n883), .A3(new_n357), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n877), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n657), .A2(new_n658), .A3(new_n358), .A4(new_n372), .ZN(new_n888));
  INV_X1    g0688(.A(new_n883), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n382), .A2(new_n883), .A3(new_n357), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n885), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n887), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n675), .A2(new_n423), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n444), .A2(new_n447), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n451), .B(new_n898), .C1(new_n899), .C2(new_n423), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n897), .B1(new_n448), .B2(new_n452), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(new_n870), .A3(new_n855), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT40), .B1(new_n896), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n902), .A2(new_n870), .A3(new_n855), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n877), .A2(new_n886), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n895), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n877), .A2(new_n886), .A3(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n904), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n872), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n872), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(G330), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT103), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI22_X1  g0717(.A1(new_n888), .A2(new_n889), .B1(new_n885), .B2(new_n892), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n908), .B1(new_n918), .B2(KEYINPUT38), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n448), .A2(new_n675), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n659), .A2(new_n882), .ZN(new_n926));
  INV_X1    g0726(.A(new_n902), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n652), .A2(new_n855), .A3(new_n675), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n850), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n926), .B1(new_n929), .B2(new_n909), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n664), .B1(new_n454), .B2(new_n711), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n866), .B1(new_n917), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n917), .B2(new_n933), .ZN(new_n935));
  INV_X1    g0735(.A(new_n600), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n936), .A2(KEYINPUT35), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(KEYINPUT35), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n937), .A2(G116), .A3(new_n217), .A4(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT36), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n220), .A2(G77), .A3(new_n324), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(G50), .B2(new_n203), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(G1), .A3(new_n735), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n935), .A2(new_n940), .A3(new_n943), .ZN(G367));
  OAI211_X1 g0744(.A(new_n617), .B(new_n621), .C1(new_n605), .C2(new_n675), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n638), .A2(new_n674), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n562), .A3(new_n688), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n621), .B1(new_n683), .B2(new_n945), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(KEYINPUT42), .B1(new_n949), .B2(new_n675), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT42), .B2(new_n948), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n674), .B1(new_n628), .B2(new_n629), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n633), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n643), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g0759(.A(new_n686), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n947), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n691), .B(KEYINPUT41), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n687), .A2(new_n689), .ZN(new_n964));
  INV_X1    g0764(.A(new_n947), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT44), .Z(new_n967));
  NOR2_X1   g0767(.A1(new_n964), .A2(new_n965), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n686), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n689), .B1(new_n685), .B2(new_n688), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n682), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n733), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT104), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n733), .A2(KEYINPUT104), .A3(new_n973), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n963), .B1(new_n978), .B2(new_n733), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n738), .A2(G1), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n962), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n811), .B1(new_n211), .B2(new_n403), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n240), .A2(new_n808), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n803), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT105), .B(KEYINPUT46), .Z(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n779), .B2(new_n478), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n529), .B2(new_n759), .C1(new_n789), .C2(new_n778), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n780), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n833), .B2(new_n768), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G294), .C2(new_n784), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n774), .A2(G97), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n366), .B1(G317), .B2(new_n766), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT106), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n994), .C1(new_n769), .C2(new_n756), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n284), .B1(new_n766), .B2(G137), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n202), .B2(new_n779), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n828), .A2(new_n289), .B1(new_n821), .B2(new_n789), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G68), .C2(new_n760), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n756), .B2(new_n822), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n783), .A2(new_n326), .B1(new_n768), .B2(new_n201), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT107), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n995), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n753), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n984), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n746), .B2(new_n955), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n981), .A2(new_n1008), .ZN(G387));
  OR2_X1    g0809(.A1(new_n685), .A2(new_n746), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n804), .A2(new_n695), .B1(G107), .B2(new_n211), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n237), .A2(new_n274), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n254), .A2(G50), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT50), .ZN(new_n1014));
  AOI211_X1 g0814(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n808), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1011), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n803), .B1(new_n1017), .B2(new_n812), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n760), .A2(new_n464), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n789), .B2(new_n201), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT109), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n779), .A2(new_n289), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G150), .B2(new_n766), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n991), .A2(new_n366), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G68), .B2(new_n819), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G159), .A2(new_n798), .B1(new_n784), .B2(new_n255), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G303), .A2(new_n819), .B1(new_n776), .B2(G317), .ZN(new_n1028));
  INV_X1    g0828(.A(G322), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1028), .B1(new_n769), .B2(new_n783), .C1(new_n756), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(G294), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n759), .A2(new_n833), .B1(new_n779), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n366), .B1(G326), .B2(new_n766), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n478), .C2(new_n828), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT49), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1027), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1018), .B1(new_n1040), .B2(new_n752), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n973), .A2(new_n980), .B1(new_n1010), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n974), .A2(new_n692), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n733), .A2(new_n973), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1042), .B1(new_n1043), .B2(new_n1044), .ZN(G393));
  XNOR2_X1  g0845(.A(new_n970), .B(new_n960), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n691), .B1(new_n1046), .B2(new_n974), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(new_n978), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n246), .A2(new_n808), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n811), .B1(new_n564), .B2(new_n211), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n803), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n284), .B1(new_n765), .B2(new_n1029), .C1(new_n779), .C2(new_n833), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n798), .A2(G317), .B1(new_n776), .B2(G311), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT52), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(G107), .C2(new_n774), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n819), .A2(G294), .B1(G116), .B2(new_n760), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n778), .B2(new_n783), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT110), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n789), .A2(new_n326), .B1(new_n821), .B2(new_n755), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n759), .A2(new_n289), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n779), .A2(new_n203), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n765), .A2(new_n822), .ZN(new_n1063));
  OR4_X1    g0863(.A1(new_n333), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n828), .A2(new_n310), .B1(new_n768), .B2(new_n254), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(G50), .C2(new_n784), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1055), .A2(new_n1058), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT111), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n753), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1051), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n746), .B2(new_n947), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n980), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1072), .B1(new_n1046), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1048), .A2(new_n1074), .ZN(G390));
  INV_X1    g0875(.A(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n870), .A2(G330), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n855), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n927), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n731), .A2(new_n902), .A3(G330), .A4(new_n855), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n709), .A2(new_n675), .A3(new_n855), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n850), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1076), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n633), .A2(new_n636), .A3(new_n634), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n705), .A2(new_n643), .A3(new_n707), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(KEYINPUT87), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n674), .B1(new_n1087), .B2(new_n708), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n847), .B1(new_n1088), .B2(new_n855), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1089), .A2(KEYINPUT112), .A3(new_n1080), .A4(new_n1079), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n902), .A2(new_n855), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n1077), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n927), .B1(new_n732), .B2(new_n1078), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n928), .A2(new_n850), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n454), .A2(new_n1077), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n664), .C1(new_n454), .C2(new_n711), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1097), .A2(new_n902), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n921), .A2(new_n924), .B1(new_n1105), .B2(new_n922), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT38), .B1(new_n890), .B2(new_n893), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n922), .B1(new_n1107), .B2(new_n887), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1083), .B2(new_n902), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1093), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1108), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n1089), .B2(new_n927), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n924), .B1(new_n896), .B2(KEYINPUT39), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1105), .A2(new_n922), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1115), .A3(new_n1080), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1110), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1104), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1099), .A2(new_n1103), .A3(new_n1116), .A4(new_n1110), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n692), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n284), .B1(new_n765), .B2(new_n1033), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n829), .A2(new_n1061), .A3(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n529), .B2(new_n783), .C1(new_n833), .C2(new_n755), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n780), .A2(G87), .B1(G116), .B2(new_n776), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n564), .B2(new_n768), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n779), .A2(new_n821), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1127), .B1(new_n768), .B2(new_n1128), .C1(new_n828), .C2(new_n201), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n798), .A2(G128), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n784), .A2(G137), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n776), .A2(G132), .ZN(new_n1132));
  INV_X1    g0932(.A(G125), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n287), .B1(new_n1133), .B2(new_n765), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G159), .B2(new_n760), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1123), .A2(new_n1125), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n752), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1138), .B(new_n803), .C1(new_n255), .C2(new_n817), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(new_n1113), .B2(new_n743), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT113), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1140), .B(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT114), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1110), .A2(new_n1116), .A3(new_n980), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1120), .B1(new_n1145), .B2(new_n1146), .ZN(G378));
  AOI21_X1  g0947(.A(new_n910), .B1(new_n905), .B2(new_n919), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n902), .A2(new_n870), .A3(new_n910), .A4(new_n855), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n908), .B2(new_n907), .ZN(new_n1150));
  OAI21_X1  g0950(.A(G330), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n302), .A2(new_n269), .A3(new_n882), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n269), .A2(new_n882), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n296), .A2(new_n301), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT118), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n925), .B2(new_n930), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G330), .B(new_n1160), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1164), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1073), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n803), .B1(new_n817), .B2(G50), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1160), .A2(new_n744), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n366), .A2(G41), .ZN(new_n1171));
  AOI211_X1 g0971(.A(G50), .B(new_n1171), .C1(new_n256), .C2(new_n271), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n776), .A2(G107), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT115), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n774), .A2(G58), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n765), .A2(new_n833), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1176), .B(new_n1022), .C1(G68), .C2(new_n760), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n819), .A2(new_n464), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .A4(new_n1171), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n564), .A2(new_n783), .B1(new_n755), .B2(new_n478), .ZN(new_n1180));
  NOR3_X1   g0980(.A1(new_n1174), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT116), .ZN(new_n1182));
  XOR2_X1   g0982(.A(new_n1182), .B(KEYINPUT58), .Z(new_n1183));
  NAND2_X1  g0983(.A1(new_n819), .A2(G137), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n821), .B2(new_n759), .C1(new_n779), .C2(new_n1128), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G128), .B2(new_n776), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1186), .B1(new_n1133), .B2(new_n755), .C1(new_n826), .C2(new_n783), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n774), .A2(G159), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n1187), .B2(KEYINPUT59), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1172), .B(new_n1183), .C1(new_n1188), .C2(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT117), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n753), .B1(new_n1193), .B2(KEYINPUT117), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1169), .B(new_n1170), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1168), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1160), .B1(new_n912), .B2(G330), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1165), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n931), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1162), .A2(new_n925), .A3(new_n930), .A4(new_n1165), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1084), .A2(new_n1090), .B1(new_n1097), .B2(new_n1096), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1103), .B1(new_n1117), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1204), .A3(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n692), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1204), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1197), .B1(new_n1206), .B2(new_n1208), .ZN(G375));
  INV_X1    g1009(.A(new_n963), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1203), .A2(new_n1102), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1104), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n803), .B1(new_n817), .B2(G68), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n781), .A2(new_n564), .B1(new_n833), .B2(new_n789), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n287), .B1(new_n766), .B2(G303), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1019), .B(new_n1215), .C1(new_n828), .C2(new_n289), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G294), .C2(new_n798), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n783), .A2(new_n478), .B1(new_n768), .B2(new_n529), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT120), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(KEYINPUT120), .B2(new_n1218), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(KEYINPUT121), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n333), .B1(G128), .B2(new_n766), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n201), .B2(new_n759), .C1(new_n783), .C2(new_n1128), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G132), .B2(new_n798), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n776), .A2(G137), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n780), .A2(G159), .B1(G150), .B2(new_n819), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n1175), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1222), .A2(KEYINPUT121), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1223), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1213), .B1(new_n1231), .B2(new_n752), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n927), .A2(new_n743), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n980), .B(KEYINPUT119), .Z(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1203), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1212), .A2(new_n1237), .ZN(G381));
  OR3_X1    g1038(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT122), .ZN(new_n1241));
  INV_X1    g1041(.A(G375), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1120), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1241), .A2(new_n1247), .ZN(G407));
  OAI211_X1 g1048(.A(G407), .B(G213), .C1(G343), .C2(new_n1247), .ZN(G409));
  NAND2_X1  g1049(.A1(new_n673), .A2(G213), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1102), .A2(new_n1091), .A3(KEYINPUT60), .A4(new_n1098), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(new_n692), .ZN(new_n1253));
  OAI21_X1  g1053(.A(KEYINPUT60), .B1(new_n1203), .B2(new_n1102), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1211), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(G384), .B1(new_n1256), .B2(new_n1237), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1236), .B(new_n864), .C1(new_n1253), .C2(new_n1255), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1252), .A2(new_n692), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1211), .B2(new_n1254), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n864), .B1(new_n1261), .B2(new_n1236), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1256), .A2(G384), .A3(new_n1237), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1259), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1080), .ZN(new_n1267));
  NOR3_X1   g1067(.A1(new_n1106), .A2(new_n1109), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1094), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1102), .B1(new_n1270), .B2(new_n1099), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1164), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1162), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1210), .A3(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1266), .B1(new_n1271), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1207), .A2(new_n1204), .A3(KEYINPUT124), .A4(new_n1210), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1235), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1196), .B1(new_n1202), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1246), .ZN(new_n1282));
  OAI211_X1 g1082(.A(G378), .B(new_n1197), .C1(new_n1206), .C2(new_n1208), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1281), .B1(new_n1280), .B2(new_n1246), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1250), .B(new_n1265), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1280), .A2(new_n1246), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT125), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1291), .A2(KEYINPUT62), .A3(new_n1250), .A4(new_n1265), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1288), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1250), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n673), .A2(G213), .A3(G2897), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(new_n1265), .B2(new_n1295), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1293), .A2(new_n1298), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1048), .A2(new_n1074), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G387), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G390), .A2(new_n981), .A3(new_n1008), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n815), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1301), .A2(new_n1304), .A3(new_n1302), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(KEYINPUT127), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1299), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1311), .B2(new_n1286), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1312), .B(new_n1298), .C1(new_n1311), .C2(new_n1286), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1310), .A2(new_n1313), .ZN(G405));
  INV_X1    g1114(.A(new_n1246), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1283), .B1(new_n1242), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1265), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1308), .ZN(G402));
endmodule


