//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(G237), .A2(G953), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(G143), .A3(G214), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n193), .A2(new_n194), .ZN(new_n200));
  AOI21_X1  g014(.A(G143), .B1(new_n196), .B2(G214), .ZN(new_n201));
  OAI211_X1 g015(.A(KEYINPUT18), .B(G131), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT77), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n203), .A2(new_n204), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n199), .B(new_n202), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n200), .B2(new_n201), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT17), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT16), .ZN(new_n213));
  INV_X1    g027(.A(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G125), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G140), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(G146), .B(new_n215), .C1(new_n219), .C2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n222));
  AOI21_X1  g036(.A(G146), .B1(new_n222), .B2(new_n215), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  AOI211_X1 g038(.A(KEYINPUT74), .B(G146), .C1(new_n222), .C2(new_n215), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n212), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n195), .A2(new_n227), .A3(new_n197), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n210), .A2(new_n211), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT94), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT94), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n210), .A2(new_n228), .A3(new_n231), .A4(new_n211), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n190), .B(new_n209), .C1(new_n226), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n215), .B1(new_n219), .B2(new_n213), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n204), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT74), .A3(new_n220), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n221), .A2(new_n223), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n240), .A2(new_n212), .A3(new_n230), .A4(new_n232), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n190), .B1(new_n241), .B2(new_n209), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n187), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT95), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT95), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n187), .C1(new_n235), .C2(new_n242), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(G475), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G475), .A2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n210), .A2(new_n228), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n250));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(new_n203), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT92), .B1(new_n219), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT19), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n203), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AND3_X1   g071(.A1(new_n257), .A2(KEYINPUT93), .A3(new_n204), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT93), .B1(new_n257), .B2(new_n204), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n220), .B(new_n249), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n190), .B1(new_n260), .B2(new_n209), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n248), .B1(new_n261), .B2(new_n235), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT20), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n248), .C1(new_n261), .C2(new_n235), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n247), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n192), .A2(G952), .ZN(new_n268));
  INV_X1    g082(.A(G234), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n191), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT72), .B(G902), .Z(new_n272));
  AOI211_X1 g086(.A(new_n192), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT21), .B(G898), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT9), .B(G234), .ZN(new_n276));
  INV_X1    g090(.A(G217), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(G953), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT96), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(G122), .ZN(new_n281));
  INV_X1    g095(.A(G122), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT96), .A3(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n280), .A2(G122), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(KEYINPUT98), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(KEYINPUT14), .B2(new_n285), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n281), .A2(new_n283), .B1(new_n285), .B2(KEYINPUT14), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT98), .ZN(new_n290));
  OAI21_X1  g104(.A(G107), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT78), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G107), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n296), .A2(new_n284), .A3(KEYINPUT97), .A4(new_n285), .ZN(new_n297));
  XNOR2_X1  g111(.A(G128), .B(G143), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n298), .B(G134), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT97), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(new_n284), .A3(new_n285), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n291), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n298), .A2(G134), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(G134), .ZN(new_n305));
  INV_X1    g119(.A(G128), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G143), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G134), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n304), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n298), .A2(new_n308), .A3(G134), .A4(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(new_n301), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n296), .B1(new_n284), .B2(new_n285), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n310), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n278), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n301), .A2(new_n300), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n304), .A3(new_n305), .A4(new_n297), .ZN(new_n317));
  OR2_X1    g131(.A1(new_n289), .A2(KEYINPUT98), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n289), .B2(KEYINPUT98), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n292), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n314), .B(new_n278), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n272), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT99), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G478), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT15), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n314), .B1(new_n317), .B2(new_n321), .ZN(new_n329));
  INV_X1    g143(.A(new_n278), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n322), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT99), .A3(new_n272), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n324), .A2(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n267), .A2(new_n275), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT2), .B(G113), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n338), .B(KEYINPUT68), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G119), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n346), .A3(G116), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G113), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n350), .A2(new_n293), .A3(new_n295), .A4(new_n351), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n350), .A2(new_n293), .A3(new_n295), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n189), .A2(G107), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n352), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT81), .B(G101), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n292), .A2(G104), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n292), .A2(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n296), .B2(G104), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G101), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  OR2_X1    g179(.A1(new_n349), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(KEYINPUT4), .ZN(new_n367));
  INV_X1    g181(.A(new_n359), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n357), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT80), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT80), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n357), .A2(new_n371), .A3(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n367), .B1(new_n373), .B2(G101), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n357), .B2(new_n368), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n350), .A2(new_n293), .A3(new_n295), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n351), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT80), .B(new_n359), .C1(new_n380), .C2(new_n352), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n376), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n343), .A2(new_n340), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n342), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n366), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G110), .B(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n366), .B(new_n387), .C1(new_n374), .C2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n392), .A3(new_n388), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT0), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n306), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n204), .A2(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n194), .A2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n306), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT64), .B1(new_n194), .B2(G146), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n204), .A3(G143), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n396), .A2(new_n403), .A3(new_n405), .A4(new_n399), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n394), .B1(new_n407), .B2(new_n217), .ZN(new_n408));
  OR2_X1    g222(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n306), .B1(new_n411), .B2(new_n398), .ZN(new_n412));
  XNOR2_X1  g226(.A(G143), .B(G146), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n405), .A3(new_n399), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n409), .A2(G128), .A3(new_n410), .ZN(new_n415));
  OAI22_X1  g229(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  MUX2_X1   g230(.A(new_n407), .B(new_n416), .S(new_n217), .Z(new_n417));
  OAI21_X1  g231(.A(new_n408), .B1(new_n417), .B2(new_n394), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT88), .B(G224), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n192), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT89), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n418), .B(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n391), .A2(new_n393), .A3(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n357), .A2(new_n360), .B1(new_n363), .B2(G101), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n349), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n387), .B(KEYINPUT8), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n348), .B1(KEYINPUT5), .B2(new_n338), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n341), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n365), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT7), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n426), .A2(new_n430), .B1(new_n417), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n418), .A2(new_n422), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(KEYINPUT7), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n390), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n424), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n424), .A2(new_n438), .A3(new_n436), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(KEYINPUT90), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n438), .B1(new_n424), .B2(new_n436), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND4_X1   g260(.A1(new_n337), .A2(new_n442), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n306), .A2(G119), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n346), .A2(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT24), .B(G110), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT73), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT23), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n456));
  OAI211_X1 g270(.A(G119), .B(new_n306), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n449), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n452), .B1(new_n459), .B2(G110), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n238), .A3(new_n239), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT75), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n238), .A2(new_n460), .A3(new_n239), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n207), .ZN(new_n466));
  INV_X1    g280(.A(G110), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n457), .A2(new_n467), .A3(new_n449), .A4(new_n458), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n450), .A2(new_n451), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n220), .B(new_n466), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT22), .B(G137), .ZN(new_n474));
  INV_X1    g288(.A(G221), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(new_n269), .A3(G953), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n474), .B(new_n476), .Z(new_n477));
  AND3_X1   g291(.A1(new_n465), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n465), .B2(new_n473), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(KEYINPUT25), .A3(new_n272), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n465), .A2(new_n473), .ZN(new_n482));
  INV_X1    g296(.A(new_n477), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n465), .A2(new_n473), .A3(new_n477), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n484), .A2(new_n272), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT25), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n277), .B1(new_n272), .B2(G234), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n480), .ZN(new_n494));
  OAI22_X1  g308(.A1(new_n489), .A2(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n341), .B1(new_n343), .B2(new_n340), .ZN(new_n496));
  INV_X1    g310(.A(G137), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G134), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(KEYINPUT11), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(KEYINPUT11), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n497), .A2(G134), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(KEYINPUT11), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n506), .A3(new_n227), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n498), .A2(KEYINPUT66), .ZN(new_n508));
  INV_X1    g322(.A(new_n504), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n497), .A3(G134), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G131), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n414), .A2(new_n415), .ZN(new_n514));
  AND2_X1   g328(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n515));
  NOR2_X1   g329(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n398), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n413), .B1(new_n517), .B2(G128), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n507), .B(new_n513), .C1(new_n514), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n402), .A2(new_n406), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n498), .A2(new_n505), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n522), .B(new_n509), .C1(new_n523), .C2(new_n498), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G131), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n525), .B2(new_n507), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT30), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n524), .A2(G131), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n227), .B1(new_n503), .B2(new_n506), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n407), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n519), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n496), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n496), .A3(new_n519), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n196), .A2(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT27), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n539), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT69), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n520), .A2(new_n526), .A3(KEYINPUT30), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n531), .B1(new_n530), .B2(new_n519), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n384), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n534), .A2(new_n535), .A3(new_n539), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n545), .A3(new_n543), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT70), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n545), .A3(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(new_n534), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n496), .B1(new_n530), .B2(new_n519), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT28), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n534), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n539), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n554), .A2(KEYINPUT31), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n564), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n553), .B2(new_n562), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n557), .A2(KEYINPUT29), .A3(new_n539), .A4(new_n559), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(new_n272), .ZN(new_n571));
  INV_X1    g385(.A(new_n556), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n558), .B1(new_n572), .B2(new_n534), .ZN(new_n573));
  INV_X1    g387(.A(new_n559), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT71), .B1(new_n575), .B2(new_n539), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n557), .A2(KEYINPUT71), .A3(new_n539), .A4(new_n559), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n561), .B1(new_n533), .B2(new_n555), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT29), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n571), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n569), .A2(KEYINPUT32), .B1(new_n581), .B2(G472), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n495), .B1(new_n567), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n375), .B1(new_n370), .B2(new_n372), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n407), .B(new_n382), .C1(new_n584), .C2(new_n367), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n361), .A2(new_n416), .A3(KEYINPUT10), .A4(new_n364), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT84), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n514), .A2(new_n518), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT84), .A3(new_n425), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n514), .A2(KEYINPUT82), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n194), .A2(G146), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT1), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT83), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT83), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n398), .A2(new_n597), .A3(KEYINPUT1), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(G128), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n414), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT82), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n414), .B2(new_n415), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n593), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n425), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n588), .A2(new_n592), .B1(new_n590), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n528), .A2(new_n529), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n585), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G140), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n192), .A2(G227), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n606), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n382), .A2(new_n407), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n374), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n604), .A2(new_n590), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n586), .A2(new_n587), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT84), .B1(new_n591), .B2(new_n425), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n613), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n365), .A2(new_n589), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n604), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n613), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT12), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(KEYINPUT12), .A3(new_n613), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n607), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n610), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n621), .A2(new_n630), .A3(G469), .ZN(new_n631));
  NAND2_X1  g445(.A1(G469), .A2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n272), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n585), .A2(new_n605), .A3(new_n606), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n606), .B1(new_n585), .B2(new_n605), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n610), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(KEYINPUT85), .B1(new_n612), .B2(new_n628), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT85), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n610), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n634), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(G469), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n633), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n276), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n475), .B1(new_n644), .B2(new_n187), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT86), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n628), .A2(new_n611), .A3(new_n607), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n611), .B1(new_n620), .B2(new_n607), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  INV_X1    g463(.A(new_n640), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n642), .B(new_n272), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n620), .A2(new_n612), .B1(new_n629), .B2(new_n610), .ZN(new_n652));
  OAI21_X1  g466(.A(G469), .B1(new_n652), .B2(G902), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n645), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n447), .A2(new_n583), .A3(new_n646), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n358), .ZN(G3));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n655), .ZN(new_n659));
  AOI211_X1 g473(.A(KEYINPUT86), .B(new_n645), .C1(new_n651), .C2(new_n653), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G472), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n634), .B1(new_n553), .B2(new_n562), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n565), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n495), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n424), .A2(new_n438), .A3(new_n436), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n443), .B1(new_n667), .B2(new_n444), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n275), .ZN(new_n671));
  OAI211_X1 g485(.A(KEYINPUT100), .B(new_n443), .C1(new_n667), .C2(new_n444), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT33), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n331), .B2(KEYINPUT101), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n332), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n634), .A2(new_n327), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n326), .A2(new_n327), .A3(new_n333), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n676), .B1(new_n675), .B2(new_n677), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n267), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n670), .A2(new_n671), .A3(new_n672), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n666), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT34), .B(G104), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G6));
  NOR2_X1   g503(.A1(new_n267), .A2(new_n275), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n670), .A2(new_n690), .A3(new_n336), .A4(new_n672), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n666), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  AOI21_X1  g509(.A(new_n491), .B1(new_n481), .B2(new_n488), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n483), .A2(KEYINPUT36), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n482), .B(new_n697), .Z(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n493), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n664), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n447), .A2(new_n646), .A3(new_n656), .A4(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT103), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n702), .B(new_n704), .ZN(G12));
  AOI21_X1  g519(.A(new_n700), .B1(new_n582), .B2(new_n567), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n670), .A2(new_n706), .A3(new_n672), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n273), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(KEYINPUT104), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n710), .A2(new_n270), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n247), .A2(new_n266), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n336), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n661), .A2(new_n707), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XOR2_X1   g532(.A(new_n712), .B(KEYINPUT39), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n661), .A2(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT40), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT40), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n696), .A2(new_n699), .ZN(new_n723));
  INV_X1    g537(.A(new_n443), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n723), .A2(new_n683), .A3(new_n715), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n563), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n572), .A2(new_n534), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n561), .ZN(new_n730));
  AOI21_X1  g544(.A(G902), .B1(new_n554), .B2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n567), .B(new_n728), .C1(new_n662), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n442), .A2(new_n446), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT38), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n725), .A2(new_n726), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n721), .A2(new_n722), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT106), .B(G143), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G45));
  NAND2_X1  g554(.A1(new_n675), .A2(new_n677), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT102), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n679), .A3(new_n678), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n267), .A3(new_n713), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n661), .A2(new_n707), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G146), .ZN(G48));
  OAI21_X1  g561(.A(new_n272), .B1(new_n649), .B2(new_n650), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n642), .A2(KEYINPUT107), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI221_X1 g564(.A(new_n272), .B1(KEYINPUT107), .B2(new_n642), .C1(new_n649), .C2(new_n650), .ZN(new_n751));
  INV_X1    g565(.A(new_n645), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n696), .B1(new_n492), .B2(new_n480), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n581), .A2(G472), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n728), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n569), .A2(KEYINPUT32), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n686), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND4_X1  g576(.A1(new_n583), .A2(new_n752), .A3(new_n751), .A4(new_n750), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n691), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n280), .ZN(G18));
  NAND3_X1  g579(.A1(new_n670), .A2(new_n706), .A3(new_n672), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n750), .A2(new_n751), .A3(new_n752), .A4(new_n337), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G119), .ZN(G21));
  AND4_X1   g583(.A1(new_n267), .A2(new_n670), .A3(new_n336), .A4(new_n672), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT108), .B1(new_n664), .B2(new_n495), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n560), .A2(new_n561), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n546), .B2(new_n552), .ZN(new_n776));
  OAI21_X1  g590(.A(G472), .B1(new_n776), .B2(new_n634), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n754), .A2(new_n772), .A3(new_n565), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n753), .A2(new_n275), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n770), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  AND2_X1   g596(.A1(new_n668), .A2(new_n669), .ZN(new_n783));
  INV_X1    g597(.A(new_n672), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n753), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n744), .A2(new_n664), .A3(new_n700), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  AOI21_X1  g602(.A(new_n724), .B1(new_n442), .B2(new_n446), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(new_n583), .A3(new_n654), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n744), .A2(KEYINPUT42), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n654), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n565), .A2(KEYINPUT109), .A3(new_n566), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT109), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n569), .B2(KEYINPUT32), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n582), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n745), .A2(new_n797), .A3(new_n754), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT42), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n227), .ZN(G33));
  NAND4_X1  g615(.A1(new_n789), .A2(new_n583), .A3(new_n654), .A4(new_n716), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  NAND2_X1  g617(.A1(new_n743), .A2(new_n683), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n683), .B2(KEYINPUT111), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n664), .A3(new_n723), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n789), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n621), .A2(new_n630), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(G469), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n632), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT110), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n651), .A3(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n817), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n752), .B(new_n719), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n811), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(KEYINPUT112), .B(G137), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(G39));
  OAI21_X1  g639(.A(new_n752), .B1(new_n820), .B2(new_n821), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n744), .A2(new_n754), .A3(new_n756), .A4(new_n757), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n789), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  NOR2_X1   g645(.A1(G952), .A2(G953), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT119), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n753), .A2(new_n443), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n735), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n779), .A2(new_n806), .A3(new_n271), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(KEYINPUT50), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n750), .A2(new_n751), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n752), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n789), .B(new_n836), .C1(new_n828), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n789), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n270), .A3(new_n753), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n732), .A2(new_n495), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n267), .A3(new_n743), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n845), .A2(new_n806), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n701), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n840), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n797), .A2(new_n754), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT48), .Z(new_n854));
  NAND2_X1  g668(.A1(new_n836), .A2(new_n785), .ZN(new_n855));
  INV_X1    g669(.A(new_n684), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n855), .B(new_n268), .C1(new_n856), .C2(new_n847), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n843), .A2(new_n859), .A3(new_n850), .A4(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n851), .B(new_n858), .C1(new_n861), .C2(KEYINPUT51), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n651), .A2(new_n653), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n696), .A2(new_n699), .A3(new_n712), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n752), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n654), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n770), .A3(new_n732), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n717), .A3(new_n746), .A4(new_n787), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT52), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n646), .A2(new_n656), .A3(new_n716), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n873), .A2(new_n707), .B1(new_n785), .B2(new_n786), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n746), .A4(new_n870), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n442), .A2(new_n443), .A3(new_n446), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n646), .A2(new_n878), .A3(new_n656), .A4(new_n665), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n684), .A2(new_n671), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n657), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n334), .A2(KEYINPUT115), .A3(new_n335), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT115), .B1(new_n334), .B2(new_n335), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n671), .A3(new_n683), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n702), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n657), .B(new_n890), .C1(new_n879), .C2(new_n880), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n882), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n763), .A2(new_n685), .B1(new_n766), .B2(new_n767), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n764), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n852), .A2(new_n654), .A3(new_n745), .A4(new_n789), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n895), .A2(KEYINPUT42), .B1(new_n790), .B2(new_n791), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n714), .A2(new_n883), .A3(new_n884), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n723), .B(new_n897), .C1(new_n756), .C2(new_n757), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n646), .A3(new_n656), .A4(new_n789), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n786), .A2(new_n654), .A3(new_n789), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n900), .A2(new_n802), .A3(new_n901), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n894), .A2(new_n896), .A3(new_n902), .A4(new_n781), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n874), .A2(new_n875), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n877), .A2(new_n904), .A3(KEYINPUT53), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT53), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n888), .B1(KEYINPUT114), .B2(new_n881), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n670), .A2(new_n672), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n910), .A2(new_n759), .A3(new_n690), .A4(new_n336), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n781), .A2(new_n760), .A3(new_n911), .A4(new_n768), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n900), .A2(new_n802), .A3(new_n901), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n800), .A2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n909), .A2(new_n913), .A3(new_n915), .A4(new_n891), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n872), .A2(new_n876), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n906), .A2(new_n907), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n916), .A2(new_n917), .A3(new_n908), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n912), .A2(new_n800), .A3(new_n914), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT116), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n922), .A3(new_n891), .A4(new_n909), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n872), .A2(new_n905), .A3(new_n876), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT116), .B1(new_n892), .B2(new_n903), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n920), .B1(new_n926), .B2(new_n908), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n919), .B1(new_n927), .B2(new_n907), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n833), .B1(new_n862), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n841), .A2(KEYINPUT49), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT113), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n841), .A2(KEYINPUT49), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n804), .A2(new_n645), .A3(new_n724), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n846), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n934), .A3(new_n735), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n929), .A2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n192), .A2(G952), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n272), .B1(new_n906), .B2(new_n918), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(new_n439), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n391), .A2(new_n393), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n423), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  OAI21_X1  g757(.A(new_n938), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(KEYINPUT120), .Z(new_n945));
  NAND2_X1  g759(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(KEYINPUT121), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G51));
  AOI211_X1 g763(.A(new_n272), .B(new_n816), .C1(new_n906), .C2(new_n918), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n632), .B(KEYINPUT57), .Z(new_n951));
  AND3_X1   g765(.A1(new_n906), .A2(new_n907), .A3(new_n918), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n907), .B1(new_n906), .B2(new_n918), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n649), .A2(new_n650), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n950), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT122), .B1(new_n957), .B2(new_n937), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n906), .A2(new_n918), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT54), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n919), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n962), .B2(new_n951), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n959), .B(new_n938), .C1(new_n963), .C2(new_n950), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n958), .A2(new_n964), .ZN(G54));
  NAND3_X1  g779(.A1(new_n939), .A2(KEYINPUT58), .A3(G475), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n261), .A2(new_n235), .ZN(new_n967));
  OR3_X1    g781(.A1(new_n966), .A2(KEYINPUT123), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT123), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n937), .B1(new_n966), .B2(new_n967), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT59), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n675), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n937), .B1(new_n962), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n675), .B1(new_n928), .B2(new_n973), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT124), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g792(.A(KEYINPUT124), .B(new_n675), .C1(new_n928), .C2(new_n973), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  NAND2_X1  g796(.A1(new_n960), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n494), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n984), .B(new_n938), .C1(new_n698), .C2(new_n983), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G66));
  INV_X1    g801(.A(new_n274), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n192), .B1(new_n988), .B2(new_n420), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n909), .A2(new_n913), .A3(new_n891), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(new_n192), .ZN(new_n991));
  INV_X1    g805(.A(G898), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n941), .B1(new_n992), .B2(G953), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n991), .B(new_n993), .ZN(G69));
  AND2_X1   g808(.A1(new_n874), .A2(new_n746), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n738), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n684), .B1(new_n683), .B2(new_n886), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n720), .A2(new_n758), .A3(new_n844), .A4(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n823), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n997), .A2(new_n830), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n192), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n547), .A2(new_n548), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(new_n257), .Z(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT125), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1003), .A2(KEYINPUT125), .A3(new_n1006), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n770), .A2(new_n852), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n822), .B1(new_n811), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n802), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1013), .A2(new_n800), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(new_n192), .A3(new_n830), .A4(new_n995), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1006), .B1(G900), .B2(G953), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1011), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1009), .A2(new_n1010), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1020), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1009), .A2(new_n1022), .A3(new_n1010), .A4(new_n1018), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(G72));
  NAND2_X1  g838(.A1(G472), .A2(G902), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1025), .B(KEYINPUT63), .Z(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n1002), .B2(new_n990), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1027), .B(new_n539), .C1(new_n555), .C2(new_n533), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1015), .A2(new_n830), .A3(new_n995), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1026), .B1(new_n1029), .B2(new_n990), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n549), .A2(new_n534), .A3(new_n561), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT127), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n937), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1028), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(new_n927), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1026), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1036), .B1(new_n578), .B2(new_n554), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(G57));
endmodule


