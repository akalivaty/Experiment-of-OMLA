

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  XOR2_X1 U320 ( .A(n373), .B(n372), .Z(n510) );
  XOR2_X1 U321 ( .A(n373), .B(n362), .Z(n538) );
  XOR2_X1 U322 ( .A(G85GAT), .B(G92GAT), .Z(n410) );
  XNOR2_X1 U323 ( .A(G106GAT), .B(G78GAT), .ZN(n288) );
  XNOR2_X1 U324 ( .A(n288), .B(G148GAT), .ZN(n374) );
  XNOR2_X1 U325 ( .A(n410), .B(n374), .ZN(n289) );
  AND2_X1 U326 ( .A1(G230GAT), .A2(G233GAT), .ZN(n290) );
  NAND2_X1 U327 ( .A1(n289), .A2(n290), .ZN(n294) );
  INV_X1 U328 ( .A(n289), .ZN(n292) );
  INV_X1 U329 ( .A(n290), .ZN(n291) );
  NAND2_X1 U330 ( .A1(n292), .A2(n291), .ZN(n293) );
  NAND2_X1 U331 ( .A1(n294), .A2(n293), .ZN(n295) );
  XNOR2_X1 U332 ( .A(n295), .B(KEYINPUT32), .ZN(n299) );
  XOR2_X1 U333 ( .A(G99GAT), .B(G71GAT), .Z(n296) );
  XOR2_X1 U334 ( .A(G120GAT), .B(n296), .Z(n363) );
  INV_X1 U335 ( .A(n363), .ZN(n297) );
  XNOR2_X1 U336 ( .A(n297), .B(KEYINPUT31), .ZN(n298) );
  XNOR2_X1 U337 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U338 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n301) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n300) );
  XOR2_X1 U340 ( .A(n301), .B(n300), .Z(n302) );
  XNOR2_X1 U341 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U342 ( .A(G57GAT), .B(KEYINPUT13), .Z(n431) );
  XOR2_X1 U343 ( .A(G204GAT), .B(G64GAT), .Z(n359) );
  XNOR2_X1 U344 ( .A(n431), .B(n359), .ZN(n304) );
  XNOR2_X1 U345 ( .A(n305), .B(n304), .ZN(n574) );
  XOR2_X1 U346 ( .A(G29GAT), .B(G36GAT), .Z(n307) );
  XNOR2_X1 U347 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n306) );
  XNOR2_X1 U348 ( .A(n307), .B(n306), .ZN(n409) );
  XOR2_X1 U349 ( .A(G141GAT), .B(G22GAT), .Z(n380) );
  XOR2_X1 U350 ( .A(n409), .B(n380), .Z(n309) );
  NAND2_X1 U351 ( .A1(G229GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U353 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n311) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U356 ( .A(n313), .B(n312), .Z(n321) );
  XOR2_X1 U357 ( .A(G1GAT), .B(G15GAT), .Z(n315) );
  XNOR2_X1 U358 ( .A(KEYINPUT69), .B(G8GAT), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U360 ( .A(KEYINPUT70), .B(n316), .Z(n439) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G43GAT), .Z(n318) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G50GAT), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U364 ( .A(n439), .B(n319), .ZN(n320) );
  XOR2_X1 U365 ( .A(n321), .B(n320), .Z(n570) );
  NOR2_X1 U366 ( .A1(n574), .A2(n570), .ZN(n462) );
  XOR2_X1 U367 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n323) );
  XNOR2_X1 U368 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n322) );
  XNOR2_X1 U369 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U370 ( .A(G127GAT), .B(KEYINPUT78), .Z(n325) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n364) );
  XOR2_X1 U373 ( .A(n364), .B(KEYINPUT5), .Z(n327) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n344) );
  XOR2_X1 U377 ( .A(KEYINPUT1), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U380 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n333) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n332) );
  XNOR2_X1 U382 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(n335), .B(n334), .Z(n342) );
  XOR2_X1 U384 ( .A(G85GAT), .B(G162GAT), .Z(n339) );
  XOR2_X1 U385 ( .A(G155GAT), .B(KEYINPUT2), .Z(n337) );
  XNOR2_X1 U386 ( .A(KEYINPUT84), .B(KEYINPUT3), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n384) );
  XNOR2_X1 U388 ( .A(G29GAT), .B(n384), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U390 ( .A(G134GAT), .B(n340), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U392 ( .A(n344), .B(n343), .ZN(n542) );
  XOR2_X1 U393 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n346) );
  XNOR2_X1 U394 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U396 ( .A(n347), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U397 ( .A(G169GAT), .B(G176GAT), .ZN(n348) );
  XNOR2_X1 U398 ( .A(n349), .B(n348), .ZN(n373) );
  XOR2_X1 U399 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n351) );
  NAND2_X1 U400 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U402 ( .A(KEYINPUT92), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(G36GAT), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U405 ( .A(n355), .B(n354), .Z(n361) );
  XOR2_X1 U406 ( .A(KEYINPUT83), .B(G218GAT), .Z(n357) );
  XNOR2_X1 U407 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U409 ( .A(G197GAT), .B(n358), .ZN(n389) );
  XOR2_X1 U410 ( .A(n389), .B(n359), .Z(n360) );
  XNOR2_X1 U411 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U412 ( .A(n364), .B(n363), .Z(n371) );
  XOR2_X1 U413 ( .A(G43GAT), .B(G134GAT), .Z(n416) );
  XOR2_X1 U414 ( .A(KEYINPUT79), .B(KEYINPUT64), .Z(n366) );
  XNOR2_X1 U415 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U417 ( .A(n416), .B(n367), .Z(n369) );
  NAND2_X1 U418 ( .A1(G227GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U421 ( .A1(n538), .A2(n510), .ZN(n391) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n415) );
  XOR2_X1 U423 ( .A(n415), .B(n374), .Z(n376) );
  NAND2_X1 U424 ( .A1(G228GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U425 ( .A(n376), .B(n375), .ZN(n388) );
  XOR2_X1 U426 ( .A(KEYINPUT81), .B(KEYINPUT22), .Z(n378) );
  XNOR2_X1 U427 ( .A(KEYINPUT24), .B(G204GAT), .ZN(n377) );
  XNOR2_X1 U428 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U429 ( .A(n379), .B(KEYINPUT86), .Z(n382) );
  XNOR2_X1 U430 ( .A(n380), .B(KEYINPUT23), .ZN(n381) );
  XNOR2_X1 U431 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U432 ( .A(n383), .B(KEYINPUT85), .Z(n386) );
  XNOR2_X1 U433 ( .A(n384), .B(KEYINPUT82), .ZN(n385) );
  XNOR2_X1 U434 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U435 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U436 ( .A(n390), .B(n389), .ZN(n543) );
  NAND2_X1 U437 ( .A1(n391), .A2(n543), .ZN(n392) );
  XOR2_X1 U438 ( .A(KEYINPUT25), .B(n392), .Z(n393) );
  XNOR2_X1 U439 ( .A(n393), .B(KEYINPUT96), .ZN(n397) );
  XOR2_X1 U440 ( .A(KEYINPUT27), .B(KEYINPUT94), .Z(n394) );
  XOR2_X1 U441 ( .A(n538), .B(n394), .Z(n401) );
  NOR2_X1 U442 ( .A1(n510), .A2(n543), .ZN(n395) );
  XNOR2_X1 U443 ( .A(KEYINPUT26), .B(n395), .ZN(n568) );
  NAND2_X1 U444 ( .A1(n401), .A2(n568), .ZN(n396) );
  NAND2_X1 U445 ( .A1(n397), .A2(n396), .ZN(n398) );
  XNOR2_X1 U446 ( .A(KEYINPUT97), .B(n398), .ZN(n399) );
  NOR2_X1 U447 ( .A1(n542), .A2(n399), .ZN(n400) );
  XNOR2_X1 U448 ( .A(n400), .B(KEYINPUT98), .ZN(n406) );
  NAND2_X1 U449 ( .A1(n401), .A2(n542), .ZN(n402) );
  XOR2_X1 U450 ( .A(KEYINPUT95), .B(n402), .Z(n507) );
  XOR2_X1 U451 ( .A(n510), .B(KEYINPUT80), .Z(n403) );
  XOR2_X1 U452 ( .A(KEYINPUT28), .B(n543), .Z(n491) );
  INV_X1 U453 ( .A(n491), .ZN(n509) );
  NAND2_X1 U454 ( .A1(n403), .A2(n509), .ZN(n404) );
  NOR2_X1 U455 ( .A1(n507), .A2(n404), .ZN(n405) );
  NOR2_X1 U456 ( .A1(n406), .A2(n405), .ZN(n459) );
  XOR2_X1 U457 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n408) );
  XNOR2_X1 U458 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n407) );
  XOR2_X1 U459 ( .A(n408), .B(n407), .Z(n414) );
  XNOR2_X1 U460 ( .A(n410), .B(n409), .ZN(n412) );
  AND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U462 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U463 ( .A(n414), .B(n413), .ZN(n418) );
  XNOR2_X1 U464 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U465 ( .A(n418), .B(n417), .ZN(n426) );
  XOR2_X1 U466 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n420) );
  XNOR2_X1 U467 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n419) );
  XNOR2_X1 U468 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U469 ( .A(KEYINPUT74), .B(G106GAT), .Z(n422) );
  XNOR2_X1 U470 ( .A(G190GAT), .B(G99GAT), .ZN(n421) );
  XNOR2_X1 U471 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U472 ( .A(n424), .B(n423), .Z(n425) );
  XOR2_X1 U473 ( .A(n426), .B(n425), .Z(n536) );
  INV_X1 U474 ( .A(n536), .ZN(n559) );
  XOR2_X1 U475 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n428) );
  XNOR2_X1 U476 ( .A(G78GAT), .B(G64GAT), .ZN(n427) );
  XNOR2_X1 U477 ( .A(n428), .B(n427), .ZN(n443) );
  XOR2_X1 U478 ( .A(G155GAT), .B(G71GAT), .Z(n430) );
  XNOR2_X1 U479 ( .A(G183GAT), .B(G127GAT), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U481 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U482 ( .A(G22GAT), .B(G211GAT), .ZN(n433) );
  XNOR2_X1 U483 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U484 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n436) );
  NAND2_X1 U485 ( .A1(G231GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U486 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U487 ( .A(n438), .B(n437), .Z(n441) );
  XNOR2_X1 U488 ( .A(n439), .B(KEYINPUT12), .ZN(n440) );
  XNOR2_X1 U489 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U490 ( .A(n443), .B(n442), .ZN(n532) );
  NOR2_X1 U491 ( .A1(n559), .A2(n532), .ZN(n444) );
  XOR2_X1 U492 ( .A(KEYINPUT16), .B(n444), .Z(n445) );
  NOR2_X1 U493 ( .A1(n459), .A2(n445), .ZN(n474) );
  NAND2_X1 U494 ( .A1(n462), .A2(n474), .ZN(n446) );
  XNOR2_X1 U495 ( .A(KEYINPUT99), .B(n446), .ZN(n455) );
  NAND2_X1 U496 ( .A1(n455), .A2(n542), .ZN(n450) );
  XOR2_X1 U497 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n448) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(G1324GAT) );
  NAND2_X1 U501 ( .A1(n455), .A2(n538), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n451), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n453) );
  NAND2_X1 U504 ( .A1(n455), .A2(n510), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(n454), .ZN(G1326GAT) );
  XOR2_X1 U507 ( .A(G22GAT), .B(KEYINPUT103), .Z(n457) );
  NAND2_X1 U508 ( .A1(n455), .A2(n491), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(G1327GAT) );
  XOR2_X1 U510 ( .A(G29GAT), .B(KEYINPUT39), .Z(n466) );
  XOR2_X1 U511 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n464) );
  INV_X1 U512 ( .A(KEYINPUT36), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(n536), .ZN(n580) );
  INV_X1 U514 ( .A(n532), .ZN(n578) );
  NOR2_X1 U515 ( .A1(n578), .A2(n459), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n580), .A2(n460), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT37), .B(n461), .ZN(n485) );
  NAND2_X1 U518 ( .A1(n462), .A2(n485), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n471) );
  NAND2_X1 U520 ( .A1(n471), .A2(n542), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n466), .B(n465), .ZN(G1328GAT) );
  XOR2_X1 U522 ( .A(G36GAT), .B(KEYINPUT105), .Z(n468) );
  NAND2_X1 U523 ( .A1(n471), .A2(n538), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n468), .B(n467), .ZN(G1329GAT) );
  NAND2_X1 U525 ( .A1(n510), .A2(n471), .ZN(n469) );
  XNOR2_X1 U526 ( .A(n469), .B(KEYINPUT40), .ZN(n470) );
  XNOR2_X1 U527 ( .A(G43GAT), .B(n470), .ZN(G1330GAT) );
  NAND2_X1 U528 ( .A1(n471), .A2(n491), .ZN(n472) );
  XNOR2_X1 U529 ( .A(G50GAT), .B(n472), .ZN(G1331GAT) );
  INV_X1 U530 ( .A(n570), .ZN(n549) );
  INV_X1 U531 ( .A(KEYINPUT41), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n574), .B(n473), .ZN(n551) );
  INV_X1 U533 ( .A(n551), .ZN(n526) );
  NOR2_X1 U534 ( .A1(n549), .A2(n526), .ZN(n484) );
  AND2_X1 U535 ( .A1(n474), .A2(n484), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n542), .A2(n480), .ZN(n475) );
  XNOR2_X1 U537 ( .A(KEYINPUT42), .B(n475), .ZN(n476) );
  XNOR2_X1 U538 ( .A(G57GAT), .B(n476), .ZN(G1332GAT) );
  NAND2_X1 U539 ( .A1(n480), .A2(n538), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n477), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U541 ( .A1(n510), .A2(n480), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n478), .B(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U543 ( .A(G71GAT), .B(n479), .ZN(G1334GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n482) );
  NAND2_X1 U545 ( .A1(n480), .A2(n491), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U547 ( .A(G78GAT), .B(n483), .Z(G1335GAT) );
  XNOR2_X1 U548 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n487) );
  AND2_X1 U549 ( .A1(n485), .A2(n484), .ZN(n490) );
  NAND2_X1 U550 ( .A1(n542), .A2(n490), .ZN(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(G1336GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n538), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n488), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U554 ( .A1(n510), .A2(n490), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n489), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U556 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n492), .B(KEYINPUT44), .ZN(n493) );
  XNOR2_X1 U558 ( .A(G106GAT), .B(n493), .ZN(G1339GAT) );
  XOR2_X1 U559 ( .A(G113GAT), .B(KEYINPUT113), .Z(n514) );
  XNOR2_X1 U560 ( .A(KEYINPUT45), .B(KEYINPUT109), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n494), .B(KEYINPUT66), .ZN(n496) );
  AND2_X1 U562 ( .A1(n578), .A2(n580), .ZN(n495) );
  XNOR2_X1 U563 ( .A(n496), .B(n495), .ZN(n497) );
  NOR2_X1 U564 ( .A1(n574), .A2(n497), .ZN(n498) );
  XOR2_X1 U565 ( .A(KEYINPUT110), .B(n498), .Z(n499) );
  NOR2_X1 U566 ( .A1(n549), .A2(n499), .ZN(n505) );
  NAND2_X1 U567 ( .A1(n549), .A2(n551), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n500), .B(KEYINPUT46), .ZN(n501) );
  NAND2_X1 U569 ( .A1(n501), .A2(n532), .ZN(n502) );
  NOR2_X1 U570 ( .A1(n559), .A2(n502), .ZN(n503) );
  XOR2_X1 U571 ( .A(n503), .B(KEYINPUT47), .Z(n504) );
  NOR2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(KEYINPUT48), .B(n506), .ZN(n540) );
  NOR2_X1 U574 ( .A1(n540), .A2(n507), .ZN(n508) );
  XOR2_X1 U575 ( .A(KEYINPUT111), .B(n508), .Z(n523) );
  NAND2_X1 U576 ( .A1(n523), .A2(n509), .ZN(n511) );
  INV_X1 U577 ( .A(n510), .ZN(n548) );
  NOR2_X1 U578 ( .A1(n511), .A2(n548), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(KEYINPUT112), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n549), .A2(n520), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1340GAT) );
  XOR2_X1 U582 ( .A(G120GAT), .B(KEYINPUT49), .Z(n516) );
  NAND2_X1 U583 ( .A1(n551), .A2(n520), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1341GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n518) );
  NAND2_X1 U586 ( .A1(n578), .A2(n520), .ZN(n517) );
  XNOR2_X1 U587 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U588 ( .A(G127GAT), .B(n519), .Z(G1342GAT) );
  XOR2_X1 U589 ( .A(G134GAT), .B(KEYINPUT51), .Z(n522) );
  NAND2_X1 U590 ( .A1(n520), .A2(n559), .ZN(n521) );
  XNOR2_X1 U591 ( .A(n522), .B(n521), .ZN(G1343GAT) );
  NAND2_X1 U592 ( .A1(n523), .A2(n568), .ZN(n535) );
  NOR2_X1 U593 ( .A1(n570), .A2(n535), .ZN(n525) );
  XNOR2_X1 U594 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1344GAT) );
  NOR2_X1 U596 ( .A1(n526), .A2(n535), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n528) );
  XNOR2_X1 U598 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n527) );
  XNOR2_X1 U599 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U600 ( .A(KEYINPUT116), .B(n529), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(G1345GAT) );
  NOR2_X1 U602 ( .A1(n532), .A2(n535), .ZN(n533) );
  XOR2_X1 U603 ( .A(KEYINPUT118), .B(n533), .Z(n534) );
  XNOR2_X1 U604 ( .A(G155GAT), .B(n534), .ZN(G1346GAT) );
  NOR2_X1 U605 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U606 ( .A(G162GAT), .B(n537), .Z(G1347GAT) );
  INV_X1 U607 ( .A(n538), .ZN(n539) );
  NOR2_X1 U608 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(KEYINPUT54), .B(n541), .ZN(n566) );
  INV_X1 U610 ( .A(n542), .ZN(n567) );
  AND2_X1 U611 ( .A1(n567), .A2(n543), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n566), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n545), .B(KEYINPUT119), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n546), .B(KEYINPUT55), .ZN(n547) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n560), .A2(n549), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n553) );
  NAND2_X1 U620 ( .A1(n560), .A2(n551), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1349GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n557) );
  NAND2_X1 U624 ( .A1(n560), .A2(n578), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G183GAT), .B(n558), .ZN(G1350GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n565) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n572) );
  AND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n576) );
  INV_X1 U639 ( .A(n573), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U643 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

