

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777;

  AND2_X1 U377 ( .A1(n427), .A2(KEYINPUT44), .ZN(n469) );
  NOR2_X2 U378 ( .A1(n616), .A2(n615), .ZN(n631) );
  NAND2_X2 U379 ( .A1(n406), .A2(n464), .ZN(n472) );
  NOR2_X2 U380 ( .A1(n669), .A2(n664), .ZN(n670) );
  XNOR2_X2 U381 ( .A(n580), .B(n579), .ZN(n669) );
  XNOR2_X2 U382 ( .A(n508), .B(n489), .ZN(n618) );
  AND2_X1 U383 ( .A1(n436), .A2(n433), .ZN(n438) );
  AND2_X1 U384 ( .A1(n394), .A2(n393), .ZN(n392) );
  AND2_X1 U385 ( .A1(n435), .A2(n433), .ZN(n443) );
  AND2_X1 U386 ( .A1(n434), .A2(n433), .ZN(n437) );
  BUF_X1 U387 ( .A(n363), .Z(n747) );
  NOR2_X1 U388 ( .A1(n469), .A2(n468), .ZN(n471) );
  OR2_X1 U389 ( .A1(n680), .A2(n388), .ZN(n482) );
  XNOR2_X1 U390 ( .A(n385), .B(n369), .ZN(n684) );
  XNOR2_X1 U391 ( .A(n632), .B(n418), .ZN(n775) );
  NOR2_X1 U392 ( .A1(n660), .A2(n659), .ZN(n444) );
  XNOR2_X1 U393 ( .A(n655), .B(KEYINPUT96), .ZN(n656) );
  XNOR2_X1 U394 ( .A(n525), .B(KEYINPUT4), .ZN(n536) );
  XNOR2_X1 U395 ( .A(G143), .B(G128), .ZN(n525) );
  INV_X2 U396 ( .A(G953), .ZN(n765) );
  OR2_X2 U397 ( .A1(n389), .A2(n680), .ZN(n454) );
  XNOR2_X2 U398 ( .A(n510), .B(n475), .ZN(n763) );
  XNOR2_X2 U399 ( .A(n409), .B(G146), .ZN(n510) );
  INV_X1 U400 ( .A(n668), .ZN(n484) );
  NAND2_X2 U401 ( .A1(n460), .A2(n457), .ZN(n614) );
  OR2_X1 U402 ( .A1(n735), .A2(n458), .ZN(n457) );
  AND2_X1 U403 ( .A1(n429), .A2(n461), .ZN(n460) );
  NAND2_X1 U404 ( .A1(n548), .A2(n459), .ZN(n458) );
  NAND2_X1 U405 ( .A1(n465), .A2(n468), .ZN(n464) );
  XNOR2_X1 U406 ( .A(n426), .B(n672), .ZN(n683) );
  NAND2_X1 U407 ( .A1(n384), .A2(n382), .ZN(n426) );
  XNOR2_X1 U408 ( .A(n383), .B(n481), .ZN(n382) );
  NOR2_X1 U409 ( .A1(G953), .A2(G237), .ZN(n538) );
  INV_X1 U410 ( .A(G125), .ZN(n409) );
  NOR2_X1 U411 ( .A1(n356), .A2(n413), .ZN(n412) );
  INV_X1 U412 ( .A(KEYINPUT69), .ZN(n636) );
  XOR2_X1 U413 ( .A(G110), .B(KEYINPUT75), .Z(n498) );
  XNOR2_X1 U414 ( .A(G137), .B(KEYINPUT68), .ZN(n559) );
  XNOR2_X1 U415 ( .A(KEYINPUT10), .B(G140), .ZN(n475) );
  XNOR2_X1 U416 ( .A(n763), .B(n559), .ZN(n408) );
  XNOR2_X1 U417 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U418 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n556) );
  XNOR2_X1 U419 ( .A(G110), .B(KEYINPUT77), .ZN(n554) );
  XNOR2_X1 U420 ( .A(n527), .B(n441), .ZN(n440) );
  INV_X1 U421 ( .A(KEYINPUT7), .ZN(n441) );
  XNOR2_X1 U422 ( .A(n430), .B(n762), .ZN(n735) );
  XNOR2_X1 U423 ( .A(n547), .B(n431), .ZN(n430) );
  XNOR2_X1 U424 ( .A(n432), .B(KEYINPUT78), .ZN(n431) );
  XNOR2_X1 U425 ( .A(n546), .B(n545), .ZN(n547) );
  NAND2_X1 U426 ( .A1(n377), .A2(n374), .ZN(n376) );
  XNOR2_X1 U427 ( .A(n424), .B(KEYINPUT39), .ZN(n648) );
  NOR2_X1 U428 ( .A1(n425), .A2(n610), .ZN(n423) );
  XOR2_X1 U429 ( .A(G478), .B(n531), .Z(n595) );
  INV_X1 U430 ( .A(KEYINPUT6), .ZN(n386) );
  XNOR2_X1 U431 ( .A(n566), .B(KEYINPUT25), .ZN(n421) );
  OR2_X1 U432 ( .A1(n749), .A2(G902), .ZN(n422) );
  NOR2_X1 U433 ( .A1(n359), .A2(KEYINPUT84), .ZN(n402) );
  AND2_X1 U434 ( .A1(n451), .A2(n447), .ZN(n446) );
  INV_X1 U435 ( .A(KEYINPUT104), .ZN(n481) );
  INV_X1 U436 ( .A(KEYINPUT47), .ZN(n420) );
  NAND2_X1 U437 ( .A1(G234), .A2(G237), .ZN(n491) );
  OR2_X1 U438 ( .A1(G237), .A2(G902), .ZN(n507) );
  INV_X1 U439 ( .A(G902), .ZN(n459) );
  NAND2_X1 U440 ( .A1(n735), .A2(G469), .ZN(n429) );
  NAND2_X1 U441 ( .A1(G469), .A2(G902), .ZN(n461) );
  NOR2_X1 U442 ( .A1(n677), .A2(n659), .ZN(n599) );
  XNOR2_X1 U443 ( .A(G902), .B(KEYINPUT15), .ZN(n506) );
  XNOR2_X1 U444 ( .A(n536), .B(n535), .ZN(n542) );
  XNOR2_X1 U445 ( .A(G131), .B(G134), .ZN(n535) );
  XNOR2_X1 U446 ( .A(G146), .B(G113), .ZN(n540) );
  XNOR2_X1 U447 ( .A(n539), .B(n362), .ZN(n381) );
  AND2_X1 U448 ( .A1(n470), .A2(n466), .ZN(n406) );
  AND2_X1 U449 ( .A1(n467), .A2(n686), .ZN(n466) );
  XOR2_X1 U450 ( .A(KEYINPUT102), .B(G122), .Z(n512) );
  XNOR2_X1 U451 ( .A(G143), .B(G131), .ZN(n511) );
  AND2_X1 U452 ( .A1(G227), .A2(n765), .ZN(n487) );
  XNOR2_X1 U453 ( .A(G146), .B(G104), .ZN(n543) );
  XOR2_X1 U454 ( .A(G110), .B(G107), .Z(n490) );
  INV_X1 U455 ( .A(G140), .ZN(n432) );
  XNOR2_X1 U456 ( .A(n542), .B(n559), .ZN(n762) );
  XNOR2_X1 U457 ( .A(n501), .B(KEYINPUT18), .ZN(n502) );
  XOR2_X1 U458 ( .A(KEYINPUT17), .B(KEYINPUT79), .Z(n500) );
  XNOR2_X1 U459 ( .A(n636), .B(KEYINPUT48), .ZN(n637) );
  NOR2_X1 U460 ( .A1(n411), .A2(n410), .ZN(n638) );
  XNOR2_X1 U461 ( .A(n509), .B(n646), .ZN(n634) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n617) );
  XOR2_X1 U463 ( .A(KEYINPUT70), .B(n612), .Z(n622) );
  AND2_X1 U464 ( .A1(n677), .A2(n611), .ZN(n612) );
  INV_X1 U465 ( .A(n681), .ZN(n453) );
  NAND2_X1 U466 ( .A1(n599), .A2(n614), .ZN(n667) );
  XNOR2_X1 U467 ( .A(n532), .B(KEYINPUT103), .ZN(n660) );
  XNOR2_X1 U468 ( .A(n378), .B(n537), .ZN(n698) );
  XNOR2_X1 U469 ( .A(n542), .B(n379), .ZN(n378) );
  XNOR2_X1 U470 ( .A(n381), .B(n380), .ZN(n379) );
  XNOR2_X1 U471 ( .A(n540), .B(KEYINPUT5), .ZN(n380) );
  XNOR2_X1 U472 ( .A(KEYINPUT16), .B(KEYINPUT74), .ZN(n497) );
  INV_X1 U473 ( .A(n359), .ZN(n405) );
  NAND2_X1 U474 ( .A1(n456), .A2(n455), .ZN(n385) );
  INV_X1 U475 ( .A(n671), .ZN(n455) );
  NOR2_X1 U476 ( .A1(n450), .A2(n449), .ZN(n448) );
  XNOR2_X1 U477 ( .A(n614), .B(n549), .ZN(n678) );
  NAND2_X1 U478 ( .A1(n666), .A2(n452), .ZN(n451) );
  NOR2_X1 U479 ( .A1(n667), .A2(n453), .ZN(n452) );
  BUF_X1 U480 ( .A(n662), .Z(n442) );
  XNOR2_X1 U481 ( .A(n358), .B(KEYINPUT71), .ZN(n757) );
  XNOR2_X1 U482 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U483 ( .A(n558), .B(n408), .ZN(n564) );
  XNOR2_X1 U484 ( .A(G128), .B(G119), .ZN(n561) );
  XNOR2_X1 U485 ( .A(n440), .B(n526), .ZN(n528) );
  INV_X1 U486 ( .A(KEYINPUT42), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n635), .B(n419), .ZN(n773) );
  INV_X1 U488 ( .A(KEYINPUT40), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n676), .B(KEYINPUT32), .ZN(n480) );
  XNOR2_X1 U490 ( .A(n738), .B(n739), .ZN(n439) );
  AND2_X1 U491 ( .A1(n398), .A2(n397), .ZN(n396) );
  AND2_X1 U492 ( .A1(n773), .A2(KEYINPUT46), .ZN(n356) );
  XOR2_X1 U493 ( .A(n498), .B(n497), .Z(n357) );
  XOR2_X1 U494 ( .A(G119), .B(KEYINPUT3), .Z(n358) );
  NAND2_X1 U495 ( .A1(n387), .A2(n476), .ZN(n359) );
  XNOR2_X1 U496 ( .A(KEYINPUT80), .B(n649), .ZN(n360) );
  XOR2_X1 U497 ( .A(n510), .B(n500), .Z(n361) );
  AND2_X1 U498 ( .A1(G210), .A2(n538), .ZN(n362) );
  AND2_X2 U499 ( .A1(n376), .A2(n359), .ZN(n363) );
  NAND2_X1 U500 ( .A1(n692), .A2(n765), .ZN(n364) );
  INV_X1 U501 ( .A(n577), .ZN(n661) );
  XNOR2_X1 U502 ( .A(n681), .B(n386), .ZN(n577) );
  AND2_X1 U503 ( .A1(n476), .A2(n697), .ZN(n365) );
  XOR2_X1 U504 ( .A(n620), .B(n420), .Z(n366) );
  AND2_X1 U505 ( .A1(n439), .A2(n433), .ZN(G54) );
  XOR2_X1 U506 ( .A(KEYINPUT31), .B(KEYINPUT100), .Z(n368) );
  XNOR2_X1 U507 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n369) );
  XOR2_X1 U508 ( .A(KEYINPUT73), .B(KEYINPUT34), .Z(n370) );
  XNOR2_X1 U509 ( .A(KEYINPUT110), .B(n699), .ZN(n371) );
  XNOR2_X1 U510 ( .A(n733), .B(n732), .ZN(n372) );
  XOR2_X1 U511 ( .A(n741), .B(n740), .Z(n373) );
  OR2_X1 U512 ( .A1(n695), .A2(n694), .ZN(n374) );
  AND2_X1 U513 ( .A1(n693), .A2(n486), .ZN(n375) );
  INV_X1 U514 ( .A(n751), .ZN(n433) );
  XNOR2_X2 U515 ( .A(n472), .B(n687), .ZN(n476) );
  NAND2_X1 U516 ( .A1(n365), .A2(n764), .ZN(n377) );
  XNOR2_X1 U517 ( .A(n757), .B(n544), .ZN(n537) );
  NAND2_X1 U518 ( .A1(n483), .A2(n482), .ZN(n383) );
  NAND2_X1 U519 ( .A1(n684), .A2(KEYINPUT44), .ZN(n384) );
  XNOR2_X2 U520 ( .A(n541), .B(G472), .ZN(n681) );
  NOR2_X1 U521 ( .A1(n689), .A2(n360), .ZN(n387) );
  NAND2_X1 U522 ( .A1(n663), .A2(n577), .ZN(n388) );
  NAND2_X1 U523 ( .A1(n675), .A2(n577), .ZN(n389) );
  NAND2_X1 U524 ( .A1(n390), .A2(n617), .ZN(n477) );
  NOR2_X1 U525 ( .A1(n639), .A2(n390), .ZN(n626) );
  NAND2_X1 U526 ( .A1(n618), .A2(n640), .ZN(n390) );
  NAND2_X1 U527 ( .A1(n396), .A2(n391), .ZN(G75) );
  NAND2_X1 U528 ( .A1(n395), .A2(n392), .ZN(n391) );
  INV_X1 U529 ( .A(n693), .ZN(n393) );
  NAND2_X1 U530 ( .A1(n399), .A2(n486), .ZN(n394) );
  INV_X1 U531 ( .A(n400), .ZN(n395) );
  NAND2_X1 U532 ( .A1(n399), .A2(n375), .ZN(n397) );
  NAND2_X1 U533 ( .A1(n400), .A2(n693), .ZN(n398) );
  INV_X1 U534 ( .A(n473), .ZN(n399) );
  NAND2_X1 U535 ( .A1(n403), .A2(n401), .ZN(n400) );
  NOR2_X1 U536 ( .A1(n364), .A2(n402), .ZN(n401) );
  NAND2_X1 U537 ( .A1(n473), .A2(n404), .ZN(n403) );
  NOR2_X1 U538 ( .A1(n486), .A2(n405), .ZN(n404) );
  NAND2_X1 U539 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U540 ( .A(n407), .B(KEYINPUT22), .ZN(n680) );
  NAND2_X1 U541 ( .A1(n477), .A2(n479), .ZN(n657) );
  NAND2_X1 U542 ( .A1(n777), .A2(n711), .ZN(n427) );
  XNOR2_X2 U543 ( .A(n454), .B(n480), .ZN(n777) );
  NAND2_X1 U544 ( .A1(n445), .A2(n444), .ZN(n407) );
  INV_X1 U545 ( .A(KEYINPUT87), .ZN(n468) );
  NAND2_X1 U546 ( .A1(n469), .A2(n468), .ZN(n467) );
  NAND2_X1 U547 ( .A1(n366), .A2(n415), .ZN(n410) );
  NAND2_X1 U548 ( .A1(n412), .A2(n628), .ZN(n411) );
  NAND2_X1 U549 ( .A1(n414), .A2(n621), .ZN(n413) );
  NAND2_X1 U550 ( .A1(n775), .A2(KEYINPUT46), .ZN(n414) );
  NAND2_X1 U551 ( .A1(n417), .A2(n416), .ZN(n415) );
  INV_X1 U552 ( .A(n773), .ZN(n416) );
  NOR2_X1 U553 ( .A1(n775), .A2(KEYINPUT46), .ZN(n417) );
  XNOR2_X2 U554 ( .A(n422), .B(n421), .ZN(n677) );
  NAND2_X1 U555 ( .A1(n606), .A2(n609), .ZN(n633) );
  NAND2_X1 U556 ( .A1(n606), .A2(n423), .ZN(n424) );
  INV_X1 U557 ( .A(n634), .ZN(n425) );
  NOR2_X1 U558 ( .A1(n427), .A2(KEYINPUT44), .ZN(n685) );
  NAND2_X1 U559 ( .A1(n666), .A2(n428), .ZN(n447) );
  AND2_X1 U560 ( .A1(n665), .A2(n368), .ZN(n428) );
  INV_X1 U561 ( .A(n664), .ZN(n666) );
  XNOR2_X1 U562 ( .A(n700), .B(n371), .ZN(n436) );
  XNOR2_X1 U563 ( .A(n734), .B(n372), .ZN(n435) );
  XNOR2_X1 U564 ( .A(n742), .B(n373), .ZN(n434) );
  INV_X1 U565 ( .A(n678), .ZN(n662) );
  NAND2_X1 U566 ( .A1(n630), .A2(n631), .ZN(n632) );
  XNOR2_X1 U567 ( .A(n437), .B(n743), .ZN(G60) );
  XNOR2_X1 U568 ( .A(n438), .B(n701), .ZN(G57) );
  XNOR2_X1 U569 ( .A(n443), .B(KEYINPUT56), .ZN(G51) );
  INV_X1 U570 ( .A(n664), .ZN(n445) );
  XNOR2_X2 U571 ( .A(n658), .B(KEYINPUT0), .ZN(n664) );
  NAND2_X1 U572 ( .A1(n448), .A2(n447), .ZN(n724) );
  NAND2_X1 U573 ( .A1(n446), .A2(n448), .ZN(n485) );
  NOR2_X1 U574 ( .A1(n666), .A2(n368), .ZN(n449) );
  NOR2_X1 U575 ( .A1(n665), .A2(n368), .ZN(n450) );
  INV_X1 U576 ( .A(n451), .ZN(n705) );
  XNOR2_X1 U577 ( .A(n670), .B(n370), .ZN(n456) );
  XNOR2_X1 U578 ( .A(n462), .B(n361), .ZN(n505) );
  XNOR2_X1 U579 ( .A(n462), .B(G101), .ZN(n756) );
  XNOR2_X2 U580 ( .A(n499), .B(n357), .ZN(n462) );
  INV_X1 U581 ( .A(n523), .ZN(n494) );
  XNOR2_X2 U582 ( .A(n463), .B(G107), .ZN(n523) );
  XNOR2_X2 U583 ( .A(G122), .B(G116), .ZN(n463) );
  INV_X1 U584 ( .A(n683), .ZN(n465) );
  NAND2_X1 U585 ( .A1(n683), .A2(n471), .ZN(n470) );
  INV_X1 U586 ( .A(n482), .ZN(n702) );
  XNOR2_X2 U587 ( .A(n474), .B(KEYINPUT81), .ZN(n473) );
  NAND2_X1 U588 ( .A1(n691), .A2(n488), .ZN(n474) );
  NOR2_X1 U589 ( .A1(n476), .A2(KEYINPUT2), .ZN(n688) );
  NAND2_X1 U590 ( .A1(n476), .A2(n765), .ZN(n755) );
  NAND2_X1 U591 ( .A1(n618), .A2(n478), .ZN(n479) );
  AND2_X1 U592 ( .A1(n640), .A2(n619), .ZN(n478) );
  NAND2_X1 U593 ( .A1(n485), .A2(n484), .ZN(n483) );
  INV_X1 U594 ( .A(KEYINPUT84), .ZN(n486) );
  NOR2_X1 U595 ( .A1(n681), .A2(n578), .ZN(n665) );
  NOR2_X1 U596 ( .A1(n442), .A2(n677), .ZN(n663) );
  OR2_X1 U597 ( .A1(KEYINPUT2), .A2(n764), .ZN(n488) );
  AND2_X1 U598 ( .A1(n507), .A2(G210), .ZN(n489) );
  XNOR2_X1 U599 ( .A(n544), .B(n487), .ZN(n545) );
  INV_X1 U600 ( .A(n525), .ZN(n526) );
  NAND2_X1 U601 ( .A1(n363), .A2(G472), .ZN(n700) );
  NOR2_X1 U602 ( .A1(G952), .A2(n765), .ZN(n751) );
  XOR2_X1 U603 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n492) );
  XNOR2_X1 U604 ( .A(n492), .B(n491), .ZN(n603) );
  NAND2_X1 U605 ( .A1(n603), .A2(G952), .ZN(n601) );
  NAND2_X1 U606 ( .A1(G214), .A2(n507), .ZN(n640) );
  XNOR2_X1 U607 ( .A(KEYINPUT76), .B(KEYINPUT38), .ZN(n509) );
  XOR2_X1 U608 ( .A(G113), .B(G104), .Z(n514) );
  NAND2_X1 U609 ( .A1(n523), .A2(n514), .ZN(n496) );
  INV_X1 U610 ( .A(n514), .ZN(n493) );
  NAND2_X1 U611 ( .A1(n494), .A2(n493), .ZN(n495) );
  NAND2_X1 U612 ( .A1(n496), .A2(n495), .ZN(n499) );
  XOR2_X1 U613 ( .A(KEYINPUT67), .B(G101), .Z(n544) );
  AND2_X1 U614 ( .A1(G224), .A2(n765), .ZN(n501) );
  XNOR2_X1 U615 ( .A(n536), .B(n502), .ZN(n503) );
  XNOR2_X1 U616 ( .A(n537), .B(n503), .ZN(n504) );
  XNOR2_X1 U617 ( .A(n505), .B(n504), .ZN(n731) );
  XNOR2_X1 U618 ( .A(n506), .B(KEYINPUT92), .ZN(n696) );
  NAND2_X1 U619 ( .A1(n731), .A2(n696), .ZN(n508) );
  INV_X1 U620 ( .A(n618), .ZN(n646) );
  NAND2_X1 U621 ( .A1(n640), .A2(n634), .ZN(n583) );
  XNOR2_X1 U622 ( .A(KEYINPUT13), .B(G475), .ZN(n522) );
  XNOR2_X1 U623 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U624 ( .A(n763), .B(n513), .ZN(n520) );
  XNOR2_X1 U625 ( .A(n514), .B(KEYINPUT12), .ZN(n518) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n516) );
  NAND2_X1 U627 ( .A1(n538), .A2(G214), .ZN(n515) );
  XNOR2_X1 U628 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U629 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U630 ( .A(n520), .B(n519), .ZN(n741) );
  NOR2_X1 U631 ( .A1(G902), .A2(n741), .ZN(n521) );
  XNOR2_X1 U632 ( .A(n522), .B(n521), .ZN(n596) );
  NAND2_X1 U633 ( .A1(G234), .A2(n765), .ZN(n524) );
  XOR2_X1 U634 ( .A(KEYINPUT8), .B(n524), .Z(n560) );
  NAND2_X1 U635 ( .A1(n560), .A2(G217), .ZN(n529) );
  XNOR2_X1 U636 ( .A(G134), .B(KEYINPUT9), .ZN(n527) );
  XNOR2_X1 U637 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U638 ( .A(n523), .B(n530), .ZN(n745) );
  NOR2_X1 U639 ( .A1(G902), .A2(n745), .ZN(n531) );
  NOR2_X1 U640 ( .A1(n596), .A2(n595), .ZN(n532) );
  NOR2_X1 U641 ( .A1(n583), .A2(n660), .ZN(n534) );
  XOR2_X1 U642 ( .A(KEYINPUT109), .B(KEYINPUT41), .Z(n533) );
  XNOR2_X1 U643 ( .A(n534), .B(n533), .ZN(n629) );
  XOR2_X1 U644 ( .A(G116), .B(G137), .Z(n539) );
  NOR2_X1 U645 ( .A1(n698), .A2(G902), .ZN(n541) );
  XNOR2_X1 U646 ( .A(n490), .B(n543), .ZN(n546) );
  INV_X1 U647 ( .A(G469), .ZN(n548) );
  INV_X1 U648 ( .A(KEYINPUT1), .ZN(n549) );
  NAND2_X1 U649 ( .A1(n696), .A2(G234), .ZN(n551) );
  XNOR2_X1 U650 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n550) );
  XNOR2_X1 U651 ( .A(n551), .B(n550), .ZN(n565) );
  NAND2_X1 U652 ( .A1(G221), .A2(n565), .ZN(n553) );
  XOR2_X1 U653 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n552) );
  XNOR2_X1 U654 ( .A(n553), .B(n552), .ZN(n659) );
  XOR2_X1 U655 ( .A(KEYINPUT23), .B(KEYINPUT97), .Z(n555) );
  XNOR2_X1 U656 ( .A(n555), .B(n554), .ZN(n557) );
  AND2_X1 U657 ( .A1(n560), .A2(G221), .ZN(n562) );
  XNOR2_X1 U658 ( .A(n564), .B(n563), .ZN(n749) );
  NAND2_X1 U659 ( .A1(G217), .A2(n565), .ZN(n566) );
  NAND2_X1 U660 ( .A1(n662), .A2(n599), .ZN(n578) );
  XOR2_X1 U661 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n568) );
  NOR2_X1 U662 ( .A1(n442), .A2(n599), .ZN(n567) );
  XOR2_X1 U663 ( .A(n568), .B(n567), .Z(n569) );
  NAND2_X1 U664 ( .A1(n681), .A2(n569), .ZN(n572) );
  AND2_X1 U665 ( .A1(n659), .A2(n677), .ZN(n570) );
  XOR2_X1 U666 ( .A(KEYINPUT49), .B(n570), .Z(n571) );
  NOR2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U668 ( .A(n573), .B(KEYINPUT118), .ZN(n574) );
  NOR2_X1 U669 ( .A1(n665), .A2(n574), .ZN(n575) );
  XOR2_X1 U670 ( .A(KEYINPUT51), .B(n575), .Z(n576) );
  NOR2_X1 U671 ( .A1(n629), .A2(n576), .ZN(n589) );
  NOR2_X1 U672 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U673 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n579) );
  NOR2_X1 U674 ( .A1(n640), .A2(n634), .ZN(n581) );
  NOR2_X1 U675 ( .A1(n660), .A2(n581), .ZN(n586) );
  INV_X1 U676 ( .A(n596), .ZN(n582) );
  NOR2_X1 U677 ( .A1(n595), .A2(n582), .ZN(n720) );
  NAND2_X1 U678 ( .A1(n582), .A2(n595), .ZN(n712) );
  INV_X1 U679 ( .A(n712), .ZN(n723) );
  NOR2_X1 U680 ( .A1(n720), .A2(n723), .ZN(n668) );
  NOR2_X1 U681 ( .A1(n668), .A2(n583), .ZN(n584) );
  XOR2_X1 U682 ( .A(KEYINPUT119), .B(n584), .Z(n585) );
  NOR2_X1 U683 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U684 ( .A1(n669), .A2(n587), .ZN(n588) );
  NOR2_X1 U685 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U686 ( .A(n590), .B(KEYINPUT52), .ZN(n591) );
  NOR2_X1 U687 ( .A1(n601), .A2(n591), .ZN(n593) );
  NOR2_X1 U688 ( .A1(n669), .A2(n629), .ZN(n592) );
  NOR2_X1 U689 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U690 ( .A(KEYINPUT120), .B(n594), .ZN(n692) );
  NAND2_X1 U691 ( .A1(n596), .A2(n595), .ZN(n671) );
  XOR2_X1 U692 ( .A(KEYINPUT107), .B(KEYINPUT30), .Z(n598) );
  NAND2_X1 U693 ( .A1(n453), .A2(n640), .ZN(n597) );
  XNOR2_X1 U694 ( .A(n598), .B(n597), .ZN(n600) );
  NOR2_X1 U695 ( .A1(n600), .A2(n667), .ZN(n606) );
  NOR2_X1 U696 ( .A1(G953), .A2(n601), .ZN(n602) );
  XOR2_X1 U697 ( .A(KEYINPUT94), .B(n602), .Z(n654) );
  NAND2_X1 U698 ( .A1(n603), .A2(G902), .ZN(n650) );
  NOR2_X1 U699 ( .A1(G900), .A2(n650), .ZN(n604) );
  NAND2_X1 U700 ( .A1(G953), .A2(n604), .ZN(n605) );
  NAND2_X1 U701 ( .A1(n654), .A2(n605), .ZN(n609) );
  NOR2_X1 U702 ( .A1(n646), .A2(n633), .ZN(n607) );
  XOR2_X1 U703 ( .A(KEYINPUT108), .B(n607), .Z(n608) );
  NOR2_X1 U704 ( .A1(n671), .A2(n608), .ZN(n715) );
  INV_X1 U705 ( .A(n715), .ZN(n621) );
  INV_X1 U706 ( .A(n609), .ZN(n610) );
  NOR2_X1 U707 ( .A1(n659), .A2(n610), .ZN(n611) );
  NOR2_X1 U708 ( .A1(n622), .A2(n681), .ZN(n613) );
  XOR2_X1 U709 ( .A(KEYINPUT28), .B(n613), .Z(n616) );
  INV_X1 U710 ( .A(n614), .ZN(n615) );
  INV_X1 U711 ( .A(n617), .ZN(n619) );
  NAND2_X1 U712 ( .A1(n631), .A2(n657), .ZN(n716) );
  NOR2_X1 U713 ( .A1(n668), .A2(n716), .ZN(n620) );
  XNOR2_X1 U714 ( .A(KEYINPUT91), .B(n442), .ZN(n673) );
  INV_X1 U715 ( .A(n720), .ZN(n717) );
  NOR2_X1 U716 ( .A1(n622), .A2(n717), .ZN(n623) );
  NAND2_X1 U717 ( .A1(n623), .A2(n661), .ZN(n624) );
  XOR2_X1 U718 ( .A(KEYINPUT105), .B(n624), .Z(n639) );
  XNOR2_X1 U719 ( .A(KEYINPUT89), .B(KEYINPUT36), .ZN(n625) );
  XNOR2_X1 U720 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X1 U721 ( .A1(n673), .A2(n627), .ZN(n727) );
  INV_X1 U722 ( .A(n727), .ZN(n628) );
  INV_X1 U723 ( .A(n629), .ZN(n630) );
  NAND2_X1 U724 ( .A1(n648), .A2(n720), .ZN(n635) );
  XNOR2_X1 U725 ( .A(n638), .B(n637), .ZN(n647) );
  XNOR2_X1 U726 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n644) );
  INV_X1 U727 ( .A(n639), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U729 ( .A1(n442), .A2(n642), .ZN(n643) );
  XOR2_X1 U730 ( .A(n644), .B(n643), .Z(n645) );
  NAND2_X1 U731 ( .A1(n646), .A2(n645), .ZN(n730) );
  NAND2_X1 U732 ( .A1(n647), .A2(n730), .ZN(n689) );
  NAND2_X1 U733 ( .A1(n723), .A2(n648), .ZN(n729) );
  NAND2_X1 U734 ( .A1(KEYINPUT2), .A2(n729), .ZN(n649) );
  INV_X1 U735 ( .A(n650), .ZN(n651) );
  NOR2_X1 U736 ( .A1(G898), .A2(n765), .ZN(n759) );
  NAND2_X1 U737 ( .A1(n651), .A2(n759), .ZN(n652) );
  XOR2_X1 U738 ( .A(KEYINPUT95), .B(n652), .Z(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n655) );
  INV_X1 U740 ( .A(n677), .ZN(n674) );
  INV_X1 U741 ( .A(KEYINPUT88), .ZN(n672) );
  INV_X1 U742 ( .A(KEYINPUT65), .ZN(n676) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U746 ( .A1(n682), .A2(n681), .ZN(n711) );
  INV_X1 U747 ( .A(n684), .ZN(n776) );
  NAND2_X1 U748 ( .A1(n685), .A2(n776), .ZN(n686) );
  XNOR2_X1 U749 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(KEYINPUT83), .ZN(n691) );
  INV_X1 U751 ( .A(n729), .ZN(n690) );
  NOR2_X2 U752 ( .A1(n690), .A2(n689), .ZN(n764) );
  XNOR2_X1 U753 ( .A(KEYINPUT121), .B(KEYINPUT53), .ZN(n693) );
  INV_X1 U754 ( .A(KEYINPUT2), .ZN(n695) );
  XOR2_X1 U755 ( .A(n696), .B(KEYINPUT85), .Z(n694) );
  INV_X1 U756 ( .A(n696), .ZN(n697) );
  XOR2_X1 U757 ( .A(n698), .B(KEYINPUT62), .Z(n699) );
  XOR2_X1 U758 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n701) );
  XOR2_X1 U759 ( .A(n702), .B(G101), .Z(G3) );
  XOR2_X1 U760 ( .A(G104), .B(KEYINPUT111), .Z(n704) );
  NAND2_X1 U761 ( .A1(n705), .A2(n720), .ZN(n703) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(G6) );
  XNOR2_X1 U763 ( .A(G107), .B(KEYINPUT27), .ZN(n709) );
  XOR2_X1 U764 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n707) );
  NAND2_X1 U765 ( .A1(n705), .A2(n723), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U767 ( .A(n709), .B(n708), .ZN(G9) );
  XOR2_X1 U768 ( .A(G110), .B(KEYINPUT113), .Z(n710) );
  XNOR2_X1 U769 ( .A(n711), .B(n710), .ZN(G12) );
  NOR2_X1 U770 ( .A1(n712), .A2(n716), .ZN(n714) );
  XNOR2_X1 U771 ( .A(G128), .B(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n714), .B(n713), .ZN(G30) );
  XOR2_X1 U773 ( .A(G143), .B(n715), .Z(G45) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT114), .B(n718), .Z(n719) );
  XNOR2_X1 U776 ( .A(G146), .B(n719), .ZN(G48) );
  XOR2_X1 U777 ( .A(G113), .B(KEYINPUT115), .Z(n722) );
  NAND2_X1 U778 ( .A1(n720), .A2(n724), .ZN(n721) );
  XNOR2_X1 U779 ( .A(n722), .B(n721), .ZN(G15) );
  NAND2_X1 U780 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT116), .ZN(n726) );
  XNOR2_X1 U782 ( .A(G116), .B(n726), .ZN(G18) );
  XNOR2_X1 U783 ( .A(G125), .B(n727), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U785 ( .A(G134), .B(n729), .ZN(G36) );
  XNOR2_X1 U786 ( .A(G140), .B(n730), .ZN(G42) );
  NAND2_X1 U787 ( .A1(n363), .A2(G210), .ZN(n734) );
  XOR2_X1 U788 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n733) );
  XNOR2_X1 U789 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  XOR2_X1 U790 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n737) );
  XNOR2_X1 U791 ( .A(n735), .B(KEYINPUT123), .ZN(n736) );
  XNOR2_X1 U792 ( .A(n737), .B(n736), .ZN(n739) );
  NAND2_X1 U793 ( .A1(n747), .A2(G469), .ZN(n738) );
  NAND2_X1 U794 ( .A1(n363), .A2(G475), .ZN(n742) );
  XOR2_X1 U795 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n740) );
  XOR2_X1 U796 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n743) );
  NAND2_X1 U797 ( .A1(G478), .A2(n747), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U799 ( .A1(n751), .A2(n746), .ZN(G63) );
  NAND2_X1 U800 ( .A1(G217), .A2(n747), .ZN(n748) );
  XNOR2_X1 U801 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(G66) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n752) );
  XNOR2_X1 U804 ( .A(KEYINPUT61), .B(n752), .ZN(n753) );
  NAND2_X1 U805 ( .A1(n753), .A2(G898), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n757), .B(n756), .ZN(n758) );
  NOR2_X1 U808 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(G69) );
  XNOR2_X1 U810 ( .A(n762), .B(n763), .ZN(n767) );
  XOR2_X1 U811 ( .A(n764), .B(n767), .Z(n766) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(n772) );
  XNOR2_X1 U813 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U814 ( .A1(n768), .A2(G900), .ZN(n769) );
  XNOR2_X1 U815 ( .A(KEYINPUT126), .B(n769), .ZN(n770) );
  NAND2_X1 U816 ( .A1(G953), .A2(n770), .ZN(n771) );
  NAND2_X1 U817 ( .A1(n772), .A2(n771), .ZN(G72) );
  XNOR2_X1 U818 ( .A(G131), .B(KEYINPUT127), .ZN(n774) );
  XNOR2_X1 U819 ( .A(n774), .B(n773), .ZN(G33) );
  XOR2_X1 U820 ( .A(G137), .B(n775), .Z(G39) );
  XNOR2_X1 U821 ( .A(G122), .B(n776), .ZN(G24) );
  XNOR2_X1 U822 ( .A(n777), .B(G119), .ZN(G21) );
endmodule

