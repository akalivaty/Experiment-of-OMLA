

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606;

  XNOR2_X2 U329 ( .A(n424), .B(n423), .ZN(n563) );
  NOR2_X2 U330 ( .A1(n421), .A2(n420), .ZN(n424) );
  XNOR2_X1 U331 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n430), .B(n299), .ZN(n317) );
  XOR2_X1 U333 ( .A(G176GAT), .B(KEYINPUT19), .Z(n426) );
  XNOR2_X1 U334 ( .A(n422), .B(KEYINPUT48), .ZN(n423) );
  XNOR2_X1 U335 ( .A(n335), .B(n334), .ZN(n496) );
  XNOR2_X1 U336 ( .A(n333), .B(n332), .ZN(n334) );
  NOR2_X1 U337 ( .A1(n544), .A2(n565), .ZN(n549) );
  XNOR2_X1 U338 ( .A(n461), .B(KEYINPUT55), .ZN(n476) );
  XNOR2_X1 U339 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U340 ( .A(KEYINPUT105), .B(n513), .Z(n297) );
  XOR2_X1 U341 ( .A(n427), .B(KEYINPUT18), .Z(n298) );
  AND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XOR2_X1 U343 ( .A(KEYINPUT10), .B(KEYINPUT80), .Z(n300) );
  INV_X1 U344 ( .A(KEYINPUT47), .ZN(n411) );
  XNOR2_X1 U345 ( .A(n411), .B(KEYINPUT114), .ZN(n412) );
  XNOR2_X1 U346 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U347 ( .A(n394), .B(n393), .ZN(n399) );
  INV_X1 U348 ( .A(n538), .ZN(n459) );
  XNOR2_X1 U349 ( .A(n401), .B(KEYINPUT66), .ZN(n402) );
  AND2_X1 U350 ( .A1(n460), .A2(n459), .ZN(n590) );
  AND2_X1 U351 ( .A1(n476), .A2(n550), .ZN(n585) );
  XNOR2_X1 U352 ( .A(KEYINPUT95), .B(n492), .ZN(n538) );
  XOR2_X1 U353 ( .A(G204GAT), .B(KEYINPUT21), .Z(n302) );
  XNOR2_X1 U354 ( .A(G197GAT), .B(G218GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n429) );
  XOR2_X1 U356 ( .A(n429), .B(KEYINPUT22), .Z(n304) );
  NAND2_X1 U357 ( .A1(G228GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U359 ( .A(n305), .B(KEYINPUT93), .Z(n307) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G141GAT), .Z(n392) );
  XNOR2_X1 U361 ( .A(n392), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U363 ( .A(KEYINPUT24), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U364 ( .A(KEYINPUT23), .B(G211GAT), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U366 ( .A(n311), .B(n310), .Z(n315) );
  XNOR2_X1 U367 ( .A(G22GAT), .B(G155GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n312), .B(G78GAT), .ZN(n352) );
  XNOR2_X1 U369 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n313), .B(KEYINPUT3), .ZN(n442) );
  XNOR2_X1 U371 ( .A(n352), .B(n442), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n486) );
  XNOR2_X1 U373 ( .A(G162GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n300), .B(n316), .ZN(n318) );
  XOR2_X1 U375 ( .A(KEYINPUT83), .B(G92GAT), .Z(n430) );
  XOR2_X1 U376 ( .A(n319), .B(G29GAT), .Z(n323) );
  XOR2_X1 U377 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n321) );
  XNOR2_X1 U378 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n400) );
  XNOR2_X1 U380 ( .A(n400), .B(G36GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n335) );
  XOR2_X1 U382 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n325) );
  XNOR2_X1 U383 ( .A(G106GAT), .B(G85GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U385 ( .A(G99GAT), .B(n326), .ZN(n377) );
  XOR2_X1 U386 ( .A(KEYINPUT82), .B(G190GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(G43GAT), .B(G50GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U389 ( .A(n377), .B(n329), .Z(n333) );
  XOR2_X1 U390 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n331) );
  XNOR2_X1 U391 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n332) );
  INV_X1 U393 ( .A(n496), .ZN(n584) );
  XOR2_X1 U394 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n337) );
  XNOR2_X1 U395 ( .A(G8GAT), .B(KEYINPUT71), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n343) );
  INV_X1 U397 ( .A(KEYINPUT13), .ZN(n338) );
  NAND2_X1 U398 ( .A1(G71GAT), .A2(n338), .ZN(n357) );
  INV_X1 U399 ( .A(G71GAT), .ZN(n339) );
  NAND2_X1 U400 ( .A1(n339), .A2(KEYINPUT13), .ZN(n358) );
  NAND2_X1 U401 ( .A1(n357), .A2(n358), .ZN(n356) );
  XOR2_X1 U402 ( .A(KEYINPUT14), .B(n356), .Z(n341) );
  XOR2_X1 U403 ( .A(G127GAT), .B(G57GAT), .Z(n443) );
  XNOR2_X1 U404 ( .A(G15GAT), .B(n443), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U406 ( .A(n343), .B(n342), .Z(n345) );
  NAND2_X1 U407 ( .A1(G231GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U409 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n347) );
  XNOR2_X1 U410 ( .A(G1GAT), .B(KEYINPUT85), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U412 ( .A(n349), .B(n348), .Z(n354) );
  XOR2_X1 U413 ( .A(G64GAT), .B(KEYINPUT84), .Z(n351) );
  XNOR2_X1 U414 ( .A(G183GAT), .B(G211GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n433) );
  XNOR2_X1 U416 ( .A(n352), .B(n433), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n599) );
  XOR2_X1 U418 ( .A(n599), .B(KEYINPUT111), .Z(n582) );
  INV_X1 U419 ( .A(KEYINPUT74), .ZN(n355) );
  NAND2_X1 U420 ( .A1(n356), .A2(n355), .ZN(n361) );
  AND2_X1 U421 ( .A1(n357), .A2(KEYINPUT74), .ZN(n359) );
  NAND2_X1 U422 ( .A1(n359), .A2(n358), .ZN(n360) );
  NAND2_X1 U423 ( .A1(n361), .A2(n360), .ZN(n363) );
  NAND2_X1 U424 ( .A1(G230GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G148GAT), .Z(n444) );
  XNOR2_X1 U427 ( .A(n364), .B(n444), .ZN(n372) );
  XOR2_X1 U428 ( .A(G92GAT), .B(G204GAT), .Z(n366) );
  XNOR2_X1 U429 ( .A(G176GAT), .B(G78GAT), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U431 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n368) );
  XNOR2_X1 U432 ( .A(G57GAT), .B(G64GAT), .ZN(n367) );
  XNOR2_X1 U433 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U434 ( .A(n370), .B(n369), .Z(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U436 ( .A(KEYINPUT79), .B(KEYINPUT33), .Z(n374) );
  XNOR2_X1 U437 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n378) );
  NAND2_X1 U440 ( .A1(n378), .A2(n377), .ZN(n382) );
  INV_X1 U441 ( .A(n377), .ZN(n380) );
  INV_X1 U442 ( .A(n378), .ZN(n379) );
  NAND2_X1 U443 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U444 ( .A1(n382), .A2(n381), .ZN(n416) );
  XOR2_X1 U445 ( .A(n416), .B(KEYINPUT65), .Z(n383) );
  XOR2_X1 U446 ( .A(n383), .B(KEYINPUT41), .Z(n575) );
  INV_X1 U447 ( .A(n575), .ZN(n554) );
  XOR2_X1 U448 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n385) );
  XNOR2_X1 U449 ( .A(KEYINPUT72), .B(KEYINPUT30), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n405) );
  XNOR2_X1 U451 ( .A(G169GAT), .B(G36GAT), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n386), .B(G8GAT), .ZN(n387) );
  INV_X1 U453 ( .A(n387), .ZN(n438) );
  XOR2_X1 U454 ( .A(G43GAT), .B(G15GAT), .Z(n463) );
  NAND2_X1 U455 ( .A1(n438), .A2(n463), .ZN(n390) );
  INV_X1 U456 ( .A(n463), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n388), .A2(n387), .ZN(n389) );
  NAND2_X1 U458 ( .A1(n390), .A2(n389), .ZN(n394) );
  NAND2_X1 U459 ( .A1(G229GAT), .A2(G233GAT), .ZN(n391) );
  XOR2_X1 U460 ( .A(KEYINPUT71), .B(G22GAT), .Z(n396) );
  XNOR2_X1 U461 ( .A(G113GAT), .B(G197GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U463 ( .A(G29GAT), .B(G1GAT), .Z(n454) );
  XOR2_X1 U464 ( .A(n397), .B(n454), .Z(n398) );
  XNOR2_X1 U465 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U466 ( .A(n400), .B(KEYINPUT68), .Z(n401) );
  XOR2_X1 U467 ( .A(n405), .B(n404), .Z(n591) );
  NAND2_X1 U468 ( .A1(n554), .A2(n591), .ZN(n407) );
  XOR2_X1 U469 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  NOR2_X1 U471 ( .A1(n582), .A2(n408), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n409), .B(KEYINPUT113), .ZN(n410) );
  NOR2_X1 U473 ( .A1(n584), .A2(n410), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n413), .B(n412), .ZN(n421) );
  XOR2_X1 U475 ( .A(KEYINPUT73), .B(n591), .Z(n552) );
  XOR2_X1 U476 ( .A(n496), .B(KEYINPUT36), .Z(n601) );
  NAND2_X1 U477 ( .A1(n599), .A2(n601), .ZN(n415) );
  XNOR2_X1 U478 ( .A(KEYINPUT45), .B(KEYINPUT115), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n417) );
  BUF_X1 U480 ( .A(n416), .Z(n595) );
  NAND2_X1 U481 ( .A1(n417), .A2(n595), .ZN(n418) );
  NOR2_X1 U482 ( .A1(n552), .A2(n418), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n419), .B(KEYINPUT116), .ZN(n420) );
  XNOR2_X1 U484 ( .A(KEYINPUT64), .B(KEYINPUT117), .ZN(n422) );
  INV_X1 U485 ( .A(n563), .ZN(n548) );
  XNOR2_X1 U486 ( .A(KEYINPUT17), .B(KEYINPUT90), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(KEYINPUT91), .B(G190GAT), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n298), .B(n428), .ZN(n473) );
  XNOR2_X1 U490 ( .A(n473), .B(n429), .ZN(n436) );
  XOR2_X1 U491 ( .A(n430), .B(KEYINPUT96), .Z(n432) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U494 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n540) );
  XNOR2_X1 U497 ( .A(n540), .B(KEYINPUT121), .ZN(n439) );
  NOR2_X1 U498 ( .A1(n548), .A2(n439), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n440), .B(KEYINPUT54), .ZN(n460) );
  XNOR2_X1 U500 ( .A(G113GAT), .B(G134GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n441), .B(KEYINPUT0), .ZN(n462) );
  XNOR2_X1 U502 ( .A(n462), .B(n442), .ZN(n458) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n446) );
  NAND2_X1 U504 ( .A1(G225GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U506 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n448) );
  XNOR2_X1 U507 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U509 ( .A(n450), .B(n449), .Z(n456) );
  XOR2_X1 U510 ( .A(KEYINPUT1), .B(G85GAT), .Z(n452) );
  XNOR2_X1 U511 ( .A(G141GAT), .B(G155GAT), .ZN(n451) );
  XNOR2_X1 U512 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U514 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U515 ( .A(n458), .B(n457), .ZN(n492) );
  NAND2_X1 U516 ( .A1(n486), .A2(n590), .ZN(n461) );
  XOR2_X1 U517 ( .A(n463), .B(n462), .Z(n465) );
  NAND2_X1 U518 ( .A1(G227GAT), .A2(G233GAT), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n465), .B(n464), .ZN(n469) );
  XOR2_X1 U520 ( .A(G127GAT), .B(G183GAT), .Z(n467) );
  XNOR2_X1 U521 ( .A(G71GAT), .B(G120GAT), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U523 ( .A(n469), .B(n468), .Z(n475) );
  XOR2_X1 U524 ( .A(KEYINPUT20), .B(KEYINPUT89), .Z(n471) );
  XNOR2_X1 U525 ( .A(G169GAT), .B(G99GAT), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U528 ( .A(n475), .B(n474), .ZN(n550) );
  NAND2_X1 U529 ( .A1(n585), .A2(n552), .ZN(n478) );
  INV_X1 U530 ( .A(KEYINPUT122), .ZN(n477) );
  XNOR2_X1 U531 ( .A(n478), .B(n477), .ZN(n480) );
  INV_X1 U532 ( .A(G169GAT), .ZN(n479) );
  XNOR2_X1 U533 ( .A(n480), .B(n479), .ZN(G1348GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n502) );
  XOR2_X1 U535 ( .A(n550), .B(KEYINPUT92), .Z(n482) );
  XOR2_X1 U536 ( .A(n486), .B(KEYINPUT28), .Z(n544) );
  XNOR2_X1 U537 ( .A(n540), .B(KEYINPUT27), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n488), .A2(n538), .ZN(n481) );
  XOR2_X1 U539 ( .A(KEYINPUT97), .B(n481), .Z(n565) );
  NAND2_X1 U540 ( .A1(n482), .A2(n549), .ZN(n494) );
  NAND2_X1 U541 ( .A1(n550), .A2(n540), .ZN(n483) );
  NAND2_X1 U542 ( .A1(n483), .A2(n486), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT25), .B(n484), .Z(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT98), .ZN(n490) );
  NOR2_X1 U545 ( .A1(n486), .A2(n550), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n487), .B(KEYINPUT26), .ZN(n589) );
  NAND2_X1 U547 ( .A1(n488), .A2(n589), .ZN(n489) );
  NAND2_X1 U548 ( .A1(n490), .A2(n489), .ZN(n491) );
  NAND2_X1 U549 ( .A1(n492), .A2(n491), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U551 ( .A(n495), .B(KEYINPUT99), .ZN(n512) );
  XOR2_X1 U552 ( .A(KEYINPUT16), .B(KEYINPUT88), .Z(n498) );
  NAND2_X1 U553 ( .A1(n599), .A2(n496), .ZN(n497) );
  XOR2_X1 U554 ( .A(n498), .B(n497), .Z(n499) );
  NOR2_X1 U555 ( .A1(n512), .A2(n499), .ZN(n500) );
  XOR2_X1 U556 ( .A(KEYINPUT100), .B(n500), .Z(n525) );
  NAND2_X1 U557 ( .A1(n552), .A2(n595), .ZN(n515) );
  NOR2_X1 U558 ( .A1(n525), .A2(n515), .ZN(n509) );
  NAND2_X1 U559 ( .A1(n509), .A2(n538), .ZN(n501) );
  XNOR2_X1 U560 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n509), .A2(n540), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G8GAT), .B(n505), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n507) );
  NAND2_X1 U566 ( .A1(n509), .A2(n550), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U568 ( .A(G15GAT), .B(n508), .Z(G1326GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n544), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(KEYINPUT104), .ZN(n511) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(n511), .ZN(G1327GAT) );
  XOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT39), .Z(n518) );
  NOR2_X1 U573 ( .A1(n599), .A2(n512), .ZN(n513) );
  NAND2_X1 U574 ( .A1(n601), .A2(n297), .ZN(n514) );
  XOR2_X1 U575 ( .A(KEYINPUT37), .B(n514), .Z(n536) );
  NOR2_X1 U576 ( .A1(n536), .A2(n515), .ZN(n516) );
  XNOR2_X1 U577 ( .A(KEYINPUT38), .B(n516), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(n538), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n518), .B(n517), .ZN(G1328GAT) );
  NAND2_X1 U580 ( .A1(n522), .A2(n540), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U582 ( .A1(n522), .A2(n550), .ZN(n520) );
  XNOR2_X1 U583 ( .A(n520), .B(KEYINPUT40), .ZN(n521) );
  XNOR2_X1 U584 ( .A(G43GAT), .B(n521), .ZN(G1330GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n544), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U587 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n528) );
  NOR2_X1 U588 ( .A1(n591), .A2(n575), .ZN(n524) );
  XOR2_X1 U589 ( .A(KEYINPUT106), .B(n524), .Z(n537) );
  NOR2_X1 U590 ( .A1(n537), .A2(n525), .ZN(n526) );
  XOR2_X1 U591 ( .A(KEYINPUT107), .B(n526), .Z(n531) );
  NAND2_X1 U592 ( .A1(n531), .A2(n538), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1332GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n540), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n529), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U596 ( .A1(n531), .A2(n550), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n530), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n533) );
  NAND2_X1 U599 ( .A1(n531), .A2(n544), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U601 ( .A(G78GAT), .B(KEYINPUT108), .Z(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1335GAT) );
  NOR2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n545), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G85GAT), .B(n539), .ZN(G1336GAT) );
  NAND2_X1 U606 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n541), .B(KEYINPUT110), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G92GAT), .B(n542), .ZN(G1337GAT) );
  NAND2_X1 U609 ( .A1(n545), .A2(n550), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n546), .B(KEYINPUT44), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G106GAT), .B(n547), .ZN(G1339GAT) );
  NAND2_X1 U614 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U615 ( .A1(n548), .A2(n551), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n559), .A2(n552), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U618 ( .A(G120GAT), .B(KEYINPUT49), .Z(n556) );
  NAND2_X1 U619 ( .A1(n559), .A2(n554), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n556), .B(n555), .ZN(G1341GAT) );
  NAND2_X1 U621 ( .A1(n559), .A2(n582), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(KEYINPUT50), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G127GAT), .B(n558), .ZN(G1342GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n561) );
  NAND2_X1 U625 ( .A1(n559), .A2(n584), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(G134GAT), .B(n562), .ZN(G1343GAT) );
  XOR2_X1 U628 ( .A(G141GAT), .B(KEYINPUT119), .Z(n567) );
  NAND2_X1 U629 ( .A1(n563), .A2(n589), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n572), .A2(n591), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1344GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n569) );
  NAND2_X1 U634 ( .A1(n572), .A2(n554), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G148GAT), .B(n570), .ZN(G1345GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n599), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U639 ( .A1(n572), .A2(n584), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(KEYINPUT120), .ZN(n574) );
  XNOR2_X1 U641 ( .A(G162GAT), .B(n574), .ZN(G1347GAT) );
  INV_X1 U642 ( .A(n585), .ZN(n581) );
  NOR2_X1 U643 ( .A1(n575), .A2(n581), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n577) );
  XNOR2_X1 U645 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U647 ( .A(KEYINPUT56), .B(n578), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n580), .B(n579), .ZN(G1349GAT) );
  NAND2_X1 U649 ( .A1(n585), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n583), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n587) );
  XOR2_X1 U652 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n586) );
  XNOR2_X1 U653 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(G190GAT), .ZN(G1351GAT) );
  AND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n602) );
  NAND2_X1 U656 ( .A1(n602), .A2(n591), .ZN(n594) );
  XOR2_X1 U657 ( .A(G197GAT), .B(KEYINPUT60), .Z(n592) );
  XNOR2_X1 U658 ( .A(KEYINPUT59), .B(n592), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n594), .B(n593), .ZN(G1352GAT) );
  XOR2_X1 U660 ( .A(G204GAT), .B(KEYINPUT61), .Z(n598) );
  INV_X1 U661 ( .A(n595), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n602), .A2(n596), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n598), .B(n597), .ZN(G1353GAT) );
  NAND2_X1 U664 ( .A1(n602), .A2(n599), .ZN(n600) );
  XNOR2_X1 U665 ( .A(n600), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U666 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n606) );
  XOR2_X1 U667 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n604) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n604), .B(n603), .ZN(n605) );
  XNOR2_X1 U670 ( .A(n606), .B(n605), .ZN(G1355GAT) );
endmodule

