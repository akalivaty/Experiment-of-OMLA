//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n591, new_n592, new_n593, new_n594, new_n595, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n470), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT66), .B1(new_n470), .B2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G101), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n466), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  INV_X1    g053(.A(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n470), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n470), .B2(G112), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n488), .B1(new_n482), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n493), .B2(G124), .ZN(G162));
  NAND3_X1  g069(.A1(KEYINPUT68), .A2(KEYINPUT4), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n480), .B2(new_n481), .ZN(new_n496));
  AND2_X1   g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n470), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n480), .B2(new_n481), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g078(.A(G138), .B(new_n470), .C1(new_n464), .C2(new_n465), .ZN(new_n504));
  XOR2_X1   g079(.A(KEYINPUT68), .B(KEYINPUT4), .Z(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n516), .A2(new_n518), .A3(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n514), .A2(G651), .B1(new_n519), .B2(G50), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n516), .B(new_n518), .C1(new_n510), .C2(new_n511), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT69), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT70), .B(G88), .Z(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT71), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n520), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n519), .A2(G51), .ZN(new_n535));
  XNOR2_X1  g110(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n534), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n522), .A2(G89), .A3(new_n526), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G64), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n512), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G651), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n522), .A2(G90), .A3(new_n526), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n519), .A2(G52), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(KEYINPUT73), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT73), .B1(new_n548), .B2(new_n549), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AND2_X1   g129(.A1(new_n522), .A2(new_n526), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G81), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n512), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n559), .A2(G651), .B1(new_n519), .B2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n522), .A2(G91), .A3(new_n526), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n512), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n516), .A2(new_n518), .A3(G53), .A4(G543), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n577));
  AND3_X1   g152(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT74), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT74), .B1(new_n576), .B2(new_n577), .ZN(new_n579));
  NOR3_X1   g154(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n576), .A2(new_n577), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n576), .A2(new_n577), .A3(KEYINPUT74), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n585), .A2(new_n586), .A3(new_n572), .A4(new_n568), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n588), .ZN(G299));
  INV_X1    g164(.A(G168), .ZN(G286));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  INV_X1    g166(.A(new_n532), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n531), .B1(new_n520), .B2(new_n528), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n532), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G303));
  NAND2_X1  g171(.A1(new_n555), .A2(G87), .ZN(new_n597));
  OAI21_X1  g172(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n519), .A2(G49), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(G288));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n517), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n522), .A2(G86), .A3(new_n526), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n519), .A2(G48), .ZN(new_n607));
  OAI21_X1  g182(.A(G61), .B1(new_n510), .B2(new_n511), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n610), .A2(KEYINPUT78), .A3(G651), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n605), .A2(new_n606), .A3(new_n607), .A4(new_n611), .ZN(G305));
  NAND2_X1  g187(.A1(new_n555), .A2(G85), .ZN(new_n613));
  NAND2_X1  g188(.A1(G72), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G60), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n512), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(new_n519), .B2(G47), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n519), .A2(G54), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n517), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n555), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n522), .A2(new_n526), .ZN(new_n625));
  INV_X1    g200(.A(G92), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n622), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n619), .B1(G868), .B2(new_n628), .ZN(G284));
  OAI21_X1  g204(.A(new_n619), .B1(G868), .B2(new_n628), .ZN(G321));
  INV_X1    g205(.A(G868), .ZN(new_n631));
  MUX2_X1   g206(.A(G286), .B(G299), .S(new_n631), .Z(G280));
  XOR2_X1   g207(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n628), .B1(new_n634), .B2(G860), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g211(.A1(new_n628), .A2(new_n634), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g215(.A(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n470), .B2(G111), .ZN(new_n643));
  OAI22_X1  g218(.A1(new_n483), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n493), .B2(G123), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(KEYINPUT82), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(KEYINPUT82), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n482), .B1(new_n471), .B2(new_n472), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n650), .A2(new_n655), .ZN(G156));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT84), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2443), .B(G2446), .Z(new_n668));
  XNOR2_X1  g243(.A(G2451), .B(G2454), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n667), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n671), .A2(G14), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT85), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  INV_X1    g250(.A(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2084), .B(G2090), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2067), .B(G2678), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2072), .B(G2078), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(KEYINPUT17), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n678), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(new_n677), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT18), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n678), .A2(new_n677), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n683), .B(new_n686), .C1(new_n681), .C2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT87), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n649), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n649), .B1(new_n690), .B2(new_n691), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n676), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n696), .A2(G2100), .A3(new_n692), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1956), .B(G2474), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1961), .B(G1966), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT20), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n701), .B(new_n702), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n700), .B1(KEYINPUT88), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT88), .B2(new_n707), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  INV_X1    g286(.A(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n710), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT89), .B(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G229));
  MUX2_X1   g293(.A(G6), .B(G305), .S(G16), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT32), .B(G1981), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G23), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT92), .Z(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(G288), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT33), .B(G1976), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(G22), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G166), .B2(new_n726), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1971), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G1971), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n729), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OR3_X1    g309(.A1(new_n723), .A2(KEYINPUT34), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT34), .B1(new_n723), .B2(new_n734), .ZN(new_n736));
  MUX2_X1   g311(.A(G24), .B(G290), .S(G16), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR3_X1   g317(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n743));
  OAI221_X1 g318(.A(G2104), .B1(G107), .B2(new_n470), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G131), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n483), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(new_n493), .B2(G119), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n740), .B1(new_n747), .B2(new_n739), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT35), .B(G1991), .Z(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n748), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n738), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n735), .A2(new_n736), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT36), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT36), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n735), .A2(new_n755), .A3(new_n736), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(KEYINPUT24), .B2(G34), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n476), .B2(G29), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  OAI21_X1  g339(.A(G105), .B1(new_n471), .B2(new_n472), .ZN(new_n765));
  INV_X1    g340(.A(G141), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n483), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n493), .B2(G129), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n768), .A2(new_n739), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n739), .B2(G32), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT27), .B(G1996), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n726), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n726), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n762), .B1(new_n770), .B2(new_n771), .C1(G1961), .C2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT99), .Z(new_n775));
  NAND2_X1  g350(.A1(G168), .A2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G16), .B2(G21), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n773), .A2(G1961), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n760), .A2(new_n761), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n739), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  NOR2_X1   g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT94), .Z(new_n787));
  INV_X1    g362(.A(G116), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n479), .B1(new_n788), .B2(G2105), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n787), .A2(new_n789), .B1(new_n474), .B2(G140), .ZN(new_n790));
  INV_X1    g365(.A(G128), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n492), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n785), .B1(new_n792), .B2(G29), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2067), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n646), .A2(G29), .A3(new_n647), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n783), .B(new_n794), .C1(KEYINPUT98), .C2(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n780), .A2(new_n781), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n739), .A2(G33), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G139), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n483), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n482), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(new_n470), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT95), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n798), .B1(new_n807), .B2(new_n739), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(G2072), .Z(new_n809));
  INV_X1    g384(.A(G19), .ZN(new_n810));
  OR3_X1    g385(.A1(new_n810), .A2(KEYINPUT93), .A3(G16), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT93), .B1(new_n810), .B2(G16), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n811), .B(new_n812), .C1(new_n562), .C2(new_n726), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1341), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n739), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n739), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT29), .Z(new_n819));
  INV_X1    g394(.A(G2090), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n739), .A2(G27), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G164), .B2(new_n739), .ZN(new_n823));
  INV_X1    g398(.A(G2078), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n770), .A2(new_n771), .ZN(new_n826));
  INV_X1    g401(.A(G28), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(KEYINPUT30), .ZN(new_n828));
  AOI21_X1  g403(.A(G29), .B1(new_n827), .B2(KEYINPUT30), .ZN(new_n829));
  OR2_X1    g404(.A1(KEYINPUT31), .A2(G11), .ZN(new_n830));
  NAND2_X1  g405(.A1(KEYINPUT31), .A2(G11), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n828), .A2(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n821), .A2(new_n825), .A3(new_n826), .A4(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n726), .A2(G4), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n628), .B2(new_n726), .ZN(new_n835));
  INV_X1    g410(.A(G1348), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n819), .B2(new_n820), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n816), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n726), .A2(G20), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT23), .Z(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G299), .B2(G16), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G1956), .ZN(new_n843));
  AND4_X1   g418(.A1(new_n775), .A2(new_n797), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n757), .A2(KEYINPUT100), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT100), .B1(new_n757), .B2(new_n844), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(G311));
  NAND2_X1  g422(.A1(new_n757), .A2(new_n844), .ZN(G150));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n512), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n519), .A2(G55), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n852), .B(new_n853), .C1(new_n625), .C2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n561), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n628), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n862), .A3(G860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(G860), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  NAND2_X1  g441(.A1(new_n474), .A2(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(new_n470), .B2(G118), .ZN(new_n869));
  INV_X1    g444(.A(G130), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n867), .B1(new_n868), .B2(new_n869), .C1(new_n492), .C2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(new_n768), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n807), .A2(new_n507), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n807), .A2(new_n507), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n792), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n807), .A2(new_n507), .ZN(new_n877));
  INV_X1    g452(.A(new_n792), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n807), .A2(new_n507), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G119), .ZN(new_n881));
  OAI221_X1 g456(.A(new_n744), .B1(new_n745), .B2(new_n483), .C1(new_n492), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT101), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n747), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n652), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n885), .A3(new_n652), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n876), .A2(new_n880), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n876), .B2(new_n880), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n873), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n876), .A2(new_n880), .ZN(new_n894));
  INV_X1    g469(.A(new_n890), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n876), .A2(new_n880), .A3(new_n890), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n872), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n648), .B(new_n476), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G162), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n893), .A3(new_n898), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g482(.A(new_n857), .B(new_n637), .ZN(new_n908));
  INV_X1    g483(.A(new_n628), .ZN(new_n909));
  NAND2_X1  g484(.A1(G299), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n582), .A2(new_n588), .A3(new_n628), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT102), .Z(new_n914));
  INV_X1    g489(.A(new_n911), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n628), .B1(new_n582), .B2(new_n588), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT41), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n910), .A2(new_n918), .A3(new_n911), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT103), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n912), .A2(new_n921), .A3(KEYINPUT41), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n908), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n914), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(G166), .B(G290), .ZN(new_n926));
  XOR2_X1   g501(.A(G288), .B(G305), .Z(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT42), .Z(new_n929));
  AND2_X1   g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n913), .B(KEYINPUT102), .ZN(new_n931));
  INV_X1    g506(.A(new_n923), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT104), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n925), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n855), .A2(new_n631), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n917), .A2(new_n919), .ZN(new_n940));
  NAND2_X1  g515(.A1(G301), .A2(G286), .ZN(new_n941));
  OAI211_X1 g516(.A(G168), .B(new_n547), .C1(new_n551), .C2(new_n552), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n561), .B(new_n855), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n857), .A2(new_n941), .A3(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n940), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT105), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n943), .A2(KEYINPUT105), .A3(new_n944), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(new_n912), .ZN(new_n952));
  INV_X1    g527(.A(new_n928), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n920), .A2(new_n949), .A3(new_n922), .A4(new_n950), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n956));
  OR3_X1    g531(.A1(new_n947), .A2(new_n956), .A3(new_n912), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n947), .B2(new_n912), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n955), .A2(new_n957), .A3(new_n928), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n939), .B1(new_n961), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n953), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n904), .A3(new_n959), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(KEYINPUT43), .B1(new_n963), .B2(new_n954), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n939), .B2(new_n970), .ZN(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n507), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n469), .A2(new_n475), .A3(G40), .A4(new_n473), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n792), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n979), .B2(new_n768), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT125), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n981), .A2(KEYINPUT47), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n977), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n768), .B(G1996), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n979), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n882), .A2(new_n750), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n747), .A2(new_n749), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n976), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n988), .A2(KEYINPUT48), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n989), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n991), .A2(new_n993), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n978), .B2(new_n878), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n999), .B2(new_n977), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT47), .B1(new_n981), .B2(new_n984), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n985), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G8), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n1005));
  INV_X1    g580(.A(G137), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n473), .B1(new_n483), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n482), .A2(G125), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n470), .B1(new_n1008), .B2(new_n463), .ZN(new_n1009));
  INV_X1    g584(.A(G40), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1005), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1004), .B1(new_n1012), .B2(new_n973), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n507), .A2(new_n972), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n975), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n507), .A2(new_n1016), .A3(new_n972), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT108), .B(G2090), .Z(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1003), .B1(new_n1013), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n592), .A2(new_n593), .A3(new_n591), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT76), .B1(new_n530), .B2(new_n532), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1024), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G303), .A2(G8), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1020), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT63), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n779), .B1(new_n1012), .B2(new_n973), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1015), .A2(new_n761), .A3(new_n1017), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT110), .B(G8), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(G168), .A3(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1028), .A2(new_n1029), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G305), .B2(G1981), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n606), .A2(new_n607), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT78), .B1(new_n610), .B2(G651), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n603), .B(new_n517), .C1(new_n608), .C2(new_n609), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1039), .A2(KEYINPUT111), .A3(new_n1042), .A4(new_n712), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G305), .A2(G1981), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT49), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1044), .A2(KEYINPUT112), .A3(KEYINPUT49), .A4(new_n1045), .ZN(new_n1052));
  OAI21_X1  g627(.A(G126), .B1(new_n464), .B2(new_n465), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n501), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(G2105), .B1(new_n504), .B2(new_n505), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1384), .B1(new_n1055), .B2(new_n498), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1033), .B1(new_n1011), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .A4(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1060), .B(new_n1057), .C1(new_n1059), .C2(G288), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1057), .B1(new_n1059), .B2(G288), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1025), .A2(new_n1027), .A3(new_n1020), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1036), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n1034), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1026), .B1(G303), .B2(G8), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1003), .B(new_n1024), .C1(new_n594), .C2(new_n595), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1058), .A2(new_n1073), .A3(new_n1066), .A4(new_n1064), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1068), .B1(new_n1074), .B2(new_n1035), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1029), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n1074), .A2(new_n1068), .A3(new_n1035), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1067), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1012), .A2(G2078), .A3(new_n973), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT53), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(KEYINPUT53), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1011), .A3(new_n1017), .ZN(new_n1083));
  INV_X1    g658(.A(G1961), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1032), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1033), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1003), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G168), .A2(new_n1033), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1092), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1093), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1095), .B1(new_n1096), .B2(new_n1089), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1087), .B1(new_n1097), .B2(KEYINPUT62), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1096), .A2(new_n1089), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1092), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1098), .A2(new_n1099), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G288), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1058), .A2(new_n1059), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1044), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1066), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1109), .A2(new_n1057), .B1(new_n1110), .B2(new_n1065), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1078), .A2(new_n1106), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1087), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1086), .A2(G171), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1114), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(new_n1087), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(new_n1099), .A3(new_n1105), .A4(new_n1097), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n562), .A2(KEYINPUT119), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1012), .A2(new_n973), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n982), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT117), .B1(new_n1014), .B2(new_n975), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1011), .A2(new_n1056), .A3(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(KEYINPUT58), .B(G1341), .Z(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1121), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n1121), .C1(new_n1123), .C2(new_n1128), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1122), .A2(new_n1133), .B1(new_n1083), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n573), .A2(KEYINPUT114), .ZN(new_n1136));
  INV_X1    g711(.A(new_n583), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT114), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n568), .A2(new_n1138), .A3(new_n572), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n580), .B2(KEYINPUT57), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n587), .A2(KEYINPUT115), .A3(new_n1141), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT61), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1083), .A2(new_n1134), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n974), .A2(new_n1011), .A3(new_n1005), .A4(new_n1133), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n573), .A2(new_n579), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1151), .A2(new_n1143), .A3(KEYINPUT57), .A4(new_n586), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT115), .B1(new_n587), .B2(new_n1141), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(new_n1153), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1131), .A2(new_n1132), .B1(new_n1147), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n628), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(G2067), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1348), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1014), .A2(new_n975), .A3(KEYINPUT117), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1125), .B1(new_n1011), .B2(new_n1056), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n978), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1011), .B1(new_n1056), .B2(new_n1016), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1017), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n836), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT118), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1159), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n628), .A2(new_n1158), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1171), .A2(new_n1172), .B1(new_n1173), .B2(new_n1157), .ZN(new_n1174));
  OAI221_X1 g749(.A(new_n1159), .B1(new_n1158), .B2(new_n628), .C1(new_n1163), .C2(new_n1170), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1156), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1150), .A2(new_n1154), .A3(KEYINPUT116), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT116), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1182), .B1(new_n1135), .B2(new_n1146), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1150), .A2(KEYINPUT120), .A3(new_n1154), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1177), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT121), .B(new_n1177), .C1(new_n1181), .C2(new_n1185), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1176), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  AOI22_X1  g765(.A1(new_n1173), .A2(new_n628), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(new_n1181), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1120), .B1(new_n1193), .B2(KEYINPUT123), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1190), .A2(new_n1195), .A3(new_n1192), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1112), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(G290), .A2(G1986), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n987), .A2(KEYINPUT107), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT107), .ZN(new_n1200));
  NAND3_X1  g775(.A1(G290), .A2(new_n1200), .A3(G1986), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1199), .A2(new_n976), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n995), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1002), .B1(new_n1197), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(G229), .A2(new_n461), .ZN(new_n1206));
  NAND4_X1  g780(.A1(new_n1206), .A2(new_n674), .A3(new_n697), .A4(new_n695), .ZN(new_n1207));
  INV_X1    g781(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n906), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g783(.A(KEYINPUT126), .B1(new_n970), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(G37), .B1(new_n899), .B2(new_n902), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1207), .B1(new_n1211), .B2(new_n905), .ZN(new_n1212));
  INV_X1    g786(.A(KEYINPUT126), .ZN(new_n1213));
  AND2_X1   g787(.A1(new_n963), .A2(new_n954), .ZN(new_n1214));
  AOI21_X1  g788(.A(new_n962), .B1(new_n965), .B2(new_n959), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n1212), .B(new_n1213), .C1(new_n1214), .C2(new_n1215), .ZN(new_n1216));
  AND2_X1   g790(.A1(new_n1210), .A2(new_n1216), .ZN(G308));
  OAI21_X1  g791(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(G225));
endmodule


