//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT27), .B(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT28), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT27), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G183gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n206), .B(new_n204), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n213), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G183gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n207), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n206), .B1(new_n219), .B2(new_n204), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n205), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(new_n223), .B2(new_n224), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n222), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT71), .B(G120gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT72), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(G113gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G113gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n233), .B1(new_n238), .B2(G120gat), .ZN(new_n239));
  INV_X1    g038(.A(new_n232), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n238), .ZN(new_n241));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT1), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(new_n243), .B2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n236), .B(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n237), .A2(new_n241), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(KEYINPUT24), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G183gat), .B2(G190gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n208), .A2(new_n204), .A3(KEYINPUT64), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G169gat), .ZN(new_n258));
  INV_X1    g057(.A(G176gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT65), .A4(KEYINPUT23), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT23), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(G169gat), .B2(G176gat), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n260), .A2(new_n227), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n227), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n270), .A3(new_n227), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(KEYINPUT25), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n218), .A2(new_n204), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n274), .B2(new_n253), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n249), .A2(new_n267), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n231), .A2(new_n248), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT73), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n221), .B2(new_n230), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n248), .ZN(new_n282));
  INV_X1    g081(.A(new_n248), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n219), .A2(new_n204), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT68), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(new_n215), .A3(new_n214), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n229), .B1(new_n286), .B2(new_n205), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n283), .B1(new_n287), .B2(new_n276), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n279), .A2(new_n282), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n290));
  AND2_X1   g089(.A1(G227gat), .A2(G233gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT32), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n292), .B2(new_n293), .ZN(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(KEYINPUT75), .ZN(new_n298));
  XOR2_X1   g097(.A(G71gat), .B(G99gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT34), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n295), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n303), .B2(new_n300), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT32), .B(new_n305), .C1(new_n292), .C2(new_n293), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n302), .B1(new_n301), .B2(new_n306), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n289), .A2(new_n291), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n301), .A2(new_n306), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT34), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n310), .B1(new_n314), .B2(new_n307), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n202), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n311), .B1(new_n308), .B2(new_n309), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n310), .A3(new_n307), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT36), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G141gat), .B(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n322), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n326), .B(new_n325), .C1(new_n321), .C2(KEYINPUT2), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT29), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT77), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT22), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n333), .A2(new_n334), .B1(G211gat), .B2(G218gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n333), .B2(new_n334), .ZN(new_n336));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G211gat), .B(G218gat), .Z(new_n340));
  OAI21_X1  g139(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n331), .B1(new_n342), .B2(KEYINPUT3), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n338), .B(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT79), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n329), .A2(new_n330), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n332), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n343), .B1(new_n352), .B2(KEYINPUT85), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n347), .A2(KEYINPUT85), .A3(new_n350), .ZN(new_n354));
  INV_X1    g153(.A(G228gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  OAI22_X1  g155(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G22gat), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n351), .A2(KEYINPUT86), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(KEYINPUT86), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n348), .B1(new_n346), .B2(KEYINPUT29), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n355), .B(new_n356), .C1(new_n361), .C2(new_n331), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n357), .A2(new_n358), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n357), .A2(new_n363), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G22gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n364), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n370), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n245), .A2(new_n247), .ZN(new_n376));
  INV_X1    g175(.A(new_n331), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n241), .A2(new_n235), .A3(new_n234), .A4(new_n236), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n331), .A2(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n349), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n379), .B(KEYINPUT4), .C1(new_n382), .C2(new_n248), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n386), .A2(KEYINPUT39), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n386), .B(KEYINPUT39), .C1(new_n385), .C2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G1gat), .B(G29gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(KEYINPUT0), .ZN(new_n393));
  XNOR2_X1  g192(.A(G57gat), .B(G85gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n395), .B(KEYINPUT89), .Z(new_n396));
  NAND3_X1  g195(.A1(new_n387), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT40), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT90), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n385), .B1(new_n380), .B2(new_n383), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT84), .B(new_n385), .C1(new_n388), .C2(new_n389), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n401), .A2(new_n404), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n396), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n397), .B2(new_n398), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT80), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n414), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n287), .B2(new_n276), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n347), .ZN(new_n418));
  INV_X1    g217(.A(new_n347), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n415), .A3(new_n416), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(KEYINPUT81), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n419), .A2(new_n415), .A3(new_n422), .A4(new_n416), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND4_X1  g227(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT30), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  AOI211_X1 g230(.A(new_n430), .B(new_n431), .C1(new_n421), .C2(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n423), .A3(new_n431), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT82), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n429), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n431), .B1(new_n421), .B2(new_n423), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT30), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(KEYINPUT88), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT88), .B1(new_n435), .B2(new_n437), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n400), .B(new_n411), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n405), .A2(new_n406), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(KEYINPUT5), .A3(new_n403), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n409), .B1(new_n443), .B2(new_n401), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n445));
  INV_X1    g244(.A(new_n395), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT6), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n444), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n410), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n395), .B1(new_n408), .B2(new_n409), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n451), .B2(KEYINPUT6), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n450), .A2(new_n452), .A3(new_n436), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n431), .A2(KEYINPUT37), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456));
  XOR2_X1   g255(.A(KEYINPUT91), .B(KEYINPUT38), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n418), .A2(new_n420), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT37), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n455), .A2(new_n456), .A3(new_n460), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n455), .A2(new_n460), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT92), .ZN(new_n464));
  INV_X1    g263(.A(new_n424), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n465), .A2(KEYINPUT37), .B1(new_n433), .B2(new_n454), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT94), .B1(new_n466), .B2(new_n457), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n455), .B1(new_n468), .B2(new_n424), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT94), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(new_n470), .A3(new_n458), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n462), .A2(new_n464), .A3(new_n467), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n375), .B1(new_n441), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n435), .A2(KEYINPUT83), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n451), .A2(KEYINPUT6), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n449), .B2(new_n451), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n437), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n374), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n320), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n374), .A2(new_n318), .A3(new_n317), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT35), .B1(new_n482), .B2(new_n479), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n312), .A2(new_n315), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n439), .A2(new_n440), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n450), .A2(new_n452), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT35), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n484), .A2(new_n374), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n481), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G57gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G64gat), .ZN(new_n492));
  INV_X1    g291(.A(G64gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G57gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(G71gat), .B(G78gat), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT101), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n492), .B2(new_n494), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT101), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n496), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT100), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n501), .B2(new_n496), .ZN(new_n505));
  AND2_X1   g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(G71gat), .A2(G78gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n508), .B(KEYINPUT100), .C1(new_n509), .C2(new_n497), .ZN(new_n510));
  AOI22_X1  g309(.A1(new_n500), .A2(new_n503), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g311(.A1(G231gat), .A2(G233gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G127gat), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G8gat), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(KEYINPUT21), .B2(new_n511), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n516), .B2(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n323), .ZN(new_n530));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n526), .A2(new_n527), .A3(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G190gat), .B(G218gat), .Z(new_n537));
  NAND2_X1  g336(.A1(G85gat), .A2(G92gat), .ZN(new_n538));
  OR2_X1    g337(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n539));
  AND3_X1   g338(.A1(KEYINPUT102), .A2(KEYINPUT103), .A3(KEYINPUT7), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT103), .B1(KEYINPUT102), .B2(KEYINPUT7), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n538), .B1(KEYINPUT102), .B2(KEYINPUT7), .ZN(new_n543));
  NAND2_X1  g342(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT103), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT102), .A2(KEYINPUT103), .A3(KEYINPUT7), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n542), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT8), .ZN(new_n551));
  OAI22_X1  g350(.A1(new_n550), .A2(new_n551), .B1(G85gat), .B2(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(G99gat), .A2(G106gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n549), .A2(new_n558), .A3(new_n553), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT17), .ZN(new_n562));
  AND2_X1   g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G43gat), .A2(G50gat), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT15), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(G29gat), .ZN(new_n568));
  INV_X1    g367(.A(G36gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT14), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G29gat), .A2(G36gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G43gat), .B(G50gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(new_n573), .B2(KEYINPUT15), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n565), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n570), .A2(new_n567), .A3(KEYINPUT95), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n572), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT95), .B1(new_n570), .B2(new_n567), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(KEYINPUT96), .B(new_n576), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n562), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n562), .A3(new_n583), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n561), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n537), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR3_X1   g397(.A1(new_n587), .A2(new_n592), .A3(new_n537), .ZN(new_n599));
  OR3_X1    g398(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n594), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n536), .A2(KEYINPUT104), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT104), .B1(new_n536), .B2(new_n602), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n523), .ZN(new_n610));
  INV_X1    g409(.A(new_n586), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n611), .B2(new_n584), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n588), .B2(new_n523), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n613), .B(new_n610), .C1(new_n611), .C2(new_n584), .ZN(new_n616));
  AOI211_X1 g415(.A(new_n607), .B(new_n609), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n610), .B(new_n588), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n608), .B(KEYINPUT13), .Z(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT98), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n523), .B1(new_n585), .B2(new_n586), .ZN(new_n623));
  INV_X1    g422(.A(new_n614), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n616), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n608), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n607), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(KEYINPUT18), .A3(new_n608), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  INV_X1    g428(.A(new_n621), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n622), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G197gat), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT11), .B(G169gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n628), .A2(new_n630), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n621), .B1(new_n640), .B2(KEYINPUT18), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n644), .A2(new_n627), .A3(KEYINPUT99), .A4(new_n637), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n632), .A2(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n505), .A2(new_n510), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n501), .A2(new_n502), .A3(new_n496), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n502), .B1(new_n501), .B2(new_n496), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n558), .B1(new_n549), .B2(new_n553), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n556), .B(new_n552), .C1(new_n542), .C2(new_n548), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n648), .A2(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n511), .A2(new_n557), .A3(new_n559), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(new_n655), .A3(KEYINPUT105), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n511), .A2(new_n557), .A3(new_n657), .A4(new_n559), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(KEYINPUT106), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n655), .A2(new_n660), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT10), .B1(new_n656), .B2(new_n658), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT106), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n647), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT107), .ZN(new_n668));
  INV_X1    g467(.A(new_n647), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n659), .A2(new_n660), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n662), .B1(new_n665), .B2(KEYINPUT106), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n647), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n668), .A2(new_n676), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n680), .B(KEYINPUT108), .Z(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n674), .B2(new_n677), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n606), .A2(new_n646), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n490), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n490), .A2(KEYINPUT110), .A3(new_n691), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n477), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(G1gat), .ZN(G1324gat));
  INV_X1    g498(.A(new_n485), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n696), .A2(KEYINPUT42), .A3(new_n700), .A4(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n696), .A2(new_n700), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(G8gat), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n706), .B2(G8gat), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n704), .B(new_n705), .C1(new_n708), .C2(new_n709), .ZN(G1325gat));
  INV_X1    g509(.A(G15gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n711), .A3(new_n484), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT36), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT36), .B1(new_n317), .B2(new_n318), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n316), .A2(KEYINPUT112), .A3(new_n319), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n694), .B2(new_n695), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n712), .B1(new_n720), .B2(new_n711), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n696), .A2(new_n375), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n400), .A2(new_n411), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n435), .A2(new_n437), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT88), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n438), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n467), .A2(new_n471), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n453), .A2(new_n464), .A3(new_n461), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n374), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n479), .A2(new_n374), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(new_n717), .A3(new_n716), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n489), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n738));
  INV_X1    g537(.A(new_n602), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI22_X1  g539(.A1(new_n735), .A2(new_n320), .B1(new_n483), .B2(new_n488), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n741), .B2(new_n602), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n690), .A2(new_n646), .A3(new_n536), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G29gat), .B1(new_n745), .B2(new_n477), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n490), .A2(new_n739), .A3(new_n744), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n697), .A2(new_n568), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n752));
  AND3_X1   g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n746), .B1(new_n753), .B2(new_n754), .ZN(G1328gat));
  NOR3_X1   g554(.A1(new_n747), .A2(G36gat), .A3(new_n485), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT46), .ZN(new_n757));
  OAI21_X1  g556(.A(G36gat), .B1(new_n745), .B2(new_n485), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(G1329gat));
  INV_X1    g558(.A(new_n484), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n747), .A2(G43gat), .A3(new_n760), .ZN(new_n761));
  AOI211_X1 g560(.A(KEYINPUT44), .B(new_n602), .C1(new_n736), .C2(new_n489), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n738), .B1(new_n490), .B2(new_n739), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n718), .B(new_n744), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(G43gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g566(.A(KEYINPUT47), .B(new_n761), .C1(new_n764), .C2(G43gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1330gat));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n375), .A2(G50gat), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n743), .A2(new_n744), .A3(new_n771), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n747), .A2(KEYINPUT115), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n374), .B1(new_n747), .B2(KEYINPUT115), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n770), .B(new_n772), .C1(new_n775), .C2(G50gat), .ZN(new_n776));
  INV_X1    g575(.A(new_n772), .ZN(new_n777));
  AOI21_X1  g576(.A(G50gat), .B1(new_n773), .B2(new_n774), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT48), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n776), .A2(new_n779), .ZN(G1331gat));
  NAND2_X1  g579(.A1(new_n632), .A2(new_n638), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n643), .A2(new_n645), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n690), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n606), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n737), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n477), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(new_n491), .ZN(G1332gat));
  NOR2_X1   g587(.A1(new_n786), .A2(new_n485), .ZN(new_n789));
  NOR2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  AND2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n792), .B1(new_n789), .B2(new_n790), .ZN(G1333gat));
  INV_X1    g592(.A(new_n786), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(G71gat), .A3(new_n718), .ZN(new_n795));
  INV_X1    g594(.A(G71gat), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n484), .B(KEYINPUT116), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n786), .B2(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n799), .B(new_n800), .ZN(G1334gat));
  NAND2_X1  g600(.A1(new_n794), .A2(new_n375), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g602(.A1(new_n783), .A2(new_n536), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n737), .A2(new_n739), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n602), .B1(new_n736), .B2(new_n489), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n808), .A2(KEYINPUT51), .A3(new_n804), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n784), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(G85gat), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n697), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n804), .A2(new_n690), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n743), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815), .B2(new_n477), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(G1336gat));
  NOR2_X1   g616(.A1(new_n485), .A2(G92gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI211_X1 g618(.A(new_n784), .B(new_n819), .C1(new_n807), .C2(new_n809), .ZN(new_n820));
  INV_X1    g619(.A(G92gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n813), .B1(new_n740), .B2(new_n742), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n700), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G92gat), .B1(new_n815), .B2(new_n485), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826));
  AND4_X1   g625(.A1(KEYINPUT51), .A2(new_n737), .A3(new_n739), .A4(new_n804), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT51), .B1(new_n808), .B2(new_n804), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n690), .B(new_n818), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n824), .A2(new_n830), .ZN(G1337gat));
  INV_X1    g630(.A(G99gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n832), .A3(new_n484), .ZN(new_n833));
  OAI21_X1  g632(.A(G99gat), .B1(new_n815), .B2(new_n719), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1338gat));
  OAI211_X1 g634(.A(new_n375), .B(new_n814), .C1(new_n762), .C2(new_n763), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n374), .A2(G106gat), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n690), .B(new_n838), .C1(new_n827), .C2(new_n828), .ZN(new_n839));
  XNOR2_X1  g638(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(G1339gat));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI211_X1 g643(.A(new_n671), .B(KEYINPUT10), .C1(new_n656), .C2(new_n658), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n666), .A2(new_n845), .A3(new_n662), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n669), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n668), .A3(new_n676), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n680), .B1(new_n674), .B2(new_n844), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n683), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n848), .B2(new_n849), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n646), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n618), .A2(new_n620), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n625), .B2(new_n608), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n636), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n782), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n688), .B2(new_n689), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n602), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n851), .A2(new_n857), .A3(new_n852), .A4(new_n602), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n536), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n605), .A2(new_n646), .A3(new_n784), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n536), .ZN(new_n866));
  INV_X1    g665(.A(new_n857), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n690), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n849), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n783), .A2(new_n871), .A3(new_n683), .A4(new_n850), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n739), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n866), .B1(new_n873), .B2(new_n860), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n863), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n865), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n482), .A2(new_n477), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n485), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(G113gat), .B1(new_n879), .B2(new_n646), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n646), .A2(G113gat), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT119), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n880), .B1(new_n879), .B2(new_n882), .ZN(G1340gat));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n876), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n477), .A3(new_n482), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n240), .A3(new_n485), .A4(new_n690), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n879), .A2(new_n784), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(G120gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT120), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n886), .B(new_n890), .C1(new_n887), .C2(G120gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1341gat));
  NOR2_X1   g691(.A1(new_n879), .A2(new_n866), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(new_n515), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n700), .A2(new_n602), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n885), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n879), .B2(new_n602), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n898), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(G1343gat));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n865), .A2(new_n876), .A3(new_n903), .A4(new_n375), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT55), .B1(new_n869), .B2(KEYINPUT121), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(KEYINPUT121), .B2(new_n869), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n851), .A2(new_n646), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n858), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n861), .B1(new_n908), .B2(new_n739), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n864), .B1(new_n909), .B2(new_n866), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT57), .B1(new_n910), .B2(new_n374), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n718), .A2(new_n477), .A3(new_n700), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n904), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G141gat), .B1(new_n913), .B2(new_n646), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n884), .A2(new_n374), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n718), .A2(new_n477), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n646), .A2(G141gat), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n915), .A2(new_n485), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n918), .B2(KEYINPUT122), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n919), .B(new_n921), .ZN(G1344gat));
  AND2_X1   g721(.A1(new_n915), .A2(new_n916), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(new_n485), .ZN(new_n924));
  INV_X1    g723(.A(G148gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n690), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(G148gat), .C1(new_n913), .C2(new_n784), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n374), .A2(new_n903), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n865), .A2(new_n876), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n865), .A2(new_n876), .A3(KEYINPUT123), .A4(new_n929), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n903), .B1(new_n910), .B2(new_n374), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n912), .A2(new_n690), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n925), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n928), .B1(new_n937), .B2(new_n927), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n926), .A2(new_n938), .ZN(G1345gat));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n323), .A3(new_n536), .ZN(new_n940));
  OAI21_X1  g739(.A(G155gat), .B1(new_n913), .B2(new_n866), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n324), .A3(new_n896), .ZN(new_n943));
  OAI21_X1  g742(.A(G162gat), .B1(new_n913), .B2(new_n602), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1347gat));
  NOR2_X1   g744(.A1(new_n485), .A2(new_n697), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n797), .A2(new_n375), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n877), .A2(new_n948), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(new_n258), .A3(new_n646), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n884), .A2(new_n697), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n482), .A2(new_n485), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n951), .A2(new_n783), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n950), .B1(new_n954), .B2(new_n258), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n949), .B2(new_n784), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n953), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n690), .A2(new_n259), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(G1349gat));
  NOR2_X1   g758(.A1(new_n949), .A2(new_n866), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n536), .A2(new_n203), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n960), .A2(new_n218), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g762(.A1(new_n739), .A2(new_n204), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n957), .A2(KEYINPUT125), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT125), .B1(new_n957), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n949), .B2(new_n602), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(G1351gat));
  NOR2_X1   g771(.A1(new_n718), .A2(new_n947), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n935), .A2(new_n783), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G197gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n718), .A2(new_n374), .A3(new_n485), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n976), .A2(new_n477), .A3(new_n876), .A4(new_n865), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT126), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n951), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n646), .A2(G197gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT127), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT127), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n975), .B1(new_n983), .B2(new_n984), .ZN(G1352gat));
  NOR2_X1   g784(.A1(new_n784), .A2(G204gat), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT62), .B1(new_n977), .B2(new_n987), .ZN(new_n988));
  OR3_X1    g787(.A1(new_n977), .A2(KEYINPUT62), .A3(new_n987), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n935), .A2(new_n690), .A3(new_n973), .ZN(new_n990));
  INV_X1    g789(.A(G204gat), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n988), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(G1353gat));
  NOR2_X1   g791(.A1(new_n866), .A2(G211gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n980), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n935), .A2(new_n536), .A3(new_n973), .ZN(new_n995));
  AND3_X1   g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  INV_X1    g797(.A(G218gat), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n978), .A2(new_n980), .A3(new_n999), .A4(new_n739), .ZN(new_n1000));
  AND3_X1   g799(.A1(new_n935), .A2(new_n739), .A3(new_n973), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n1001), .B2(new_n999), .ZN(G1355gat));
endmodule


