

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752;

  AND2_X1 U371 ( .A1(n591), .A2(n592), .ZN(n608) );
  NOR2_X1 U372 ( .A1(n707), .A2(n691), .ZN(n526) );
  NAND2_X1 U373 ( .A1(n377), .A2(n577), .ZN(n580) );
  XNOR2_X1 U374 ( .A(n576), .B(n575), .ZN(n377) );
  OR2_X1 U375 ( .A1(n624), .A2(n521), .ZN(n634) );
  NAND2_X1 U376 ( .A1(n350), .A2(n349), .ZN(n576) );
  AND2_X1 U377 ( .A1(n396), .A2(n397), .ZN(n353) );
  INV_X1 U378 ( .A(n581), .ZN(n349) );
  XNOR2_X1 U379 ( .A(n439), .B(n495), .ZN(n737) );
  INV_X1 U380 ( .A(n593), .ZN(n350) );
  NAND2_X1 U381 ( .A1(n570), .A2(n571), .ZN(n593) );
  XNOR2_X2 U382 ( .A(KEYINPUT77), .B(G143), .ZN(n375) );
  NAND2_X1 U383 ( .A1(n351), .A2(n537), .ZN(n539) );
  NOR2_X1 U384 ( .A1(n527), .A2(n688), .ZN(n351) );
  XNOR2_X1 U385 ( .A(n353), .B(n354), .ZN(n649) );
  INV_X1 U386 ( .A(G953), .ZN(n746) );
  INV_X1 U387 ( .A(n492), .ZN(n545) );
  AND2_X1 U388 ( .A1(n390), .A2(n408), .ZN(n391) );
  XNOR2_X2 U389 ( .A(n441), .B(n440), .ZN(n731) );
  XOR2_X2 U390 ( .A(G101), .B(KEYINPUT93), .Z(n441) );
  XNOR2_X2 U391 ( .A(n358), .B(n730), .ZN(n373) );
  XNOR2_X2 U392 ( .A(n509), .B(n409), .ZN(n730) );
  XNOR2_X2 U393 ( .A(n511), .B(n510), .ZN(n669) );
  XNOR2_X2 U394 ( .A(n737), .B(G146), .ZN(n511) );
  INV_X1 U395 ( .A(n397), .ZN(n624) );
  NAND2_X1 U396 ( .A1(n587), .A2(n528), .ZN(n569) );
  AND2_X1 U397 ( .A1(n381), .A2(n389), .ZN(n382) );
  AND2_X1 U398 ( .A1(n376), .A2(n616), .ZN(n742) );
  NAND2_X1 U399 ( .A1(n414), .A2(n412), .ZN(n666) );
  AND2_X1 U400 ( .A1(n417), .A2(n415), .ZN(n414) );
  BUF_X1 U401 ( .A(n519), .Z(n530) );
  XNOR2_X1 U402 ( .A(n577), .B(KEYINPUT106), .ZN(n704) );
  AND2_X1 U403 ( .A1(n561), .A2(n528), .ZN(n396) );
  XNOR2_X1 U404 ( .A(n451), .B(KEYINPUT90), .ZN(n374) );
  NAND2_X2 U405 ( .A1(n382), .A2(n385), .ZN(n584) );
  XNOR2_X1 U406 ( .A(n370), .B(n449), .ZN(n572) );
  XNOR2_X1 U407 ( .A(n375), .B(n438), .ZN(n471) );
  INV_X1 U408 ( .A(n659), .ZN(n660) );
  NOR2_X2 U409 ( .A1(n392), .A2(n391), .ZN(n352) );
  NOR2_X2 U410 ( .A1(n392), .A2(n391), .ZN(n720) );
  XOR2_X1 U411 ( .A(n529), .B(KEYINPUT68), .Z(n354) );
  XNOR2_X1 U412 ( .A(n544), .B(n543), .ZN(n751) );
  NAND2_X1 U413 ( .A1(n545), .A2(n541), .ZN(n544) );
  OR2_X1 U414 ( .A1(n669), .A2(n386), .ZN(n385) );
  XNOR2_X1 U415 ( .A(n374), .B(n421), .ZN(n597) );
  NAND2_X1 U416 ( .A1(n359), .A2(n387), .ZN(n502) );
  INV_X1 U417 ( .A(n683), .ZN(n359) );
  NAND2_X1 U418 ( .A1(n365), .A2(n363), .ZN(n362) );
  AND2_X1 U419 ( .A1(n601), .A2(n600), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n666), .B(n364), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n405), .B(n403), .ZN(n464) );
  XNOR2_X1 U422 ( .A(KEYINPUT82), .B(KEYINPUT8), .ZN(n405) );
  NOR2_X1 U423 ( .A1(n404), .A2(G953), .ZN(n403) );
  INV_X1 U424 ( .A(G234), .ZN(n404) );
  NOR2_X1 U425 ( .A1(G953), .A2(G237), .ZN(n503) );
  XNOR2_X1 U426 ( .A(n731), .B(n442), .ZN(n499) );
  XNOR2_X1 U427 ( .A(n367), .B(G146), .ZN(n445) );
  INV_X1 U428 ( .A(G125), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n610), .B(n609), .ZN(n376) );
  NAND2_X1 U430 ( .A1(n385), .A2(n383), .ZN(n565) );
  INV_X1 U431 ( .A(n523), .ZN(n528) );
  XNOR2_X1 U432 ( .A(G128), .B(G119), .ZN(n425) );
  XOR2_X1 U433 ( .A(KEYINPUT7), .B(KEYINPUT102), .Z(n466) );
  XNOR2_X1 U434 ( .A(KEYINPUT103), .B(KEYINPUT9), .ZN(n465) );
  INV_X1 U435 ( .A(G128), .ZN(n438) );
  XNOR2_X1 U436 ( .A(G116), .B(G122), .ZN(n469) );
  XOR2_X1 U437 ( .A(G134), .B(G107), .Z(n470) );
  XNOR2_X1 U438 ( .A(n445), .B(n366), .ZN(n736) );
  XNOR2_X1 U439 ( .A(G140), .B(KEYINPUT10), .ZN(n366) );
  XNOR2_X1 U440 ( .A(n586), .B(n585), .ZN(n369) );
  NAND2_X1 U441 ( .A1(n572), .A2(n641), .ZN(n451) );
  XNOR2_X1 U442 ( .A(n612), .B(KEYINPUT112), .ZN(n402) );
  NOR2_X1 U443 ( .A1(n573), .A2(KEYINPUT109), .ZN(n416) );
  XNOR2_X1 U444 ( .A(n436), .B(n422), .ZN(n546) );
  OR2_X1 U445 ( .A1(G902), .A2(n661), .ZN(n436) );
  XNOR2_X1 U446 ( .A(n407), .B(n406), .ZN(n532) );
  XNOR2_X1 U447 ( .A(G478), .B(KEYINPUT104), .ZN(n406) );
  NOR2_X1 U448 ( .A1(n722), .A2(G902), .ZN(n407) );
  INV_X1 U449 ( .A(n391), .ZN(n378) );
  INV_X1 U450 ( .A(KEYINPUT81), .ZN(n364) );
  XNOR2_X1 U451 ( .A(n362), .B(KEYINPUT79), .ZN(n361) );
  AND2_X1 U452 ( .A1(n381), .A2(n379), .ZN(n383) );
  NOR2_X1 U453 ( .A1(n384), .A2(n380), .ZN(n379) );
  INV_X1 U454 ( .A(n389), .ZN(n380) );
  INV_X1 U455 ( .A(n641), .ZN(n384) );
  XNOR2_X1 U456 ( .A(KEYINPUT5), .B(G101), .ZN(n504) );
  XNOR2_X1 U457 ( .A(G137), .B(G134), .ZN(n494) );
  XNOR2_X1 U458 ( .A(G131), .B(KEYINPUT66), .ZN(n493) );
  INV_X1 U459 ( .A(KEYINPUT44), .ZN(n549) );
  XOR2_X1 U460 ( .A(KEYINPUT18), .B(KEYINPUT91), .Z(n444) );
  XNOR2_X1 U461 ( .A(n411), .B(n410), .ZN(n509) );
  XNOR2_X1 U462 ( .A(G119), .B(G116), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n437), .B(G113), .ZN(n411) );
  INV_X2 U464 ( .A(KEYINPUT3), .ZN(n437) );
  XNOR2_X1 U465 ( .A(G122), .B(G104), .ZN(n481) );
  NAND2_X1 U466 ( .A1(n669), .A2(n513), .ZN(n381) );
  NAND2_X1 U467 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U468 ( .A(KEYINPUT0), .ZN(n458) );
  AND2_X1 U469 ( .A1(n597), .A2(n457), .ZN(n459) );
  XNOR2_X1 U470 ( .A(G110), .B(G107), .ZN(n440) );
  XNOR2_X1 U471 ( .A(G902), .B(KEYINPUT15), .ZN(n659) );
  XNOR2_X1 U472 ( .A(G143), .B(G131), .ZN(n477) );
  XOR2_X1 U473 ( .A(KEYINPUT100), .B(G113), .Z(n478) );
  XOR2_X1 U474 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n476) );
  XNOR2_X1 U475 ( .A(n471), .B(KEYINPUT4), .ZN(n439) );
  XNOR2_X1 U476 ( .A(n481), .B(KEYINPUT16), .ZN(n409) );
  INV_X1 U477 ( .A(KEYINPUT33), .ZN(n529) );
  XNOR2_X1 U478 ( .A(n398), .B(KEYINPUT85), .ZN(n390) );
  NOR2_X1 U479 ( .A1(n742), .A2(KEYINPUT2), .ZN(n617) );
  NOR2_X1 U480 ( .A1(n643), .A2(n644), .ZN(n582) );
  NAND2_X1 U481 ( .A1(n596), .A2(n597), .ZN(n598) );
  XNOR2_X1 U482 ( .A(n488), .B(n487), .ZN(n533) );
  XNOR2_X1 U483 ( .A(n486), .B(G475), .ZN(n487) );
  XOR2_X1 U484 ( .A(n433), .B(n432), .Z(n661) );
  XNOR2_X1 U485 ( .A(n474), .B(n473), .ZN(n722) );
  AND2_X1 U486 ( .A1(n663), .A2(G953), .ZN(n725) );
  NOR2_X1 U487 ( .A1(n399), .A2(n624), .ZN(n710) );
  XNOR2_X1 U488 ( .A(n401), .B(n400), .ZN(n399) );
  INV_X1 U489 ( .A(KEYINPUT36), .ZN(n400) );
  NAND2_X1 U490 ( .A1(n593), .A2(n413), .ZN(n412) );
  INV_X1 U491 ( .A(KEYINPUT109), .ZN(n413) );
  AND2_X1 U492 ( .A1(n657), .A2(n623), .ZN(n419) );
  INV_X1 U493 ( .A(n368), .ZN(n596) );
  AND2_X1 U494 ( .A1(n573), .A2(KEYINPUT109), .ZN(n355) );
  AND2_X1 U495 ( .A1(n616), .A2(KEYINPUT2), .ZN(n356) );
  INV_X1 U496 ( .A(G902), .ZN(n387) );
  XNOR2_X1 U497 ( .A(n446), .B(n357), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n424), .B(n445), .ZN(n357) );
  XNOR2_X2 U499 ( .A(n584), .B(KEYINPUT6), .ZN(n561) );
  INV_X1 U500 ( .A(n439), .ZN(n358) );
  NAND2_X1 U501 ( .A1(n715), .A2(n659), .ZN(n370) );
  XNOR2_X2 U502 ( .A(n371), .B(n373), .ZN(n715) );
  NAND2_X1 U503 ( .A1(n376), .A2(n356), .ZN(n398) );
  XNOR2_X2 U504 ( .A(n501), .B(n500), .ZN(n683) );
  XNOR2_X1 U505 ( .A(n360), .B(n687), .ZN(G54) );
  NOR2_X2 U506 ( .A1(n686), .A2(n725), .ZN(n360) );
  NAND2_X1 U507 ( .A1(n361), .A2(n605), .ZN(n606) );
  INV_X1 U508 ( .A(n598), .ZN(n702) );
  NAND2_X1 U509 ( .A1(n369), .A2(n587), .ZN(n368) );
  XNOR2_X2 U510 ( .A(n372), .B(n447), .ZN(n371) );
  INV_X1 U511 ( .A(n499), .ZN(n372) );
  NOR2_X1 U512 ( .A1(n402), .A2(n374), .ZN(n401) );
  NAND2_X1 U513 ( .A1(n377), .A2(n706), .ZN(n667) );
  NAND2_X1 U514 ( .A1(n621), .A2(n378), .ZN(n420) );
  INV_X1 U515 ( .A(n513), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n513), .A2(G902), .ZN(n389) );
  NAND2_X1 U517 ( .A1(n393), .A2(n660), .ZN(n392) );
  NAND2_X1 U518 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U519 ( .A(KEYINPUT2), .ZN(n394) );
  NAND2_X1 U520 ( .A1(n408), .A2(n742), .ZN(n395) );
  XNOR2_X2 U521 ( .A(n555), .B(KEYINPUT45), .ZN(n408) );
  XNOR2_X2 U522 ( .A(n587), .B(KEYINPUT1), .ZN(n397) );
  XNOR2_X2 U523 ( .A(n502), .B(G469), .ZN(n587) );
  AND2_X1 U524 ( .A1(n568), .A2(n567), .ZN(n571) );
  XNOR2_X2 U525 ( .A(n580), .B(n579), .ZN(n668) );
  NOR2_X1 U526 ( .A1(n408), .A2(KEYINPUT2), .ZN(n556) );
  NAND2_X1 U527 ( .A1(n408), .A2(n746), .ZN(n729) );
  NOR2_X1 U528 ( .A1(n416), .A2(n595), .ZN(n415) );
  NAND2_X1 U529 ( .A1(n594), .A2(n355), .ZN(n417) );
  XNOR2_X1 U530 ( .A(n418), .B(n658), .ZN(G75) );
  NAND2_X1 U531 ( .A1(n420), .A2(n419), .ZN(n418) );
  INV_X1 U532 ( .A(n546), .ZN(n626) );
  NAND2_X1 U533 ( .A1(n546), .A2(n520), .ZN(n523) );
  XOR2_X1 U534 ( .A(KEYINPUT19), .B(KEYINPUT73), .Z(n421) );
  XOR2_X1 U535 ( .A(n435), .B(KEYINPUT25), .Z(n422) );
  XOR2_X1 U536 ( .A(KEYINPUT86), .B(KEYINPUT46), .Z(n423) );
  AND2_X1 U537 ( .A1(G224), .A2(n746), .ZN(n424) );
  AND2_X1 U538 ( .A1(n558), .A2(n456), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n542), .B(KEYINPUT76), .ZN(n543) );
  XOR2_X1 U540 ( .A(G137), .B(G110), .Z(n426) );
  XNOR2_X1 U541 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U542 ( .A(n736), .B(n427), .ZN(n433) );
  XOR2_X1 U543 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U544 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n428) );
  XNOR2_X1 U545 ( .A(n429), .B(n428), .ZN(n431) );
  NAND2_X1 U546 ( .A1(n464), .A2(G221), .ZN(n430) );
  XOR2_X1 U547 ( .A(n431), .B(n430), .Z(n432) );
  NAND2_X1 U548 ( .A1(G234), .A2(n659), .ZN(n434) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n434), .ZN(n460) );
  NAND2_X1 U550 ( .A1(n460), .A2(G217), .ZN(n435) );
  INV_X1 U551 ( .A(KEYINPUT67), .ZN(n442) );
  XNOR2_X1 U552 ( .A(KEYINPUT74), .B(KEYINPUT17), .ZN(n443) );
  XNOR2_X1 U553 ( .A(n444), .B(n443), .ZN(n446) );
  NOR2_X1 U554 ( .A1(G237), .A2(G902), .ZN(n448) );
  XNOR2_X1 U555 ( .A(KEYINPUT71), .B(n448), .ZN(n450) );
  AND2_X1 U556 ( .A1(n450), .A2(G210), .ZN(n449) );
  NAND2_X1 U557 ( .A1(n450), .A2(G214), .ZN(n641) );
  NAND2_X1 U558 ( .A1(G237), .A2(G234), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n452), .B(KEYINPUT14), .ZN(n653) );
  OR2_X1 U560 ( .A1(n746), .A2(G902), .ZN(n453) );
  NAND2_X1 U561 ( .A1(n653), .A2(n453), .ZN(n455) );
  NOR2_X1 U562 ( .A1(G953), .A2(G952), .ZN(n454) );
  NOR2_X1 U563 ( .A1(n455), .A2(n454), .ZN(n558) );
  NAND2_X1 U564 ( .A1(G953), .A2(G898), .ZN(n456) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n460), .A2(G221), .ZN(n461) );
  XNOR2_X1 U567 ( .A(KEYINPUT21), .B(n461), .ZN(n627) );
  INV_X1 U568 ( .A(KEYINPUT96), .ZN(n462) );
  XNOR2_X1 U569 ( .A(n627), .B(n462), .ZN(n520) );
  INV_X1 U570 ( .A(n520), .ZN(n463) );
  NOR2_X1 U571 ( .A1(n519), .A2(n463), .ZN(n490) );
  NAND2_X1 U572 ( .A1(G217), .A2(n464), .ZN(n468) );
  XNOR2_X1 U573 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U574 ( .A(n468), .B(n467), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n470), .B(n469), .ZN(n472) );
  XOR2_X1 U576 ( .A(n471), .B(n472), .Z(n473) );
  NAND2_X1 U577 ( .A1(n503), .A2(G214), .ZN(n475) );
  XNOR2_X1 U578 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U580 ( .A(n480), .B(n479), .ZN(n484) );
  INV_X1 U581 ( .A(n481), .ZN(n482) );
  XNOR2_X1 U582 ( .A(n482), .B(KEYINPUT11), .ZN(n483) );
  XNOR2_X1 U583 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U584 ( .A(n736), .B(n485), .ZN(n676) );
  NOR2_X1 U585 ( .A1(G902), .A2(n676), .ZN(n488) );
  XNOR2_X1 U586 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n486) );
  NAND2_X1 U587 ( .A1(n532), .A2(n533), .ZN(n643) );
  INV_X1 U588 ( .A(n643), .ZN(n489) );
  NAND2_X1 U589 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U590 ( .A(n491), .B(KEYINPUT22), .ZN(n492) );
  XNOR2_X1 U591 ( .A(n494), .B(n493), .ZN(n495) );
  INV_X1 U592 ( .A(n511), .ZN(n501) );
  XNOR2_X1 U593 ( .A(G140), .B(G104), .ZN(n497) );
  NAND2_X1 U594 ( .A1(n746), .A2(G227), .ZN(n496) );
  XNOR2_X1 U595 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U596 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U597 ( .A1(n503), .A2(G210), .ZN(n505) );
  XNOR2_X1 U598 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U599 ( .A(KEYINPUT72), .B(KEYINPUT97), .ZN(n506) );
  XNOR2_X1 U600 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U601 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U602 ( .A(KEYINPUT98), .ZN(n512) );
  XNOR2_X1 U603 ( .A(n512), .B(G472), .ZN(n513) );
  NOR2_X1 U604 ( .A1(n397), .A2(n561), .ZN(n514) );
  NAND2_X1 U605 ( .A1(n545), .A2(n514), .ZN(n515) );
  NOR2_X1 U606 ( .A1(n626), .A2(n515), .ZN(n688) );
  INV_X1 U607 ( .A(n532), .ZN(n516) );
  NAND2_X1 U608 ( .A1(n516), .A2(n533), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n517), .B(KEYINPUT105), .ZN(n706) );
  INV_X1 U610 ( .A(n533), .ZN(n518) );
  AND2_X1 U611 ( .A1(n518), .A2(n532), .ZN(n577) );
  OR2_X1 U612 ( .A1(n706), .A2(n577), .ZN(n603) );
  INV_X1 U613 ( .A(n603), .ZN(n645) );
  OR2_X1 U614 ( .A1(n584), .A2(n523), .ZN(n521) );
  OR2_X2 U615 ( .A1(n530), .A2(n634), .ZN(n522) );
  XNOR2_X2 U616 ( .A(n522), .B(KEYINPUT31), .ZN(n707) );
  INV_X1 U617 ( .A(n569), .ZN(n524) );
  NAND2_X1 U618 ( .A1(n524), .A2(n584), .ZN(n525) );
  NOR2_X1 U619 ( .A1(n530), .A2(n525), .ZN(n691) );
  NOR2_X1 U620 ( .A1(n645), .A2(n526), .ZN(n527) );
  NOR2_X1 U621 ( .A1(n530), .A2(n649), .ZN(n531) );
  XNOR2_X1 U622 ( .A(n531), .B(KEYINPUT34), .ZN(n535) );
  OR2_X1 U623 ( .A1(n533), .A2(n532), .ZN(n595) );
  XNOR2_X1 U624 ( .A(KEYINPUT75), .B(n595), .ZN(n534) );
  NAND2_X1 U625 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X2 U626 ( .A(n536), .B(KEYINPUT35), .ZN(n750) );
  NAND2_X1 U627 ( .A1(n750), .A2(KEYINPUT44), .ZN(n537) );
  XNOR2_X1 U628 ( .A(n539), .B(KEYINPUT89), .ZN(n554) );
  NAND2_X1 U629 ( .A1(n397), .A2(n626), .ZN(n540) );
  NOR2_X1 U630 ( .A1(n540), .A2(n561), .ZN(n541) );
  XOR2_X1 U631 ( .A(KEYINPUT32), .B(KEYINPUT64), .Z(n542) );
  INV_X1 U632 ( .A(n584), .ZN(n629) );
  NOR2_X1 U633 ( .A1(n629), .A2(n546), .ZN(n547) );
  NAND2_X1 U634 ( .A1(n624), .A2(n547), .ZN(n548) );
  NOR2_X1 U635 ( .A1(n492), .A2(n548), .ZN(n698) );
  NOR2_X2 U636 ( .A1(n751), .A2(n698), .ZN(n550) );
  XNOR2_X1 U637 ( .A(n550), .B(n549), .ZN(n552) );
  NAND2_X1 U638 ( .A1(n550), .A2(n750), .ZN(n551) );
  NAND2_X1 U639 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U640 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U641 ( .A(KEYINPUT83), .B(n556), .ZN(n619) );
  INV_X1 U642 ( .A(n704), .ZN(n560) );
  NAND2_X1 U643 ( .A1(G953), .A2(G900), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n558), .A2(n557), .ZN(n566) );
  NOR2_X1 U645 ( .A1(n627), .A2(n566), .ZN(n559) );
  NAND2_X1 U646 ( .A1(n626), .A2(n559), .ZN(n583) );
  NOR2_X1 U647 ( .A1(n560), .A2(n583), .ZN(n562) );
  NAND2_X1 U648 ( .A1(n562), .A2(n561), .ZN(n612) );
  XNOR2_X1 U649 ( .A(n710), .B(KEYINPUT87), .ZN(n592) );
  INV_X1 U650 ( .A(KEYINPUT108), .ZN(n563) );
  XNOR2_X1 U651 ( .A(n563), .B(KEYINPUT30), .ZN(n564) );
  XNOR2_X1 U652 ( .A(n565), .B(n564), .ZN(n568) );
  INV_X1 U653 ( .A(n566), .ZN(n567) );
  XNOR2_X1 U654 ( .A(n569), .B(KEYINPUT107), .ZN(n570) );
  BUF_X1 U655 ( .A(n572), .Z(n573) );
  XNOR2_X1 U656 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n573), .B(n574), .ZN(n581) );
  XNOR2_X1 U658 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n575) );
  INV_X1 U659 ( .A(KEYINPUT111), .ZN(n578) );
  XNOR2_X1 U660 ( .A(n578), .B(KEYINPUT40), .ZN(n579) );
  INV_X1 U661 ( .A(n581), .ZN(n640) );
  NAND2_X1 U662 ( .A1(n641), .A2(n640), .ZN(n644) );
  XNOR2_X1 U663 ( .A(KEYINPUT41), .B(n582), .ZN(n639) );
  OR2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n586) );
  XOR2_X1 U665 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n585) );
  NOR2_X1 U666 ( .A1(n639), .A2(n368), .ZN(n589) );
  INV_X1 U667 ( .A(KEYINPUT42), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n589), .B(n588), .ZN(n752) );
  NAND2_X1 U669 ( .A1(n668), .A2(n752), .ZN(n590) );
  XNOR2_X1 U670 ( .A(n590), .B(n423), .ZN(n591) );
  INV_X1 U671 ( .A(n593), .ZN(n594) );
  INV_X1 U672 ( .A(n573), .ZN(n614) );
  NAND2_X1 U673 ( .A1(n598), .A2(KEYINPUT47), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n645), .A2(KEYINPUT47), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT80), .B(n599), .ZN(n600) );
  INV_X1 U676 ( .A(KEYINPUT47), .ZN(n602) );
  AND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n702), .A2(n604), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT69), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U681 ( .A(KEYINPUT48), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n624), .A2(n641), .ZN(n611) );
  OR2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U684 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n712) );
  AND2_X1 U686 ( .A1(n667), .A2(n712), .ZN(n616) );
  XOR2_X1 U687 ( .A(n617), .B(KEYINPUT84), .Z(n618) );
  AND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT78), .ZN(n621) );
  NOR2_X1 U690 ( .A1(n639), .A2(n649), .ZN(n622) );
  XOR2_X1 U691 ( .A(KEYINPUT120), .B(n622), .Z(n623) );
  NAND2_X1 U692 ( .A1(n624), .A2(n523), .ZN(n625) );
  XNOR2_X1 U693 ( .A(n625), .B(KEYINPUT50), .ZN(n632) );
  AND2_X1 U694 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U695 ( .A(KEYINPUT49), .B(n628), .Z(n630) );
  NOR2_X1 U696 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U697 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U698 ( .A(n633), .B(KEYINPUT119), .ZN(n636) );
  INV_X1 U699 ( .A(n634), .ZN(n635) );
  NOR2_X1 U700 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U701 ( .A(KEYINPUT51), .B(n637), .Z(n638) );
  NOR2_X1 U702 ( .A1(n639), .A2(n638), .ZN(n651) );
  NOR2_X1 U703 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U704 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U705 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U706 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U707 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U708 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U709 ( .A(KEYINPUT52), .B(n652), .ZN(n655) );
  NAND2_X1 U710 ( .A1(n653), .A2(G952), .ZN(n654) );
  NOR2_X1 U711 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U712 ( .A1(n656), .A2(G953), .ZN(n657) );
  INV_X1 U713 ( .A(KEYINPUT53), .ZN(n658) );
  NAND2_X1 U714 ( .A1(n720), .A2(G217), .ZN(n662) );
  XNOR2_X1 U715 ( .A(n662), .B(n661), .ZN(n664) );
  INV_X1 U716 ( .A(G952), .ZN(n663) );
  NOR2_X2 U717 ( .A1(n664), .A2(n725), .ZN(n665) );
  XNOR2_X1 U718 ( .A(n665), .B(KEYINPUT124), .ZN(G66) );
  XNOR2_X1 U719 ( .A(n666), .B(G143), .ZN(G45) );
  XNOR2_X1 U720 ( .A(n667), .B(G134), .ZN(G36) );
  XNOR2_X1 U721 ( .A(n668), .B(G131), .ZN(G33) );
  AND2_X1 U722 ( .A1(n720), .A2(G472), .ZN(n671) );
  XOR2_X1 U723 ( .A(n669), .B(KEYINPUT62), .Z(n670) );
  XNOR2_X1 U724 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U725 ( .A1(n672), .A2(n725), .ZN(n674) );
  XOR2_X1 U726 ( .A(KEYINPUT92), .B(KEYINPUT63), .Z(n673) );
  XNOR2_X1 U727 ( .A(n674), .B(n673), .ZN(G57) );
  NAND2_X1 U728 ( .A1(n352), .A2(G475), .ZN(n678) );
  XNOR2_X1 U729 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n675) );
  XNOR2_X1 U730 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U731 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U732 ( .A1(n679), .A2(n725), .ZN(n680) );
  XNOR2_X1 U733 ( .A(n680), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U734 ( .A(KEYINPUT123), .ZN(n687) );
  NAND2_X1 U735 ( .A1(n352), .A2(G469), .ZN(n685) );
  XOR2_X1 U736 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n681) );
  XNOR2_X1 U737 ( .A(n681), .B(KEYINPUT58), .ZN(n682) );
  XNOR2_X1 U738 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U739 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U740 ( .A(G101), .B(n688), .Z(G3) );
  XOR2_X1 U741 ( .A(G104), .B(KEYINPUT113), .Z(n690) );
  NAND2_X1 U742 ( .A1(n691), .A2(n704), .ZN(n689) );
  XNOR2_X1 U743 ( .A(n690), .B(n689), .ZN(G6) );
  NAND2_X1 U744 ( .A1(n691), .A2(n706), .ZN(n697) );
  XOR2_X1 U745 ( .A(KEYINPUT116), .B(KEYINPUT27), .Z(n693) );
  XNOR2_X1 U746 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n693), .B(n692), .ZN(n695) );
  XOR2_X1 U748 ( .A(G107), .B(KEYINPUT26), .Z(n694) );
  XNOR2_X1 U749 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U750 ( .A(n697), .B(n696), .ZN(G9) );
  XOR2_X1 U751 ( .A(G110), .B(n698), .Z(G12) );
  XOR2_X1 U752 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n700) );
  NAND2_X1 U753 ( .A1(n702), .A2(n706), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U755 ( .A(G128), .B(n701), .Z(G30) );
  NAND2_X1 U756 ( .A1(n704), .A2(n702), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(G146), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n704), .A2(n707), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n705), .B(G113), .ZN(G15) );
  NAND2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n708), .B(KEYINPUT118), .ZN(n709) );
  XNOR2_X1 U762 ( .A(G116), .B(n709), .ZN(G18) );
  XNOR2_X1 U763 ( .A(G125), .B(n710), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n711), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U765 ( .A(G140), .B(n712), .ZN(G42) );
  AND2_X1 U766 ( .A1(n720), .A2(G210), .ZN(n717) );
  XNOR2_X1 U767 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n713) );
  XOR2_X1 U768 ( .A(n713), .B(KEYINPUT55), .Z(n714) );
  XOR2_X1 U769 ( .A(n715), .B(n714), .Z(n716) );
  XNOR2_X1 U770 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n718), .A2(n725), .ZN(n719) );
  XNOR2_X1 U772 ( .A(n719), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U773 ( .A(n352), .Z(n721) );
  NAND2_X1 U774 ( .A1(n721), .A2(G478), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U776 ( .A1(n725), .A2(n724), .ZN(G63) );
  NAND2_X1 U777 ( .A1(G953), .A2(G224), .ZN(n726) );
  XNOR2_X1 U778 ( .A(KEYINPUT61), .B(n726), .ZN(n727) );
  NAND2_X1 U779 ( .A1(n727), .A2(G898), .ZN(n728) );
  NAND2_X1 U780 ( .A1(n729), .A2(n728), .ZN(n735) );
  XOR2_X1 U781 ( .A(n731), .B(n730), .Z(n733) );
  NOR2_X1 U782 ( .A1(G898), .A2(n746), .ZN(n732) );
  NOR2_X1 U783 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(G69) );
  XNOR2_X1 U785 ( .A(n736), .B(KEYINPUT125), .ZN(n738) );
  XOR2_X1 U786 ( .A(n738), .B(n737), .Z(n743) );
  XNOR2_X1 U787 ( .A(n743), .B(G227), .ZN(n739) );
  NAND2_X1 U788 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U789 ( .A1(G953), .A2(n740), .ZN(n741) );
  XOR2_X1 U790 ( .A(KEYINPUT127), .B(n741), .Z(n749) );
  INV_X1 U791 ( .A(n742), .ZN(n745) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT126), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U796 ( .A(n750), .B(G122), .Z(G24) );
  XOR2_X1 U797 ( .A(G119), .B(n751), .Z(G21) );
  XNOR2_X1 U798 ( .A(G137), .B(n752), .ZN(G39) );
endmodule

