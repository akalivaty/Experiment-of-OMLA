

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT64), .B(n523), .ZN(n660) );
  BUF_X1 U552 ( .A(n614), .Z(n615) );
  OR2_X1 U553 ( .A1(G2105), .A2(n536), .ZN(n537) );
  NOR2_X1 U554 ( .A1(n703), .A2(n702), .ZN(n708) );
  XNOR2_X2 U555 ( .A(n531), .B(KEYINPUT65), .ZN(n532) );
  AND2_X1 U556 ( .A1(n805), .A2(n804), .ZN(n515) );
  OR2_X1 U557 ( .A1(n741), .A2(n740), .ZN(n516) );
  OR2_X1 U558 ( .A1(n706), .A2(n705), .ZN(n709) );
  INV_X1 U559 ( .A(n729), .ZN(n714) );
  XNOR2_X1 U560 ( .A(n736), .B(KEYINPUT32), .ZN(n742) );
  AND2_X1 U561 ( .A1(n742), .A2(n516), .ZN(n764) );
  INV_X1 U562 ( .A(n817), .ZN(n805) );
  XNOR2_X1 U563 ( .A(n591), .B(KEYINPUT15), .ZN(n959) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  XNOR2_X1 U565 ( .A(KEYINPUT85), .B(n542), .ZN(G164) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n654) );
  NAND2_X1 U567 ( .A1(n654), .A2(G89), .ZN(n517) );
  XNOR2_X1 U568 ( .A(n517), .B(KEYINPUT4), .ZN(n519) );
  INV_X1 U569 ( .A(G651), .ZN(n521) );
  NOR2_X1 U570 ( .A1(n634), .A2(n521), .ZN(n655) );
  NAND2_X1 U571 ( .A1(G76), .A2(n655), .ZN(n518) );
  NAND2_X1 U572 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U573 ( .A(n520), .B(KEYINPUT5), .ZN(n529) );
  XNOR2_X1 U574 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n527) );
  NOR2_X1 U575 ( .A1(G543), .A2(n521), .ZN(n522) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n522), .Z(n653) );
  NAND2_X1 U577 ( .A1(G63), .A2(n653), .ZN(n525) );
  NOR2_X1 U578 ( .A1(G651), .A2(n634), .ZN(n523) );
  NAND2_X1 U579 ( .A1(G51), .A2(n660), .ZN(n524) );
  NAND2_X1 U580 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U581 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U583 ( .A(KEYINPUT7), .B(n530), .ZN(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U585 ( .A(G2104), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n536), .A2(G2105), .ZN(n531) );
  NAND2_X1 U587 ( .A1(G126), .A2(n532), .ZN(n535) );
  NOR2_X1 U588 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XOR2_X1 U589 ( .A(KEYINPUT17), .B(n533), .Z(n613) );
  NAND2_X1 U590 ( .A1(G138), .A2(n613), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n541) );
  AND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U593 ( .A1(G114), .A2(n881), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n537), .B(KEYINPUT67), .ZN(n614) );
  NAND2_X1 U595 ( .A1(G102), .A2(n614), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  OR2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U598 ( .A1(G137), .A2(n613), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G113), .A2(n881), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G125), .A2(n532), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n545), .B(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G101), .A2(n614), .ZN(n546) );
  XOR2_X1 U604 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U605 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X2 U606 ( .A1(n550), .A2(n549), .ZN(G160) );
  NAND2_X1 U607 ( .A1(G64), .A2(n653), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G52), .A2(n660), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n559) );
  NAND2_X1 U610 ( .A1(n654), .A2(G90), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U612 ( .A1(G77), .A2(n655), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n556), .ZN(n557) );
  XNOR2_X1 U615 ( .A(KEYINPUT69), .B(n557), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n559), .A2(n558), .ZN(G171) );
  XNOR2_X1 U617 ( .A(G2446), .B(G2443), .ZN(n569) );
  XOR2_X1 U618 ( .A(G2430), .B(KEYINPUT105), .Z(n561) );
  XNOR2_X1 U619 ( .A(G2454), .B(G2435), .ZN(n560) );
  XNOR2_X1 U620 ( .A(n561), .B(n560), .ZN(n565) );
  XOR2_X1 U621 ( .A(G2438), .B(G2427), .Z(n563) );
  XNOR2_X1 U622 ( .A(G1341), .B(G1348), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(n565), .B(n564), .Z(n567) );
  XNOR2_X1 U625 ( .A(KEYINPUT104), .B(G2451), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n569), .B(n568), .ZN(n570) );
  AND2_X1 U628 ( .A1(n570), .A2(G14), .ZN(G401) );
  AND2_X1 U629 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U630 ( .A(G57), .ZN(G237) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n571), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n826) );
  NAND2_X1 U634 ( .A1(n826), .A2(G567), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n572), .Z(G234) );
  NAND2_X1 U636 ( .A1(G56), .A2(n653), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n573), .Z(n580) );
  NAND2_X1 U638 ( .A1(G81), .A2(n654), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT12), .B(n574), .Z(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT71), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G68), .A2(n655), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G43), .A2(n660), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n958) );
  INV_X1 U647 ( .A(G860), .ZN(n603) );
  NOR2_X1 U648 ( .A1(n958), .A2(n603), .ZN(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT72), .B(n583), .Z(G153) );
  XNOR2_X1 U650 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G66), .A2(n653), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G92), .A2(n654), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U655 ( .A1(G54), .A2(n660), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G79), .A2(n655), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT74), .ZN(n589) );
  NOR2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U660 ( .A(G868), .ZN(n672) );
  NAND2_X1 U661 ( .A1(n959), .A2(n672), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U663 ( .A1(G65), .A2(n653), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G78), .A2(n655), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n654), .A2(G91), .ZN(n596) );
  XOR2_X1 U667 ( .A(KEYINPUT70), .B(n596), .Z(n597) );
  NOR2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G53), .A2(n660), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G299) );
  NOR2_X1 U671 ( .A1(G286), .A2(n672), .ZN(n602) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U675 ( .A(n959), .ZN(n895) );
  NAND2_X1 U676 ( .A1(n604), .A2(n895), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n958), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n606), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G868), .A2(n895), .ZN(n607) );
  NOR2_X1 U681 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U683 ( .A1(n532), .A2(G123), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G111), .A2(n881), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n619) );
  BUF_X1 U687 ( .A(n613), .Z(n878) );
  NAND2_X1 U688 ( .A1(G135), .A2(n878), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G99), .A2(n615), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n918) );
  XNOR2_X1 U692 ( .A(G2096), .B(n918), .ZN(n621) );
  INV_X1 U693 ( .A(G2100), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G93), .A2(n654), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G80), .A2(n655), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G55), .A2(n660), .ZN(n624) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(n624), .ZN(n625) );
  NOR2_X1 U700 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n653), .A2(G67), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n673) );
  NAND2_X1 U703 ( .A1(n895), .A2(G559), .ZN(n670) );
  XNOR2_X1 U704 ( .A(n958), .B(n670), .ZN(n629) );
  NOR2_X1 U705 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U706 ( .A(n673), .B(n630), .Z(G145) );
  NAND2_X1 U707 ( .A1(G651), .A2(G74), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G49), .A2(n660), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U710 ( .A1(n653), .A2(n633), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U713 ( .A1(n653), .A2(G62), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(KEYINPUT78), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G50), .A2(n660), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT79), .B(n640), .ZN(n645) );
  NAND2_X1 U718 ( .A1(G88), .A2(n654), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G75), .A2(n655), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U721 ( .A(KEYINPUT80), .B(n643), .Z(n644) );
  NAND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(G303) );
  NAND2_X1 U723 ( .A1(G61), .A2(n653), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G86), .A2(n654), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n655), .A2(G73), .ZN(n648) );
  XOR2_X1 U727 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G48), .A2(n660), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(G305) );
  AND2_X1 U731 ( .A1(n653), .A2(G60), .ZN(n659) );
  NAND2_X1 U732 ( .A1(G85), .A2(n654), .ZN(n657) );
  NAND2_X1 U733 ( .A1(G72), .A2(n655), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n662) );
  NAND2_X1 U736 ( .A1(G47), .A2(n660), .ZN(n661) );
  NAND2_X1 U737 ( .A1(n662), .A2(n661), .ZN(G290) );
  XOR2_X1 U738 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n663) );
  XNOR2_X1 U739 ( .A(n673), .B(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(n664), .B(G288), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n958), .B(G303), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n665), .B(G305), .ZN(n666) );
  XNOR2_X1 U743 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U744 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U745 ( .A(n669), .B(G299), .ZN(n896) );
  XOR2_X1 U746 ( .A(n896), .B(n670), .Z(n671) );
  NAND2_X1 U747 ( .A1(G868), .A2(n671), .ZN(n675) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n677), .ZN(n679) );
  XNOR2_X1 U753 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n678) );
  XNOR2_X1 U754 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U755 ( .A1(G2072), .A2(n680), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U757 ( .A1(G108), .A2(G120), .ZN(n681) );
  NOR2_X1 U758 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U759 ( .A1(G69), .A2(n682), .ZN(n833) );
  NAND2_X1 U760 ( .A1(n833), .A2(G567), .ZN(n689) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n684) );
  NAND2_X1 U762 ( .A1(G132), .A2(G82), .ZN(n683) );
  XNOR2_X1 U763 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U764 ( .A1(n685), .A2(G218), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G96), .A2(n686), .ZN(n832) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n832), .ZN(n687) );
  XNOR2_X1 U767 ( .A(KEYINPUT84), .B(n687), .ZN(n688) );
  NAND2_X1 U768 ( .A1(n689), .A2(n688), .ZN(n834) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n690) );
  NOR2_X1 U770 ( .A1(n834), .A2(n690), .ZN(n831) );
  NAND2_X1 U771 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U772 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U773 ( .A(G1981), .B(KEYINPUT98), .ZN(n691) );
  XNOR2_X1 U774 ( .A(n691), .B(G305), .ZN(n976) );
  NOR2_X1 U775 ( .A1(G1976), .A2(G288), .ZN(n968) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n782) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n781) );
  INV_X1 U778 ( .A(n781), .ZN(n692) );
  NAND2_X2 U779 ( .A1(n782), .A2(n692), .ZN(n729) );
  AND2_X1 U780 ( .A1(n714), .A2(G1996), .ZN(n693) );
  XOR2_X1 U781 ( .A(n693), .B(KEYINPUT26), .Z(n696) );
  AND2_X1 U782 ( .A1(n729), .A2(G1341), .ZN(n694) );
  NOR2_X1 U783 ( .A1(n694), .A2(n958), .ZN(n695) );
  AND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n729), .ZN(n698) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n714), .ZN(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U788 ( .A1(n959), .A2(n701), .ZN(n699) );
  NOR2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n703) );
  AND2_X1 U790 ( .A1(n959), .A2(n701), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n714), .A2(G2072), .ZN(n704) );
  XNOR2_X1 U792 ( .A(n704), .B(KEYINPUT27), .ZN(n706) );
  AND2_X1 U793 ( .A1(G1956), .A2(n729), .ZN(n705) );
  NOR2_X1 U794 ( .A1(G299), .A2(n709), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n712) );
  NAND2_X1 U796 ( .A1(G299), .A2(n709), .ZN(n710) );
  XOR2_X1 U797 ( .A(KEYINPUT28), .B(n710), .Z(n711) );
  NOR2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U799 ( .A(n713), .B(KEYINPUT29), .ZN(n718) );
  XNOR2_X1 U800 ( .A(G1961), .B(KEYINPUT93), .ZN(n984) );
  NAND2_X1 U801 ( .A1(n729), .A2(n984), .ZN(n716) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n945) );
  NAND2_X1 U803 ( .A1(n714), .A2(n945), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n722) );
  NAND2_X1 U805 ( .A1(G171), .A2(n722), .ZN(n717) );
  NAND2_X1 U806 ( .A1(n718), .A2(n717), .ZN(n727) );
  NAND2_X1 U807 ( .A1(G8), .A2(n729), .ZN(n748) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n748), .ZN(n741) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n729), .ZN(n737) );
  NOR2_X1 U810 ( .A1(n741), .A2(n737), .ZN(n719) );
  NAND2_X1 U811 ( .A1(G8), .A2(n719), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(G168), .A2(n721), .ZN(n724) );
  NOR2_X1 U814 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U816 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U818 ( .A1(n739), .A2(G286), .ZN(n728) );
  XNOR2_X1 U819 ( .A(n728), .B(KEYINPUT94), .ZN(n734) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n748), .ZN(n731) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n729), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n732), .A2(G303), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U825 ( .A1(n735), .A2(G8), .ZN(n736) );
  NAND2_X1 U826 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n968), .A2(n764), .ZN(n747) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n743) );
  XNOR2_X1 U830 ( .A(n743), .B(KEYINPUT95), .ZN(n745) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n744) );
  AND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n751) );
  NAND2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n966) );
  INV_X1 U835 ( .A(n748), .ZN(n765) );
  AND2_X1 U836 ( .A1(n966), .A2(n765), .ZN(n749) );
  OR2_X1 U837 ( .A1(KEYINPUT33), .A2(n749), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT96), .ZN(n753) );
  NOR2_X1 U840 ( .A1(n976), .A2(n753), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n968), .A2(KEYINPUT33), .ZN(n754) );
  XNOR2_X1 U842 ( .A(KEYINPUT97), .B(n754), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n755), .A2(n765), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n761) );
  NOR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n758) );
  XNOR2_X1 U846 ( .A(n758), .B(KEYINPUT24), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n759), .A2(n765), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n768) );
  NAND2_X1 U849 ( .A1(G166), .A2(G8), .ZN(n762) );
  NOR2_X1 U850 ( .A1(G2090), .A2(n762), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  INV_X1 U854 ( .A(n769), .ZN(n806) );
  NAND2_X1 U855 ( .A1(n615), .A2(G104), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT86), .ZN(n772) );
  NAND2_X1 U857 ( .A1(G140), .A2(n878), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n773), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n881), .A2(G116), .ZN(n774) );
  XOR2_X1 U861 ( .A(KEYINPUT87), .B(n774), .Z(n776) );
  NAND2_X1 U862 ( .A1(n532), .A2(G128), .ZN(n775) );
  NAND2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U866 ( .A(KEYINPUT36), .B(n780), .ZN(n891) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U868 ( .A1(n891), .A2(n819), .ZN(n915) );
  NOR2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n821) );
  NAND2_X1 U870 ( .A1(n915), .A2(n821), .ZN(n783) );
  XOR2_X1 U871 ( .A(KEYINPUT88), .B(n783), .Z(n817) );
  NAND2_X1 U872 ( .A1(G129), .A2(n532), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G117), .A2(n881), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U875 ( .A(KEYINPUT90), .B(n786), .ZN(n790) );
  NAND2_X1 U876 ( .A1(G105), .A2(n615), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(KEYINPUT91), .ZN(n788) );
  XNOR2_X1 U878 ( .A(n788), .B(KEYINPUT38), .ZN(n789) );
  NOR2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n878), .A2(G141), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n871) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n871), .ZN(n793) );
  XOR2_X1 U883 ( .A(KEYINPUT92), .B(n793), .Z(n802) );
  NAND2_X1 U884 ( .A1(G131), .A2(n878), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G95), .A2(n615), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G119), .A2(n532), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G107), .A2(n881), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT89), .B(n798), .Z(n799) );
  NOR2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n870) );
  INV_X1 U892 ( .A(G1991), .ZN(n939) );
  NOR2_X1 U893 ( .A1(n870), .A2(n939), .ZN(n801) );
  NOR2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n910) );
  XOR2_X1 U895 ( .A(G1986), .B(G290), .Z(n970) );
  NAND2_X1 U896 ( .A1(n910), .A2(n970), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n803), .A2(n821), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n806), .A2(n515), .ZN(n824) );
  XNOR2_X1 U899 ( .A(KEYINPUT39), .B(KEYINPUT102), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT101), .ZN(n815) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n871), .ZN(n926) );
  INV_X1 U902 ( .A(n910), .ZN(n812) );
  AND2_X1 U903 ( .A1(n939), .A2(n870), .ZN(n808) );
  XOR2_X1 U904 ( .A(KEYINPUT99), .B(n808), .Z(n919) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n919), .A2(n809), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT100), .ZN(n811) );
  NOR2_X1 U908 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n926), .A2(n813), .ZN(n814) );
  XNOR2_X1 U910 ( .A(n815), .B(n814), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT103), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n891), .A2(n819), .ZN(n917) );
  NAND2_X1 U914 ( .A1(n820), .A2(n917), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT106), .B(n827), .Z(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  XOR2_X1 U923 ( .A(KEYINPUT107), .B(n829), .Z(n830) );
  NAND2_X1 U924 ( .A1(n831), .A2(n830), .ZN(G188) );
  XOR2_X1 U925 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  NOR2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G325) );
  XNOR2_X1 U927 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G108), .ZN(G238) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G82), .ZN(G220) );
  INV_X1 U933 ( .A(n834), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2096), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2072), .B(KEYINPUT42), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n837), .B(G2678), .Z(n839) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U940 ( .A(KEYINPUT110), .B(G2100), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U944 ( .A(G1981), .B(G1956), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1961), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U947 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U950 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U951 ( .A(G2474), .B(KEYINPUT111), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U953 ( .A(G1966), .B(KEYINPUT41), .Z(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U955 ( .A1(n532), .A2(G124), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U957 ( .A1(G136), .A2(n878), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(KEYINPUT112), .B(n857), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G112), .A2(n881), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G100), .A2(n615), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U963 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G130), .A2(n532), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G118), .A2(n881), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n615), .A2(G106), .ZN(n864) );
  XOR2_X1 U968 ( .A(KEYINPUT113), .B(n864), .Z(n866) );
  NAND2_X1 U969 ( .A1(n878), .A2(G142), .ZN(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n867), .Z(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n890) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(n873) );
  XNOR2_X1 U974 ( .A(G164), .B(G160), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n873), .B(n872), .ZN(n877) );
  XOR2_X1 U976 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n875) );
  XNOR2_X1 U977 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(n877), .B(n876), .Z(n888) );
  NAND2_X1 U980 ( .A1(G139), .A2(n878), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G103), .A2(n615), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G127), .A2(n532), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G115), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n906) );
  XNOR2_X1 U988 ( .A(n918), .B(n906), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n891), .B(G162), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U993 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n895), .B(G286), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n898), .B(G171), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G37), .A2(n899), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n900), .Z(n901) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n901), .ZN(n902) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n902), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(n903), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  INV_X1 U1007 ( .A(KEYINPUT55), .ZN(n954) );
  XOR2_X1 U1008 ( .A(G2072), .B(n906), .Z(n908) );
  XOR2_X1 U1009 ( .A(G164), .B(G2078), .Z(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(KEYINPUT50), .B(n909), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G2084), .B(G160), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(KEYINPUT117), .B(n912), .ZN(n913) );
  NOR2_X1 U1015 ( .A1(n914), .A2(n913), .ZN(n924) );
  INV_X1 U1016 ( .A(n915), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1019 ( .A(KEYINPUT118), .B(n920), .Z(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n927), .Z(n929) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n929), .B(n928), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n932), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n954), .A2(n933), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1031 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(G34), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(G2084), .B(n936), .ZN(n952) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G35), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G25), .B(n939), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n940), .A2(G28), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G26), .B(G2067), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1043 ( .A(G27), .B(n945), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n954), .B(n953), .ZN(n956) );
  INV_X1 U1049 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n957), .ZN(n1013) );
  XNOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .ZN(n983) );
  XNOR2_X1 U1053 ( .A(n958), .B(G1341), .ZN(n964) );
  XOR2_X1 U1054 ( .A(G171), .B(G1961), .Z(n961) );
  XNOR2_X1 U1055 ( .A(n959), .B(G1348), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT123), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n981) );
  XOR2_X1 U1059 ( .A(G1956), .B(G299), .Z(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G1971), .B(G166), .Z(n971) );
  NOR2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1065 ( .A(KEYINPUT124), .B(n973), .Z(n979) );
  XOR2_X1 U1066 ( .A(G1966), .B(G168), .Z(n974) );
  XNOR2_X1 U1067 ( .A(KEYINPUT122), .B(n974), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(KEYINPUT57), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n1011) );
  INV_X1 U1073 ( .A(G16), .ZN(n1009) );
  XNOR2_X1 U1074 ( .A(G5), .B(n984), .ZN(n999) );
  XOR2_X1 U1075 ( .A(KEYINPUT126), .B(G4), .Z(n986) );
  XNOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(n989) );
  XOR2_X1 U1078 ( .A(KEYINPUT125), .B(G1981), .Z(n987) );
  XNOR2_X1 U1079 ( .A(G6), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(G1956), .B(G20), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(KEYINPUT60), .ZN(n997) );
  XOR2_X1 U1086 ( .A(KEYINPUT127), .B(G1966), .Z(n995) );
  XNOR2_X1 U1087 ( .A(G21), .B(n995), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1003) );
  XOR2_X1 U1093 ( .A(G1986), .B(G24), .Z(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT61), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1016), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

