

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U553 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X2 U554 ( .A1(n664), .A2(n598), .ZN(n600) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n647) );
  NOR2_X1 U556 ( .A1(n655), .A2(n654), .ZN(n657) );
  INV_X1 U557 ( .A(KEYINPUT98), .ZN(n621) );
  XNOR2_X1 U558 ( .A(n631), .B(KEYINPUT27), .ZN(n633) );
  XNOR2_X1 U559 ( .A(n660), .B(KEYINPUT102), .ZN(n677) );
  AND2_X1 U560 ( .A1(n701), .A2(n700), .ZN(n702) );
  INV_X1 U561 ( .A(G2104), .ZN(n524) );
  XOR2_X1 U562 ( .A(KEYINPUT96), .B(n632), .Z(n517) );
  AND2_X1 U563 ( .A1(G8), .A2(n674), .ZN(n518) );
  NOR2_X1 U564 ( .A1(n674), .A2(n650), .ZN(n651) );
  XNOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n656) );
  XNOR2_X1 U566 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X1 U567 ( .A1(n675), .A2(n518), .ZN(n676) );
  AND2_X1 U568 ( .A1(n677), .A2(n676), .ZN(n678) );
  INV_X1 U569 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U570 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U571 ( .A1(G651), .A2(n561), .ZN(n799) );
  NOR2_X1 U572 ( .A1(n561), .A2(n533), .ZN(n795) );
  NOR2_X1 U573 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U574 ( .A(G2105), .ZN(n522) );
  AND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n885) );
  NAND2_X1 U576 ( .A1(n885), .A2(G113), .ZN(n521) );
  AND2_X4 U577 ( .A1(n522), .A2(G2104), .ZN(n880) );
  NAND2_X1 U578 ( .A1(G101), .A2(n880), .ZN(n519) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n519), .Z(n520) );
  NAND2_X1 U580 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X2 U581 ( .A1(G2104), .A2(n522), .ZN(n884) );
  NAND2_X1 U582 ( .A1(G125), .A2(n884), .ZN(n527) );
  XNOR2_X2 U583 ( .A(n525), .B(KEYINPUT17), .ZN(n881) );
  NAND2_X1 U584 ( .A1(G137), .A2(n881), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U586 ( .A1(n533), .A2(G543), .ZN(n530) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n530), .Z(n604) );
  BUF_X1 U588 ( .A(n604), .Z(n802) );
  NAND2_X1 U589 ( .A1(G64), .A2(n802), .ZN(n532) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n561) );
  NAND2_X1 U591 ( .A1(G52), .A2(n799), .ZN(n531) );
  AND2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT64), .B(KEYINPUT9), .ZN(n537) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n794) );
  NAND2_X1 U595 ( .A1(G90), .A2(n794), .ZN(n535) );
  INV_X1 U596 ( .A(G651), .ZN(n533) );
  NAND2_X1 U597 ( .A1(G77), .A2(n795), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U600 ( .A1(n539), .A2(n538), .ZN(G301) );
  NAND2_X1 U601 ( .A1(n794), .A2(G89), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  NAND2_X1 U603 ( .A1(G76), .A2(n795), .ZN(n541) );
  NAND2_X1 U604 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT5), .ZN(n549) );
  XNOR2_X1 U606 ( .A(KEYINPUT6), .B(KEYINPUT69), .ZN(n547) );
  NAND2_X1 U607 ( .A1(G63), .A2(n802), .ZN(n545) );
  NAND2_X1 U608 ( .A1(G51), .A2(n799), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(KEYINPUT7), .B(n550), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G88), .A2(n794), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G75), .A2(n795), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G62), .A2(n802), .ZN(n554) );
  NAND2_X1 U618 ( .A1(G50), .A2(n799), .ZN(n553) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(KEYINPUT77), .B(n555), .Z(n556) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(G166) );
  XNOR2_X1 U622 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U623 ( .A1(G49), .A2(n799), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G74), .A2(G651), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U626 ( .A1(n802), .A2(n560), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(G87), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(G288) );
  NAND2_X1 U629 ( .A1(G73), .A2(n795), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT2), .ZN(n571) );
  NAND2_X1 U631 ( .A1(G61), .A2(n802), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G86), .A2(n794), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G48), .A2(n799), .ZN(n567) );
  XNOR2_X1 U635 ( .A(KEYINPUT75), .B(n567), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT76), .B(n572), .ZN(G305) );
  NAND2_X1 U639 ( .A1(G85), .A2(n794), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G72), .A2(n795), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G60), .A2(n802), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G47), .A2(n799), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  OR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(G290) );
  NAND2_X1 U646 ( .A1(G56), .A2(n604), .ZN(n579) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n579), .Z(n585) );
  NAND2_X1 U648 ( .A1(n794), .A2(G81), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT12), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G68), .A2(n795), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(n583), .Z(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n799), .A2(G43), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n924) );
  NAND2_X1 U656 ( .A1(G138), .A2(n881), .ZN(n589) );
  INV_X1 U657 ( .A(KEYINPUT88), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n589), .B(n588), .ZN(n596) );
  NAND2_X1 U659 ( .A1(G114), .A2(n885), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT87), .B(n590), .Z(n594) );
  NAND2_X1 U661 ( .A1(G126), .A2(n884), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G102), .A2(n880), .ZN(n591) );
  AND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(G164) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NAND2_X1 U667 ( .A1(G160), .A2(G40), .ZN(n710) );
  INV_X1 U668 ( .A(n710), .ZN(n597) );
  NAND2_X2 U669 ( .A1(n711), .A2(n597), .ZN(n664) );
  INV_X1 U670 ( .A(G1996), .ZN(n598) );
  INV_X1 U671 ( .A(KEYINPUT26), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n600), .B(n599), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n664), .A2(G1341), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U675 ( .A1(n924), .A2(n603), .ZN(n620) );
  INV_X1 U676 ( .A(KEYINPUT67), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n604), .A2(G66), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n606), .B(n605), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n794), .A2(G92), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U681 ( .A(KEYINPUT68), .B(n609), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G79), .A2(n795), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G54), .A2(n799), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  XOR2_X1 U686 ( .A(KEYINPUT15), .B(n614), .Z(n927) );
  NAND2_X1 U687 ( .A1(n620), .A2(n927), .ZN(n619) );
  NAND2_X1 U688 ( .A1(G1348), .A2(n664), .ZN(n616) );
  INV_X1 U689 ( .A(n664), .ZN(n642) );
  NAND2_X1 U690 ( .A1(G2067), .A2(n642), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT97), .B(n617), .Z(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n620), .A2(n927), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n635) );
  NAND2_X1 U697 ( .A1(G65), .A2(n802), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G53), .A2(n799), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G91), .A2(n794), .ZN(n628) );
  NAND2_X1 U701 ( .A1(G78), .A2(n795), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n928) );
  NAND2_X1 U704 ( .A1(n642), .A2(G2072), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G1956), .A2(n664), .ZN(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n517), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n928), .A2(n636), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n639) );
  NOR2_X1 U709 ( .A1(n928), .A2(n636), .ZN(n637) );
  XOR2_X1 U710 ( .A(n637), .B(KEYINPUT28), .Z(n638) );
  NAND2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n641) );
  XOR2_X1 U712 ( .A(KEYINPUT99), .B(KEYINPUT29), .Z(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n646) );
  NAND2_X1 U714 ( .A1(G1961), .A2(n664), .ZN(n644) );
  XOR2_X1 U715 ( .A(G2078), .B(KEYINPUT25), .Z(n974) );
  NAND2_X1 U716 ( .A1(n642), .A2(n974), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n653), .A2(G301), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n648) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(n659) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n664), .ZN(n674) );
  NAND2_X1 U722 ( .A1(G8), .A2(n664), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n662), .A2(G1966), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(KEYINPUT95), .ZN(n673) );
  NAND2_X1 U725 ( .A1(G8), .A2(n673), .ZN(n650) );
  XOR2_X1 U726 ( .A(KEYINPUT30), .B(n651), .Z(n652) );
  NOR2_X1 U727 ( .A1(G168), .A2(n652), .ZN(n655) );
  AND2_X1 U728 ( .A1(G301), .A2(n653), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  AND2_X1 U730 ( .A1(G286), .A2(G8), .ZN(n661) );
  NAND2_X1 U731 ( .A1(n677), .A2(n661), .ZN(n671) );
  INV_X1 U732 ( .A(G8), .ZN(n669) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n662), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(KEYINPUT104), .ZN(n666) );
  NOR2_X1 U735 ( .A1(n664), .A2(G2090), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n667), .A2(G303), .ZN(n668) );
  OR2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  AND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U740 ( .A(KEYINPUT32), .B(n672), .ZN(n680) );
  INV_X1 U741 ( .A(n673), .ZN(n675) );
  XNOR2_X1 U742 ( .A(KEYINPUT103), .B(n678), .ZN(n679) );
  NAND2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n697) );
  NOR2_X1 U744 ( .A1(G1976), .A2(G288), .ZN(n681) );
  XOR2_X1 U745 ( .A(KEYINPUT105), .B(n681), .Z(n684) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n684), .A2(n682), .ZN(n934) );
  NAND2_X1 U748 ( .A1(n697), .A2(n934), .ZN(n683) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n929) );
  NAND2_X1 U750 ( .A1(n683), .A2(n929), .ZN(n692) );
  NAND2_X1 U751 ( .A1(KEYINPUT33), .A2(n684), .ZN(n685) );
  XNOR2_X1 U752 ( .A(KEYINPUT106), .B(n685), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n662), .A2(n686), .ZN(n689) );
  XNOR2_X1 U754 ( .A(KEYINPUT107), .B(G1981), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(G305), .ZN(n920) );
  INV_X1 U756 ( .A(n920), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n694) );
  INV_X1 U758 ( .A(n694), .ZN(n690) );
  OR2_X1 U759 ( .A1(n662), .A2(n690), .ZN(n691) );
  NOR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n703) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U762 ( .A1(G8), .A2(n693), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n694), .A2(KEYINPUT33), .ZN(n698) );
  AND2_X1 U764 ( .A1(n695), .A2(n698), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n701) );
  INV_X1 U766 ( .A(n698), .ZN(n699) );
  OR2_X1 U767 ( .A1(n699), .A2(n662), .ZN(n700) );
  XNOR2_X1 U768 ( .A(n704), .B(KEYINPUT108), .ZN(n709) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XOR2_X1 U770 ( .A(n705), .B(KEYINPUT24), .Z(n706) );
  NOR2_X1 U771 ( .A1(n662), .A2(n706), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT94), .ZN(n708) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n743) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n755) );
  XNOR2_X1 U775 ( .A(KEYINPUT37), .B(G2067), .ZN(n746) );
  NAND2_X1 U776 ( .A1(n880), .A2(G104), .ZN(n712) );
  XNOR2_X1 U777 ( .A(n712), .B(KEYINPUT90), .ZN(n714) );
  NAND2_X1 U778 ( .A1(G140), .A2(n881), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U780 ( .A(KEYINPUT34), .B(n715), .ZN(n720) );
  NAND2_X1 U781 ( .A1(G128), .A2(n884), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G116), .A2(n885), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U784 ( .A(KEYINPUT35), .B(n718), .Z(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(KEYINPUT36), .B(n721), .ZN(n867) );
  NOR2_X1 U787 ( .A1(n746), .A2(n867), .ZN(n1007) );
  NAND2_X1 U788 ( .A1(n755), .A2(n1007), .ZN(n752) );
  XOR2_X1 U789 ( .A(KEYINPUT92), .B(KEYINPUT38), .Z(n723) );
  NAND2_X1 U790 ( .A1(G105), .A2(n880), .ZN(n722) );
  XNOR2_X1 U791 ( .A(n723), .B(n722), .ZN(n727) );
  NAND2_X1 U792 ( .A1(G117), .A2(n885), .ZN(n725) );
  NAND2_X1 U793 ( .A1(G141), .A2(n881), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U795 ( .A1(n727), .A2(n726), .ZN(n729) );
  NAND2_X1 U796 ( .A1(n884), .A2(G129), .ZN(n728) );
  NAND2_X1 U797 ( .A1(n729), .A2(n728), .ZN(n893) );
  NAND2_X1 U798 ( .A1(G1996), .A2(n893), .ZN(n730) );
  XNOR2_X1 U799 ( .A(n730), .B(KEYINPUT93), .ZN(n739) );
  NAND2_X1 U800 ( .A1(G119), .A2(n884), .ZN(n732) );
  NAND2_X1 U801 ( .A1(G131), .A2(n881), .ZN(n731) );
  NAND2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n736) );
  NAND2_X1 U803 ( .A1(G95), .A2(n880), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G107), .A2(n885), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U807 ( .A(n737), .B(KEYINPUT91), .ZN(n868) );
  AND2_X1 U808 ( .A1(G1991), .A2(n868), .ZN(n738) );
  NOR2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n1015) );
  INV_X1 U810 ( .A(n755), .ZN(n740) );
  NOR2_X1 U811 ( .A1(n1015), .A2(n740), .ZN(n749) );
  INV_X1 U812 ( .A(n749), .ZN(n741) );
  NAND2_X1 U813 ( .A1(n752), .A2(n741), .ZN(n742) );
  NOR2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n936) );
  NAND2_X1 U816 ( .A1(n936), .A2(n755), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n745), .A2(n744), .ZN(n758) );
  NAND2_X1 U818 ( .A1(n746), .A2(n867), .ZN(n1014) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n893), .ZN(n1010) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n868), .ZN(n1001) );
  NOR2_X1 U821 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U822 ( .A1(n1001), .A2(n747), .ZN(n748) );
  NOR2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U824 ( .A1(n1010), .A2(n750), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(KEYINPUT39), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n1014), .A2(n754), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U831 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U832 ( .A(KEYINPUT66), .B(G132), .Z(G219) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U834 ( .A(KEYINPUT65), .B(G57), .ZN(G237) );
  NOR2_X1 U835 ( .A1(G219), .A2(G220), .ZN(n761) );
  XNOR2_X1 U836 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n760) );
  XNOR2_X1 U837 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U838 ( .A(KEYINPUT22), .B(n762), .ZN(n763) );
  NOR2_X1 U839 ( .A1(G218), .A2(n763), .ZN(n764) );
  NAND2_X1 U840 ( .A1(G96), .A2(n764), .ZN(n917) );
  NAND2_X1 U841 ( .A1(n917), .A2(G2106), .ZN(n769) );
  NAND2_X1 U842 ( .A1(G69), .A2(G120), .ZN(n765) );
  NOR2_X1 U843 ( .A1(G237), .A2(n765), .ZN(n766) );
  XNOR2_X1 U844 ( .A(KEYINPUT84), .B(n766), .ZN(n767) );
  NAND2_X1 U845 ( .A1(n767), .A2(G108), .ZN(n918) );
  NAND2_X1 U846 ( .A1(n918), .A2(G567), .ZN(n768) );
  AND2_X1 U847 ( .A1(n769), .A2(n768), .ZN(G319) );
  AND2_X1 U848 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U849 ( .A1(G7), .A2(G661), .ZN(n771) );
  XNOR2_X1 U850 ( .A(n771), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U851 ( .A(G223), .ZN(n832) );
  NAND2_X1 U852 ( .A1(n832), .A2(G567), .ZN(n772) );
  XOR2_X1 U853 ( .A(KEYINPUT11), .B(n772), .Z(G234) );
  INV_X1 U854 ( .A(G860), .ZN(n777) );
  OR2_X1 U855 ( .A1(n924), .A2(n777), .ZN(G153) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n774) );
  OR2_X1 U857 ( .A1(n927), .A2(G868), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n774), .A2(n773), .ZN(G284) );
  INV_X1 U859 ( .A(n928), .ZN(G299) );
  INV_X1 U860 ( .A(G868), .ZN(n820) );
  NOR2_X1 U861 ( .A1(G286), .A2(n820), .ZN(n776) );
  NOR2_X1 U862 ( .A1(G868), .A2(G299), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(G297) );
  NAND2_X1 U864 ( .A1(G559), .A2(n777), .ZN(n778) );
  XNOR2_X1 U865 ( .A(KEYINPUT70), .B(n778), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n779), .A2(n927), .ZN(n780) );
  XNOR2_X1 U867 ( .A(KEYINPUT16), .B(n780), .ZN(G148) );
  NOR2_X1 U868 ( .A1(G868), .A2(n924), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n927), .A2(G868), .ZN(n781) );
  NOR2_X1 U870 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U872 ( .A1(G99), .A2(n880), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G111), .A2(n885), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n786), .B(KEYINPUT71), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G135), .A2(n881), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U878 ( .A1(n884), .A2(G123), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT18), .B(n789), .Z(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n1000) );
  XNOR2_X1 U881 ( .A(n1000), .B(G2096), .ZN(n793) );
  INV_X1 U882 ( .A(G2100), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(G156) );
  NAND2_X1 U884 ( .A1(G93), .A2(n794), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G80), .A2(n795), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(KEYINPUT73), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G55), .A2(n799), .ZN(n800) );
  NAND2_X1 U889 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n802), .A2(G67), .ZN(n803) );
  XOR2_X1 U891 ( .A(KEYINPUT74), .B(n803), .Z(n804) );
  OR2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n819) );
  XNOR2_X1 U893 ( .A(KEYINPUT72), .B(n924), .ZN(n806) );
  NAND2_X1 U894 ( .A1(n927), .A2(G559), .ZN(n816) );
  XNOR2_X1 U895 ( .A(n806), .B(n816), .ZN(n807) );
  NOR2_X1 U896 ( .A1(G860), .A2(n807), .ZN(n808) );
  XOR2_X1 U897 ( .A(n819), .B(n808), .Z(G145) );
  XNOR2_X1 U898 ( .A(KEYINPUT19), .B(KEYINPUT78), .ZN(n810) );
  XNOR2_X1 U899 ( .A(G288), .B(n928), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n810), .B(n809), .ZN(n813) );
  XNOR2_X1 U901 ( .A(G166), .B(n819), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n924), .B(n811), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n813), .B(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(n814), .B(G290), .ZN(n815) );
  XNOR2_X1 U905 ( .A(G305), .B(n815), .ZN(n855) );
  XNOR2_X1 U906 ( .A(KEYINPUT79), .B(n816), .ZN(n817) );
  XNOR2_X1 U907 ( .A(n855), .B(n817), .ZN(n818) );
  NAND2_X1 U908 ( .A1(n818), .A2(G868), .ZN(n822) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n822), .A2(n821), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2084), .A2(G2078), .ZN(n824) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n823) );
  XNOR2_X1 U913 ( .A(n824), .B(n823), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n825), .A2(G2090), .ZN(n826) );
  XOR2_X1 U915 ( .A(KEYINPUT21), .B(n826), .Z(n827) );
  XNOR2_X1 U916 ( .A(KEYINPUT81), .B(n827), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(G2072), .ZN(G158) );
  NAND2_X1 U918 ( .A1(G661), .A2(G483), .ZN(n829) );
  XNOR2_X1 U919 ( .A(KEYINPUT85), .B(n829), .ZN(n830) );
  NAND2_X1 U920 ( .A1(n830), .A2(G319), .ZN(n831) );
  XOR2_X1 U921 ( .A(KEYINPUT86), .B(n831), .Z(n835) );
  NAND2_X1 U922 ( .A1(G36), .A2(n835), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U925 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n835), .A2(n834), .ZN(G188) );
  XOR2_X1 U928 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U929 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U931 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n842) );
  XNOR2_X1 U936 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U937 ( .A(KEYINPUT111), .B(G1956), .Z(n845) );
  XNOR2_X1 U938 ( .A(G1971), .B(G1961), .ZN(n844) );
  XNOR2_X1 U939 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U940 ( .A(n846), .B(G2474), .Z(n848) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U943 ( .A(G1966), .B(G1976), .Z(n850) );
  XNOR2_X1 U944 ( .A(G1986), .B(G1981), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U946 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U947 ( .A(KEYINPUT41), .B(KEYINPUT112), .ZN(n853) );
  XNOR2_X1 U948 ( .A(n854), .B(n853), .ZN(G229) );
  XNOR2_X1 U949 ( .A(n927), .B(G286), .ZN(n856) );
  XNOR2_X1 U950 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U951 ( .A(G301), .B(n857), .Z(n858) );
  NOR2_X1 U952 ( .A1(G37), .A2(n858), .ZN(n859) );
  XOR2_X1 U953 ( .A(KEYINPUT115), .B(n859), .Z(G397) );
  NAND2_X1 U954 ( .A1(n884), .A2(G124), .ZN(n860) );
  XNOR2_X1 U955 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U956 ( .A1(G112), .A2(n885), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U958 ( .A1(G100), .A2(n880), .ZN(n864) );
  NAND2_X1 U959 ( .A1(G136), .A2(n881), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U961 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U962 ( .A(G164), .B(n867), .ZN(n869) );
  XNOR2_X1 U963 ( .A(n869), .B(n868), .ZN(n879) );
  NAND2_X1 U964 ( .A1(G130), .A2(n884), .ZN(n871) );
  NAND2_X1 U965 ( .A1(G118), .A2(n885), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U967 ( .A1(n880), .A2(G106), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT113), .B(n872), .Z(n874) );
  NAND2_X1 U969 ( .A1(n881), .A2(G142), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U971 ( .A(KEYINPUT45), .B(n875), .Z(n876) );
  NOR2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U973 ( .A(n879), .B(n878), .Z(n892) );
  NAND2_X1 U974 ( .A1(G103), .A2(n880), .ZN(n883) );
  NAND2_X1 U975 ( .A1(G139), .A2(n881), .ZN(n882) );
  NAND2_X1 U976 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U977 ( .A1(G127), .A2(n884), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G115), .A2(n885), .ZN(n886) );
  NAND2_X1 U979 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U981 ( .A1(n890), .A2(n889), .ZN(n995) );
  XNOR2_X1 U982 ( .A(n995), .B(n1000), .ZN(n891) );
  XNOR2_X1 U983 ( .A(n892), .B(n891), .ZN(n898) );
  XNOR2_X1 U984 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n895) );
  XNOR2_X1 U985 ( .A(n893), .B(G162), .ZN(n894) );
  XNOR2_X1 U986 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U987 ( .A(G160), .B(n896), .Z(n897) );
  XNOR2_X1 U988 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U989 ( .A1(G37), .A2(n899), .ZN(n900) );
  XNOR2_X1 U990 ( .A(KEYINPUT114), .B(n900), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G2451), .B(G2443), .ZN(n910) );
  XOR2_X1 U992 ( .A(G2446), .B(KEYINPUT109), .Z(n902) );
  XNOR2_X1 U993 ( .A(KEYINPUT110), .B(G2438), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U998 ( .A(n906), .B(n905), .Z(n908) );
  XNOR2_X1 U999 ( .A(G2430), .B(G2427), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(n911), .A2(G14), .ZN(n919) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n919), .ZN(n914) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n912), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1007 ( .A1(G397), .A2(G395), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(G225) );
  XOR2_X1 U1009 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  INV_X1 U1013 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G325) );
  INV_X1 U1015 ( .A(G325), .ZN(G261) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(n919), .ZN(G401) );
  XNOR2_X1 U1018 ( .A(G16), .B(KEYINPUT56), .ZN(n944) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT57), .ZN(n942) );
  XOR2_X1 U1022 ( .A(G1341), .B(KEYINPUT124), .Z(n923) );
  XNOR2_X1 U1023 ( .A(n924), .B(n923), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n940) );
  XNOR2_X1 U1026 ( .A(n927), .B(G1348), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1956), .B(n928), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(G1961), .B(G301), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n970) );
  INV_X1 U1037 ( .A(G16), .ZN(n968) );
  XOR2_X1 U1038 ( .A(G1956), .B(G20), .Z(n950) );
  XOR2_X1 U1039 ( .A(G1341), .B(G19), .Z(n945) );
  XNOR2_X1 U1040 ( .A(KEYINPUT125), .B(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(G6), .B(G1981), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT126), .B(n948), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1045 ( .A(KEYINPUT59), .B(G1348), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G4), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n954), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G21), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G5), .B(G1961), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n965) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n962) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT61), .B(n966), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n993) );
  XOR2_X1 U1063 ( .A(G29), .B(KEYINPUT122), .Z(n989) );
  XOR2_X1 U1064 ( .A(G25), .B(G1991), .Z(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(G28), .ZN(n980) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G26), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G33), .B(G2072), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G32), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G27), .B(n974), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1074 ( .A(KEYINPUT53), .B(n981), .Z(n984) );
  XOR2_X1 U1075 ( .A(KEYINPUT54), .B(G34), .Z(n982) );
  XNOR2_X1 U1076 ( .A(G2084), .B(n982), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G35), .B(G2090), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n987), .B(KEYINPUT55), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(G11), .A2(n990), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT123), .B(n991), .Z(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(n994), .B(KEYINPUT127), .ZN(n1026) );
  INV_X1 U1086 ( .A(G29), .ZN(n1024) );
  XOR2_X1 U1087 ( .A(G2072), .B(n995), .Z(n997) );
  XOR2_X1 U1088 ( .A(G164), .B(G2078), .Z(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1090 ( .A(n998), .B(KEYINPUT50), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(n999), .B(KEYINPUT121), .ZN(n1020) );
  XOR2_X1 U1092 ( .A(G160), .B(G2084), .Z(n1004) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(KEYINPUT117), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT118), .B(n1005), .Z(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT119), .B(n1008), .Z(n1013) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1101 ( .A(KEYINPUT51), .B(n1011), .Z(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT120), .B(n1018), .Z(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1107 ( .A(KEYINPUT52), .B(n1021), .Z(n1022) );
  NOR2_X1 U1108 ( .A1(KEYINPUT55), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
  INV_X1 U1113 ( .A(G301), .ZN(G171) );
endmodule

