

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U558 ( .A(KEYINPUT13), .B(n579), .Z(n522) );
  NOR2_X2 U559 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n781) );
  NOR2_X2 U561 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X2 U562 ( .A(n706), .B(n705), .ZN(n707) );
  INV_X1 U563 ( .A(KEYINPUT98), .ZN(n705) );
  AND2_X1 U564 ( .A1(n716), .A2(G1341), .ZN(n523) );
  INV_X1 U565 ( .A(G168), .ZN(n720) );
  XNOR2_X1 U566 ( .A(n715), .B(n714), .ZN(n777) );
  NAND2_X1 U567 ( .A1(G160), .A2(G40), .ZN(n780) );
  NOR2_X2 U568 ( .A1(n639), .A2(n548), .ZN(n646) );
  NAND2_X1 U569 ( .A1(n582), .A2(n581), .ZN(n972) );
  XNOR2_X1 U570 ( .A(n524), .B(KEYINPUT64), .ZN(n526) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n525) );
  XNOR2_X1 U572 ( .A(n526), .B(n525), .ZN(n606) );
  NAND2_X1 U573 ( .A1(n606), .A2(G138), .ZN(n534) );
  INV_X1 U574 ( .A(G2104), .ZN(n527) );
  AND2_X1 U575 ( .A1(n527), .A2(G2105), .ZN(n898) );
  NAND2_X1 U576 ( .A1(G126), .A2(n898), .ZN(n529) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n899) );
  NAND2_X1 U578 ( .A1(G114), .A2(n899), .ZN(n528) );
  AND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n532) );
  INV_X1 U580 ( .A(G2105), .ZN(n530) );
  AND2_X4 U581 ( .A1(n530), .A2(G2104), .ZN(n537) );
  NAND2_X1 U582 ( .A1(n537), .A2(G102), .ZN(n531) );
  AND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n533) );
  AND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(G164) );
  NAND2_X1 U585 ( .A1(G137), .A2(n606), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n899), .A2(G113), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U588 ( .A1(n898), .A2(G125), .ZN(n540) );
  NAND2_X1 U589 ( .A1(G101), .A2(n537), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT23), .B(n538), .Z(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U592 ( .A1(n542), .A2(n541), .ZN(G160) );
  NOR2_X1 U593 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U594 ( .A1(n650), .A2(G89), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT4), .ZN(n546) );
  XNOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n544), .B(KEYINPUT67), .ZN(n639) );
  INV_X1 U598 ( .A(G651), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G76), .A2(n646), .ZN(n545) );
  NAND2_X1 U600 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U601 ( .A(KEYINPUT5), .B(n547), .ZN(n556) );
  XNOR2_X1 U602 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n554) );
  NOR2_X2 U603 ( .A1(G651), .A2(n639), .ZN(n647) );
  NAND2_X1 U604 ( .A1(n647), .A2(G51), .ZN(n552) );
  NOR2_X1 U605 ( .A1(G543), .A2(n548), .ZN(n549) );
  XOR2_X2 U606 ( .A(KEYINPUT1), .B(n549), .Z(n654) );
  NAND2_X1 U607 ( .A1(n654), .A2(G63), .ZN(n550) );
  XOR2_X1 U608 ( .A(KEYINPUT73), .B(n550), .Z(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(n554), .B(n553), .Z(n555) );
  NAND2_X1 U611 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U612 ( .A(KEYINPUT7), .B(n557), .ZN(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U614 ( .A1(G65), .A2(n654), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G53), .A2(n647), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U617 ( .A1(G91), .A2(n650), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G78), .A2(n646), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  OR2_X1 U620 ( .A1(n563), .A2(n562), .ZN(G299) );
  NAND2_X1 U621 ( .A1(G64), .A2(n654), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G52), .A2(n647), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U624 ( .A(KEYINPUT68), .B(n566), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G90), .A2(n650), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G77), .A2(n646), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n569), .Z(n570) );
  NOR2_X1 U629 ( .A1(n571), .A2(n570), .ZN(G171) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G57), .ZN(G237) );
  XOR2_X1 U632 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n573) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n573), .B(n572), .ZN(G223) );
  INV_X1 U635 ( .A(G223), .ZN(n834) );
  NAND2_X1 U636 ( .A1(n834), .A2(G567), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n654), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n575), .Z(n580) );
  NAND2_X1 U640 ( .A1(n650), .A2(G81), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G68), .A2(n646), .ZN(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n522), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n647), .A2(G43), .ZN(n581) );
  INV_X1 U646 ( .A(G860), .ZN(n614) );
  OR2_X1 U647 ( .A1(n972), .A2(n614), .ZN(G153) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G79), .A2(n646), .ZN(n584) );
  NAND2_X1 U650 ( .A1(G54), .A2(n647), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U652 ( .A1(G92), .A2(n650), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G66), .A2(n654), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n589), .B(KEYINPUT15), .ZN(n699) );
  NOR2_X1 U657 ( .A1(G868), .A2(n699), .ZN(n591) );
  INV_X1 U658 ( .A(G868), .ZN(n666) );
  NOR2_X1 U659 ( .A1(n666), .A2(G301), .ZN(n590) );
  NOR2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U661 ( .A(KEYINPUT72), .B(n592), .ZN(G284) );
  NOR2_X1 U662 ( .A1(G286), .A2(n666), .ZN(n593) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n593), .Z(n595) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n614), .A2(G559), .ZN(n596) );
  INV_X1 U667 ( .A(n699), .ZN(n981) );
  NAND2_X1 U668 ( .A1(n596), .A2(n981), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U670 ( .A1(n981), .A2(G868), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G559), .A2(n598), .ZN(n599) );
  XNOR2_X1 U672 ( .A(n599), .B(KEYINPUT76), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n972), .A2(G868), .ZN(n600) );
  NOR2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G123), .A2(n898), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT77), .B(n602), .Z(n603) );
  XNOR2_X1 U677 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G99), .A2(n537), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n899), .A2(G111), .ZN(n608) );
  BUF_X1 U681 ( .A(n606), .Z(n902) );
  NAND2_X1 U682 ( .A1(G135), .A2(n902), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n930) );
  XNOR2_X1 U685 ( .A(G2096), .B(n930), .ZN(n612) );
  INV_X1 U686 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(G156) );
  XOR2_X1 U688 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n616) );
  NAND2_X1 U689 ( .A1(G559), .A2(n981), .ZN(n613) );
  XOR2_X1 U690 ( .A(n972), .B(n613), .Z(n663) );
  NAND2_X1 U691 ( .A1(n663), .A2(n614), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n616), .B(n615), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G93), .A2(n650), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G67), .A2(n654), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G80), .A2(n646), .ZN(n619) );
  XNOR2_X1 U697 ( .A(KEYINPUT79), .B(n619), .ZN(n620) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n647), .A2(G55), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n665) );
  XOR2_X1 U701 ( .A(n624), .B(n665), .Z(G145) );
  NAND2_X1 U702 ( .A1(G88), .A2(n650), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G75), .A2(n646), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G62), .A2(n654), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G50), .A2(n647), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U708 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G61), .A2(n654), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT82), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G86), .A2(n650), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G48), .A2(n647), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n646), .A2(G73), .ZN(n634) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n634), .Z(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G87), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U721 ( .A1(n654), .A2(n642), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G49), .A2(n647), .ZN(n643) );
  XOR2_X1 U723 ( .A(KEYINPUT81), .B(n643), .Z(n644) );
  NAND2_X1 U724 ( .A1(n645), .A2(n644), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G72), .A2(n646), .ZN(n649) );
  NAND2_X1 U726 ( .A1(G47), .A2(n647), .ZN(n648) );
  NAND2_X1 U727 ( .A1(n649), .A2(n648), .ZN(n653) );
  NAND2_X1 U728 ( .A1(G85), .A2(n650), .ZN(n651) );
  XOR2_X1 U729 ( .A(KEYINPUT66), .B(n651), .Z(n652) );
  NOR2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n654), .A2(G60), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(G290) );
  XOR2_X1 U733 ( .A(G305), .B(G288), .Z(n657) );
  XNOR2_X1 U734 ( .A(n665), .B(n657), .ZN(n658) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(n658), .ZN(n660) );
  XNOR2_X1 U736 ( .A(G290), .B(KEYINPUT83), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U738 ( .A(G166), .B(n661), .Z(n662) );
  XNOR2_X1 U739 ( .A(G299), .B(n662), .ZN(n914) );
  XNOR2_X1 U740 ( .A(n663), .B(n914), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U743 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U745 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U746 ( .A1(n670), .A2(G2090), .ZN(n671) );
  XNOR2_X1 U747 ( .A(n671), .B(KEYINPUT84), .ZN(n672) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U749 ( .A1(G2072), .A2(n673), .ZN(G158) );
  XOR2_X1 U750 ( .A(KEYINPUT85), .B(G44), .Z(n674) );
  XNOR2_X1 U751 ( .A(KEYINPUT3), .B(n674), .ZN(G218) );
  XOR2_X1 U752 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  XNOR2_X1 U753 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n676) );
  XNOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT86), .ZN(n675) );
  XNOR2_X1 U756 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n677), .A2(G96), .ZN(n678) );
  NOR2_X1 U758 ( .A1(G218), .A2(n678), .ZN(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT87), .B(n679), .ZN(n839) );
  NAND2_X1 U760 ( .A1(n839), .A2(G2106), .ZN(n683) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G108), .A2(n681), .ZN(n840) );
  NAND2_X1 U764 ( .A1(n840), .A2(G567), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n872) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n872), .A2(n684), .ZN(n838) );
  NAND2_X1 U768 ( .A1(n838), .A2(G36), .ZN(G176) );
  XOR2_X1 U769 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  INV_X1 U770 ( .A(n780), .ZN(n686) );
  AND2_X1 U771 ( .A1(n781), .A2(n686), .ZN(n693) );
  NAND2_X1 U772 ( .A1(n693), .A2(G2072), .ZN(n685) );
  XOR2_X1 U773 ( .A(KEYINPUT27), .B(n685), .Z(n688) );
  NAND2_X1 U774 ( .A1(n781), .A2(n686), .ZN(n716) );
  NAND2_X1 U775 ( .A1(G1956), .A2(n716), .ZN(n687) );
  NAND2_X1 U776 ( .A1(n688), .A2(n687), .ZN(n702) );
  NAND2_X1 U777 ( .A1(G299), .A2(n702), .ZN(n689) );
  XOR2_X1 U778 ( .A(KEYINPUT28), .B(n689), .Z(n708) );
  NOR2_X1 U779 ( .A1(n972), .A2(n523), .ZN(n692) );
  AND2_X1 U780 ( .A1(n693), .A2(G1996), .ZN(n690) );
  XOR2_X1 U781 ( .A(n690), .B(KEYINPUT26), .Z(n691) );
  AND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n697) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n716), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G2067), .A2(n693), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n701) );
  AND2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U790 ( .A1(G299), .A2(n702), .ZN(n703) );
  OR2_X2 U791 ( .A1(n704), .A2(n703), .ZN(n706) );
  NOR2_X2 U792 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U793 ( .A(n709), .B(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U794 ( .A(G2078), .B(KEYINPUT25), .ZN(n957) );
  NOR2_X1 U795 ( .A1(n716), .A2(n957), .ZN(n711) );
  INV_X1 U796 ( .A(G1961), .ZN(n999) );
  NOR2_X1 U797 ( .A1(n693), .A2(n999), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n722) );
  NAND2_X1 U799 ( .A1(n722), .A2(G171), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n727) );
  NAND2_X1 U801 ( .A1(n716), .A2(G8), .ZN(n715) );
  INV_X1 U802 ( .A(KEYINPUT95), .ZN(n714) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n777), .ZN(n741) );
  NOR2_X1 U804 ( .A1(n716), .A2(G2084), .ZN(n717) );
  XNOR2_X1 U805 ( .A(n717), .B(KEYINPUT97), .ZN(n737) );
  NAND2_X1 U806 ( .A1(G8), .A2(n737), .ZN(n718) );
  NOR2_X1 U807 ( .A1(n741), .A2(n718), .ZN(n719) );
  XNOR2_X1 U808 ( .A(n719), .B(KEYINPUT30), .ZN(n721) );
  AND2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n724) );
  NOR2_X1 U810 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U811 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U812 ( .A(KEYINPUT31), .B(n725), .Z(n726) );
  NAND2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n739), .A2(G286), .ZN(n733) );
  NOR2_X1 U815 ( .A1(G2090), .A2(n716), .ZN(n728) );
  XOR2_X1 U816 ( .A(KEYINPUT99), .B(n728), .Z(n730) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n777), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n731), .A2(G303), .ZN(n732) );
  NAND2_X1 U820 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT100), .ZN(n735) );
  NAND2_X1 U822 ( .A1(n735), .A2(G8), .ZN(n736) );
  XNOR2_X1 U823 ( .A(n736), .B(KEYINPUT32), .ZN(n745) );
  INV_X1 U824 ( .A(n737), .ZN(n738) );
  NAND2_X1 U825 ( .A1(G8), .A2(n738), .ZN(n743) );
  INV_X1 U826 ( .A(n739), .ZN(n740) );
  NOR2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n753) );
  NOR2_X1 U830 ( .A1(G2090), .A2(G303), .ZN(n746) );
  NAND2_X1 U831 ( .A1(G8), .A2(n746), .ZN(n747) );
  NAND2_X1 U832 ( .A1(n753), .A2(n747), .ZN(n749) );
  INV_X1 U833 ( .A(KEYINPUT104), .ZN(n748) );
  XNOR2_X1 U834 ( .A(n749), .B(n748), .ZN(n751) );
  INV_X1 U835 ( .A(n777), .ZN(n750) );
  XNOR2_X1 U836 ( .A(n752), .B(KEYINPUT105), .ZN(n772) );
  INV_X1 U837 ( .A(n753), .ZN(n758) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n754) );
  XOR2_X1 U839 ( .A(KEYINPUT101), .B(n754), .Z(n977) );
  NOR2_X1 U840 ( .A1(G303), .A2(G1971), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n977), .A2(n755), .ZN(n756) );
  XOR2_X1 U842 ( .A(KEYINPUT102), .B(n756), .Z(n757) );
  NOR2_X1 U843 ( .A1(n758), .A2(n757), .ZN(n761) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U845 ( .A1(KEYINPUT103), .A2(n777), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n978), .A2(n759), .ZN(n760) );
  NOR2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n762), .ZN(n769) );
  INV_X1 U849 ( .A(KEYINPUT103), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n977), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n977), .A2(KEYINPUT103), .ZN(n765) );
  NAND2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n777), .A2(n767), .ZN(n768) );
  NOR2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U856 ( .A(G1981), .B(G305), .Z(n973) );
  NAND2_X1 U857 ( .A1(n770), .A2(n973), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT106), .ZN(n779) );
  NOR2_X1 U860 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U861 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  XNOR2_X1 U862 ( .A(KEYINPUT96), .B(n775), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n779), .A2(n778), .ZN(n815) );
  NOR2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n828) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  XNOR2_X1 U867 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n793) );
  NAND2_X1 U868 ( .A1(G128), .A2(n898), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G116), .A2(n899), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(KEYINPUT35), .B(n784), .ZN(n791) );
  XNOR2_X1 U872 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n789) );
  NAND2_X1 U873 ( .A1(n537), .A2(G104), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G140), .A2(n902), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U876 ( .A(n787), .B(KEYINPUT34), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n789), .B(n788), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n793), .B(n792), .ZN(n911) );
  NOR2_X1 U880 ( .A1(n826), .A2(n911), .ZN(n946) );
  NAND2_X1 U881 ( .A1(n828), .A2(n946), .ZN(n824) );
  NAND2_X1 U882 ( .A1(G119), .A2(n898), .ZN(n794) );
  XNOR2_X1 U883 ( .A(n794), .B(KEYINPUT92), .ZN(n801) );
  NAND2_X1 U884 ( .A1(n537), .A2(G95), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G131), .A2(n902), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G107), .A2(n899), .ZN(n797) );
  XNOR2_X1 U888 ( .A(KEYINPUT93), .B(n797), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n801), .A2(n800), .ZN(n888) );
  AND2_X1 U891 ( .A1(n888), .A2(G1991), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G105), .A2(n537), .ZN(n802) );
  XNOR2_X1 U893 ( .A(n802), .B(KEYINPUT38), .ZN(n809) );
  NAND2_X1 U894 ( .A1(n899), .A2(G117), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G141), .A2(n902), .ZN(n803) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n898), .A2(G129), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT94), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n889) );
  AND2_X1 U901 ( .A1(n889), .A2(G1996), .ZN(n810) );
  NOR2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n937) );
  INV_X1 U903 ( .A(n828), .ZN(n812) );
  NOR2_X1 U904 ( .A1(n937), .A2(n812), .ZN(n821) );
  INV_X1 U905 ( .A(n821), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n824), .A2(n813), .ZN(n814) );
  NOR2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n817) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n983) );
  NAND2_X1 U909 ( .A1(n983), .A2(n828), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n831) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n889), .ZN(n818) );
  XOR2_X1 U912 ( .A(KEYINPUT107), .B(n818), .Z(n939) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n888), .ZN(n931) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n931), .A2(n819), .ZN(n820) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n939), .A2(n822), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n826), .A2(n911), .ZN(n943) );
  NAND2_X1 U921 ( .A1(n827), .A2(n943), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n833) );
  XNOR2_X1 U924 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n834), .ZN(G217) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n835) );
  XNOR2_X1 U928 ( .A(KEYINPUT111), .B(n835), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n836), .A2(G661), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(KEYINPUT112), .B(KEYINPUT114), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2678), .B(G2096), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n843), .B(KEYINPUT113), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U944 ( .A(G2100), .B(G2090), .Z(n847) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U950 ( .A(G1956), .B(G1961), .Z(n853) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1976), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U953 ( .A(n854), .B(KEYINPUT41), .Z(n856) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U956 ( .A(G2474), .B(G1971), .Z(n858) );
  XNOR2_X1 U957 ( .A(G1981), .B(G1966), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U960 ( .A(G2430), .B(G2451), .Z(n862) );
  XNOR2_X1 U961 ( .A(G2446), .B(G2427), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n869) );
  XOR2_X1 U963 ( .A(G2438), .B(G2435), .Z(n864) );
  XNOR2_X1 U964 ( .A(G2443), .B(KEYINPUT109), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U966 ( .A(n865), .B(G2454), .Z(n867) );
  XNOR2_X1 U967 ( .A(G1341), .B(G1348), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n870), .A2(G14), .ZN(n871) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n871), .Z(G401) );
  INV_X1 U972 ( .A(n872), .ZN(G319) );
  NAND2_X1 U973 ( .A1(G124), .A2(n898), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n537), .A2(G100), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n899), .A2(G112), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G136), .A2(n902), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U980 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U981 ( .A1(n537), .A2(G103), .ZN(n881) );
  NAND2_X1 U982 ( .A1(G139), .A2(n902), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n887) );
  NAND2_X1 U984 ( .A1(G127), .A2(n898), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G115), .A2(n899), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U987 ( .A(KEYINPUT116), .B(n884), .Z(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n885), .ZN(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n926) );
  XNOR2_X1 U990 ( .A(n926), .B(n888), .ZN(n891) );
  XOR2_X1 U991 ( .A(G160), .B(n889), .Z(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U993 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  XNOR2_X1 U994 ( .A(n930), .B(KEYINPUT115), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U996 ( .A(n895), .B(n894), .Z(n897) );
  XNOR2_X1 U997 ( .A(G164), .B(G162), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n909) );
  NAND2_X1 U999 ( .A1(G130), .A2(n898), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n899), .ZN(n900) );
  NAND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n537), .A2(G106), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n902), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(n905), .B(KEYINPUT45), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(n909), .B(n908), .Z(n910) );
  XOR2_X1 U1008 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n912), .ZN(n913) );
  XOR2_X1 U1010 ( .A(KEYINPUT117), .B(n913), .Z(G395) );
  XOR2_X1 U1011 ( .A(n914), .B(G286), .Z(n916) );
  XNOR2_X1 U1012 ( .A(G171), .B(n981), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1014 ( .A(n917), .B(n972), .Z(n918) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(n919), .Z(n920) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n920), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n921) );
  XOR2_X1 U1020 ( .A(KEYINPUT119), .B(n921), .Z(n922) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(G401), .A2(n923), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1026 ( .A(G2072), .B(n926), .Z(n928) );
  XOR2_X1 U1027 ( .A(G164), .B(G2078), .Z(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n929), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G160), .B(G2084), .Z(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n940), .B(KEYINPUT51), .ZN(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n967), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n956) );
  XOR2_X1 U1049 ( .A(G25), .B(G1991), .Z(n952) );
  NAND2_X1 U1050 ( .A1(n952), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1054 ( .A(G27), .B(n957), .Z(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(n967), .B(n966), .ZN(n969) );
  INV_X1 U1062 ( .A(G29), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n970), .ZN(n1028) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XOR2_X1 U1066 ( .A(G1341), .B(KEYINPUT124), .Z(n971) );
  XNOR2_X1 U1067 ( .A(n972), .B(n971), .ZN(n996) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n974) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(KEYINPUT120), .ZN(n976) );
  XOR2_X1 U1071 ( .A(KEYINPUT57), .B(n976), .Z(n994) );
  XNOR2_X1 U1072 ( .A(n977), .B(KEYINPUT121), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(n980), .B(KEYINPUT122), .ZN(n991) );
  XNOR2_X1 U1075 ( .A(G171), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(n981), .B(G1348), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(G1956), .B(G299), .ZN(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G303), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1026) );
  INV_X1 U1088 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1089 ( .A(G5), .B(n999), .ZN(n1013) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1000), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(n1001), .B(G1348), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(G20), .B(G1956), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1099 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1100 ( .A(n1008), .B(KEYINPUT126), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(G1986), .B(G24), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(G22), .B(G1971), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G1976), .B(KEYINPUT127), .ZN(n1016) );
  XNOR2_X1 U1108 ( .A(n1016), .B(G23), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1110 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

