

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X4 U551 ( .A1(n531), .A2(n530), .ZN(G160) );
  NOR2_X1 U552 ( .A1(n815), .A2(n796), .ZN(n517) );
  AND2_X1 U553 ( .A1(n806), .A2(n805), .ZN(n518) );
  OR2_X1 U554 ( .A1(n787), .A2(n768), .ZN(n769) );
  XNOR2_X1 U555 ( .A(n769), .B(KEYINPUT30), .ZN(n770) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n751) );
  XNOR2_X1 U557 ( .A(n752), .B(n751), .ZN(n757) );
  AND2_X1 U558 ( .A1(n785), .A2(n776), .ZN(n775) );
  INV_X1 U559 ( .A(KEYINPUT106), .ZN(n799) );
  INV_X1 U560 ( .A(KEYINPUT17), .ZN(n521) );
  XNOR2_X1 U561 ( .A(n521), .B(KEYINPUT66), .ZN(n522) );
  NOR2_X1 U562 ( .A1(n821), .A2(n820), .ZN(n823) );
  NOR2_X1 U563 ( .A1(G651), .A2(n629), .ZN(n660) );
  XOR2_X1 U564 ( .A(KEYINPUT64), .B(G2104), .Z(n527) );
  NOR2_X4 U565 ( .A1(n527), .A2(G2105), .ZN(n993) );
  NAND2_X1 U566 ( .A1(G101), .A2(n993), .ZN(n519) );
  XNOR2_X1 U567 ( .A(n519), .B(KEYINPUT65), .ZN(n520) );
  XNOR2_X1 U568 ( .A(KEYINPUT23), .B(n520), .ZN(n526) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X2 U570 ( .A(n523), .B(n522), .ZN(n994) );
  NAND2_X1 U571 ( .A1(n994), .A2(G137), .ZN(n524) );
  XOR2_X1 U572 ( .A(KEYINPUT67), .B(n524), .Z(n525) );
  NAND2_X1 U573 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U574 ( .A1(n527), .A2(G2105), .ZN(n989) );
  NAND2_X1 U575 ( .A1(G125), .A2(n989), .ZN(n529) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n990) );
  NAND2_X1 U577 ( .A1(G113), .A2(n990), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U580 ( .A1(n653), .A2(G89), .ZN(n532) );
  XNOR2_X1 U581 ( .A(n532), .B(KEYINPUT4), .ZN(n535) );
  XNOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .ZN(n533) );
  XNOR2_X1 U583 ( .A(n533), .B(KEYINPUT69), .ZN(n629) );
  INV_X1 U584 ( .A(G651), .ZN(n538) );
  NOR2_X1 U585 ( .A1(n629), .A2(n538), .ZN(n650) );
  NAND2_X1 U586 ( .A1(G76), .A2(n650), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U588 ( .A(KEYINPUT5), .B(n536), .ZN(n544) );
  NAND2_X1 U589 ( .A1(n660), .A2(G51), .ZN(n537) );
  XOR2_X1 U590 ( .A(KEYINPUT81), .B(n537), .Z(n541) );
  NOR2_X1 U591 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n539), .Z(n654) );
  NAND2_X1 U593 ( .A1(n654), .A2(G63), .ZN(n540) );
  NAND2_X1 U594 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U597 ( .A(KEYINPUT7), .B(n545), .ZN(G168) );
  XOR2_X1 U598 ( .A(G2443), .B(G2446), .Z(n547) );
  XNOR2_X1 U599 ( .A(G2427), .B(G2451), .ZN(n546) );
  XNOR2_X1 U600 ( .A(n547), .B(n546), .ZN(n553) );
  XOR2_X1 U601 ( .A(G2430), .B(G2454), .Z(n549) );
  XNOR2_X1 U602 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U604 ( .A(G2435), .B(G2438), .Z(n550) );
  XNOR2_X1 U605 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U606 ( .A(n553), .B(n552), .Z(n554) );
  AND2_X1 U607 ( .A1(G14), .A2(n554), .ZN(G401) );
  NAND2_X1 U608 ( .A1(n989), .A2(G126), .ZN(n556) );
  NAND2_X1 U609 ( .A1(G138), .A2(n994), .ZN(n555) );
  NAND2_X1 U610 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U611 ( .A1(G114), .A2(n990), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G102), .A2(n993), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n560), .A2(n559), .ZN(G164) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  XOR2_X1 U616 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U617 ( .A1(G94), .A2(G452), .ZN(n561) );
  XNOR2_X1 U618 ( .A(n561), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n562), .B(KEYINPUT10), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT78), .B(n563), .ZN(G223) );
  INV_X1 U622 ( .A(G223), .ZN(n840) );
  NAND2_X1 U623 ( .A1(n840), .A2(G567), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U625 ( .A1(G56), .A2(n654), .ZN(n565) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(n565), .Z(n572) );
  NAND2_X1 U627 ( .A1(G81), .A2(n653), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT79), .B(n566), .Z(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G68), .A2(n650), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n570), .Z(n571) );
  NOR2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n660), .A2(G43), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n1018) );
  INV_X1 U636 ( .A(G860), .ZN(n620) );
  OR2_X1 U637 ( .A1(n1018), .A2(n620), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G90), .A2(n653), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G77), .A2(n650), .ZN(n575) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT9), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G64), .A2(n654), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G52), .A2(n660), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT71), .B(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(KEYINPUT72), .B(n583), .ZN(G171) );
  INV_X1 U648 ( .A(G171), .ZN(G301) );
  NAND2_X1 U649 ( .A1(G301), .A2(G868), .ZN(n593) );
  NAND2_X1 U650 ( .A1(G92), .A2(n653), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G66), .A2(n654), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G79), .A2(n650), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G54), .A2(n660), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT80), .B(n588), .ZN(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT15), .ZN(n1021) );
  INV_X1 U659 ( .A(G868), .ZN(n671) );
  NAND2_X1 U660 ( .A1(n1021), .A2(n671), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U662 ( .A1(n653), .A2(G91), .ZN(n594) );
  XNOR2_X1 U663 ( .A(n594), .B(KEYINPUT74), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G65), .A2(n654), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U666 ( .A1(G78), .A2(n650), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G53), .A2(n660), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n909) );
  XNOR2_X1 U670 ( .A(n909), .B(KEYINPUT75), .ZN(G299) );
  NAND2_X1 U671 ( .A1(G286), .A2(G868), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G299), .A2(n671), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n620), .A2(G559), .ZN(n603) );
  INV_X1 U675 ( .A(n1021), .ZN(n618) );
  NAND2_X1 U676 ( .A1(n603), .A2(n618), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U678 ( .A1(n618), .A2(G868), .ZN(n605) );
  NOR2_X1 U679 ( .A1(G559), .A2(n605), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT82), .ZN(n608) );
  NOR2_X1 U681 ( .A1(n1018), .A2(G868), .ZN(n607) );
  NOR2_X1 U682 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U683 ( .A1(n990), .A2(G111), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G135), .A2(n994), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U686 ( .A1(n989), .A2(G123), .ZN(n611) );
  XNOR2_X1 U687 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G99), .A2(n993), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n1005) );
  XNOR2_X1 U691 ( .A(n1005), .B(G2096), .ZN(n617) );
  INV_X1 U692 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G559), .A2(n618), .ZN(n619) );
  XOR2_X1 U695 ( .A(n1018), .B(n619), .Z(n669) );
  NAND2_X1 U696 ( .A1(n620), .A2(n669), .ZN(n628) );
  NAND2_X1 U697 ( .A1(G93), .A2(n653), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G67), .A2(n654), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G55), .A2(n660), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT83), .B(n623), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n650), .A2(G80), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n672) );
  XNOR2_X1 U705 ( .A(n628), .B(n672), .ZN(G145) );
  NAND2_X1 U706 ( .A1(G49), .A2(n660), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G87), .A2(n629), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U709 ( .A1(n654), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G651), .A2(G74), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G72), .A2(n650), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G47), .A2(n660), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G85), .A2(n653), .ZN(n637) );
  XOR2_X1 U716 ( .A(KEYINPUT68), .B(n637), .Z(n638) );
  NOR2_X1 U717 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n654), .A2(G60), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U720 ( .A(KEYINPUT70), .B(n642), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G75), .A2(n650), .ZN(n644) );
  NAND2_X1 U722 ( .A1(G50), .A2(n660), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G88), .A2(n653), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G62), .A2(n654), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(KEYINPUT86), .ZN(G166) );
  XOR2_X1 U729 ( .A(KEYINPUT84), .B(KEYINPUT2), .Z(n652) );
  NAND2_X1 U730 ( .A1(G73), .A2(n650), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n652), .B(n651), .ZN(n658) );
  NAND2_X1 U732 ( .A1(G86), .A2(n653), .ZN(n656) );
  NAND2_X1 U733 ( .A1(G61), .A2(n654), .ZN(n655) );
  NAND2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT85), .B(n659), .Z(n662) );
  NAND2_X1 U737 ( .A1(n660), .A2(G48), .ZN(n661) );
  NAND2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G305) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(G288), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n663), .B(n672), .ZN(n666) );
  XNOR2_X1 U741 ( .A(G290), .B(G166), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n664), .B(G299), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n668) );
  XNOR2_X1 U744 ( .A(G305), .B(KEYINPUT87), .ZN(n667) );
  XNOR2_X1 U745 ( .A(n668), .B(n667), .ZN(n1017) );
  XNOR2_X1 U746 ( .A(n669), .B(n1017), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n678), .A2(G2072), .ZN(n679) );
  XNOR2_X1 U755 ( .A(KEYINPUT88), .B(n679), .ZN(G158) );
  XOR2_X1 U756 ( .A(KEYINPUT76), .B(G57), .Z(G237) );
  XOR2_X1 U757 ( .A(KEYINPUT89), .B(G44), .Z(n680) );
  XNOR2_X1 U758 ( .A(KEYINPUT3), .B(n680), .ZN(G218) );
  XNOR2_X1 U759 ( .A(KEYINPUT77), .B(G82), .ZN(G220) );
  NAND2_X1 U760 ( .A1(G108), .A2(G120), .ZN(n681) );
  NOR2_X1 U761 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(G69), .A2(n682), .ZN(n968) );
  NAND2_X1 U763 ( .A1(n968), .A2(G567), .ZN(n687) );
  NOR2_X1 U764 ( .A1(G219), .A2(G220), .ZN(n683) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U766 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G96), .A2(n685), .ZN(n967) );
  NAND2_X1 U768 ( .A1(n967), .A2(G2106), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n687), .A2(n686), .ZN(n988) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n988), .A2(n688), .ZN(n844) );
  NAND2_X1 U772 ( .A1(n844), .A2(G36), .ZN(G176) );
  INV_X1 U773 ( .A(G166), .ZN(G303) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n727) );
  AND2_X2 U775 ( .A1(G160), .A2(G40), .ZN(n728) );
  INV_X1 U776 ( .A(n728), .ZN(n690) );
  NOR2_X1 U777 ( .A1(n727), .A2(n690), .ZN(n834) );
  NAND2_X1 U778 ( .A1(n993), .A2(G104), .ZN(n692) );
  NAND2_X1 U779 ( .A1(G140), .A2(n994), .ZN(n691) );
  NAND2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT34), .B(n693), .ZN(n701) );
  XNOR2_X1 U782 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n990), .A2(G116), .ZN(n694) );
  XNOR2_X1 U784 ( .A(n694), .B(KEYINPUT90), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G128), .A2(n989), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n697), .B(KEYINPUT35), .ZN(n698) );
  XNOR2_X1 U788 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U790 ( .A(n702), .B(KEYINPUT36), .ZN(n1010) );
  XNOR2_X1 U791 ( .A(G2067), .B(KEYINPUT37), .ZN(n832) );
  NOR2_X1 U792 ( .A1(n1010), .A2(n832), .ZN(n854) );
  NAND2_X1 U793 ( .A1(n834), .A2(n854), .ZN(n830) );
  NAND2_X1 U794 ( .A1(n990), .A2(G107), .ZN(n704) );
  NAND2_X1 U795 ( .A1(G131), .A2(n994), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X1 U797 ( .A1(G119), .A2(n989), .ZN(n706) );
  NAND2_X1 U798 ( .A1(G95), .A2(n993), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  OR2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n1006) );
  NAND2_X1 U801 ( .A1(G1991), .A2(n1006), .ZN(n718) );
  NAND2_X1 U802 ( .A1(G105), .A2(n993), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n709), .B(KEYINPUT38), .ZN(n716) );
  NAND2_X1 U804 ( .A1(n989), .A2(G129), .ZN(n711) );
  NAND2_X1 U805 ( .A1(G141), .A2(n994), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U807 ( .A1(G117), .A2(n990), .ZN(n712) );
  XNOR2_X1 U808 ( .A(KEYINPUT93), .B(n712), .ZN(n713) );
  NOR2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n1004) );
  NAND2_X1 U811 ( .A1(G1996), .A2(n1004), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U813 ( .A(KEYINPUT94), .B(n719), .Z(n857) );
  INV_X1 U814 ( .A(n857), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n834), .A2(n720), .ZN(n824) );
  NAND2_X1 U816 ( .A1(n830), .A2(n824), .ZN(n821) );
  NAND2_X1 U817 ( .A1(n727), .A2(n728), .ZN(n758) );
  INV_X1 U818 ( .A(G2072), .ZN(n871) );
  NOR2_X1 U819 ( .A1(n758), .A2(n871), .ZN(n724) );
  INV_X1 U820 ( .A(n724), .ZN(n722) );
  XNOR2_X1 U821 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n723) );
  INV_X1 U822 ( .A(n723), .ZN(n721) );
  NAND2_X1 U823 ( .A1(n722), .A2(n721), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n730) );
  AND2_X1 U826 ( .A1(n728), .A2(n727), .ZN(n738) );
  INV_X1 U827 ( .A(n738), .ZN(n760) );
  NAND2_X1 U828 ( .A1(n760), .A2(G1956), .ZN(n729) );
  NAND2_X1 U829 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U830 ( .A(n731), .B(KEYINPUT99), .ZN(n746) );
  NOR2_X1 U831 ( .A1(n746), .A2(n909), .ZN(n733) );
  XOR2_X1 U832 ( .A(KEYINPUT28), .B(KEYINPUT100), .Z(n732) );
  XNOR2_X1 U833 ( .A(n733), .B(n732), .ZN(n750) );
  INV_X1 U834 ( .A(G1996), .ZN(n890) );
  NOR2_X1 U835 ( .A1(n758), .A2(n890), .ZN(n734) );
  XOR2_X1 U836 ( .A(n734), .B(KEYINPUT26), .Z(n736) );
  NAND2_X1 U837 ( .A1(n760), .A2(G1341), .ZN(n735) );
  NAND2_X1 U838 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U839 ( .A1(n1018), .A2(n737), .ZN(n742) );
  BUF_X1 U840 ( .A(n758), .Z(n767) );
  NAND2_X1 U841 ( .A1(G1348), .A2(n767), .ZN(n740) );
  NAND2_X1 U842 ( .A1(G2067), .A2(n738), .ZN(n739) );
  NAND2_X1 U843 ( .A1(n740), .A2(n739), .ZN(n743) );
  NOR2_X1 U844 ( .A1(n1021), .A2(n743), .ZN(n741) );
  OR2_X1 U845 ( .A1(n742), .A2(n741), .ZN(n745) );
  NAND2_X1 U846 ( .A1(n1021), .A2(n743), .ZN(n744) );
  NAND2_X1 U847 ( .A1(n745), .A2(n744), .ZN(n748) );
  NAND2_X1 U848 ( .A1(n746), .A2(n909), .ZN(n747) );
  NAND2_X1 U849 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U850 ( .A1(n750), .A2(n749), .ZN(n752) );
  XOR2_X1 U851 ( .A(G2078), .B(KEYINPUT25), .Z(n753) );
  XNOR2_X1 U852 ( .A(KEYINPUT97), .B(n753), .ZN(n889) );
  NOR2_X1 U853 ( .A1(n767), .A2(n889), .ZN(n755) );
  AND2_X1 U854 ( .A1(n767), .A2(G1961), .ZN(n754) );
  NOR2_X1 U855 ( .A1(n755), .A2(n754), .ZN(n766) );
  NAND2_X1 U856 ( .A1(G171), .A2(n766), .ZN(n756) );
  NAND2_X1 U857 ( .A1(n757), .A2(n756), .ZN(n785) );
  INV_X1 U858 ( .A(G8), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n758), .A2(G8), .ZN(n759) );
  XOR2_X2 U860 ( .A(KEYINPUT95), .B(n759), .Z(n815) );
  NOR2_X1 U861 ( .A1(G1971), .A2(n815), .ZN(n762) );
  NOR2_X1 U862 ( .A1(G2090), .A2(n760), .ZN(n761) );
  NOR2_X1 U863 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U864 ( .A1(G303), .A2(n763), .ZN(n764) );
  OR2_X1 U865 ( .A1(n765), .A2(n764), .ZN(n776) );
  NOR2_X1 U866 ( .A1(n766), .A2(G171), .ZN(n772) );
  NOR2_X1 U867 ( .A1(n815), .A2(G1966), .ZN(n787) );
  NOR2_X1 U868 ( .A1(G2084), .A2(n767), .ZN(n788) );
  OR2_X1 U869 ( .A1(n788), .A2(n765), .ZN(n768) );
  NOR2_X1 U870 ( .A1(n770), .A2(G168), .ZN(n771) );
  NOR2_X1 U871 ( .A1(n772), .A2(n771), .ZN(n774) );
  XNOR2_X1 U872 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n773) );
  XNOR2_X1 U873 ( .A(n774), .B(n773), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n775), .A2(n784), .ZN(n780) );
  INV_X1 U875 ( .A(n776), .ZN(n778) );
  AND2_X1 U876 ( .A1(G286), .A2(G8), .ZN(n777) );
  OR2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n783) );
  XOR2_X1 U879 ( .A(KEYINPUT32), .B(KEYINPUT102), .Z(n781) );
  XNOR2_X1 U880 ( .A(KEYINPUT103), .B(n781), .ZN(n782) );
  XNOR2_X1 U881 ( .A(n783), .B(n782), .ZN(n792) );
  AND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G8), .A2(n788), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n813) );
  NOR2_X1 U887 ( .A1(G1976), .A2(G288), .ZN(n801) );
  NOR2_X1 U888 ( .A1(G303), .A2(G1971), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n801), .A2(n793), .ZN(n913) );
  NAND2_X1 U890 ( .A1(n813), .A2(n913), .ZN(n794) );
  XNOR2_X1 U891 ( .A(n794), .B(KEYINPUT104), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G288), .A2(G1976), .ZN(n795) );
  XOR2_X1 U893 ( .A(KEYINPUT105), .B(n795), .Z(n912) );
  INV_X1 U894 ( .A(n912), .ZN(n796) );
  AND2_X1 U895 ( .A1(n797), .A2(n517), .ZN(n798) );
  NOR2_X2 U896 ( .A1(KEYINPUT33), .A2(n798), .ZN(n800) );
  XNOR2_X1 U897 ( .A(n800), .B(n799), .ZN(n806) );
  XOR2_X1 U898 ( .A(G1981), .B(G305), .Z(n906) );
  INV_X1 U899 ( .A(n906), .ZN(n804) );
  NAND2_X1 U900 ( .A1(KEYINPUT33), .A2(n801), .ZN(n802) );
  NOR2_X1 U901 ( .A1(n815), .A2(n802), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT24), .ZN(n809) );
  INV_X1 U905 ( .A(n815), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U907 ( .A(n810), .B(KEYINPUT96), .ZN(n818) );
  NOR2_X1 U908 ( .A1(G303), .A2(G2090), .ZN(n811) );
  XOR2_X1 U909 ( .A(KEYINPUT107), .B(n811), .Z(n812) );
  NAND2_X1 U910 ( .A1(n812), .A2(G8), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n518), .A2(n819), .ZN(n820) );
  XNOR2_X1 U915 ( .A(G1986), .B(G290), .ZN(n911) );
  NAND2_X1 U916 ( .A1(n911), .A2(n834), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n837) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n1004), .ZN(n876) );
  INV_X1 U919 ( .A(n824), .ZN(n827) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n1006), .ZN(n860) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n860), .A2(n825), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n876), .A2(n828), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n1010), .A2(n832), .ZN(n853) );
  NAND2_X1 U928 ( .A1(n833), .A2(n853), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n837), .A2(n836), .ZN(n839) );
  XNOR2_X1 U931 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n838) );
  XNOR2_X1 U932 ( .A(n839), .B(n838), .ZN(G329) );
  NAND2_X1 U933 ( .A1(n840), .A2(G2106), .ZN(n841) );
  XOR2_X1 U934 ( .A(KEYINPUT109), .B(n841), .Z(G217) );
  AND2_X1 U935 ( .A1(G15), .A2(G2), .ZN(n842) );
  NAND2_X1 U936 ( .A1(G661), .A2(n842), .ZN(G259) );
  NAND2_X1 U937 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U938 ( .A1(n844), .A2(n843), .ZN(G188) );
  XOR2_X1 U939 ( .A(G120), .B(KEYINPUT110), .Z(G236) );
  NAND2_X1 U941 ( .A1(n990), .A2(G112), .ZN(n846) );
  NAND2_X1 U942 ( .A1(G136), .A2(n994), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n846), .A2(n845), .ZN(n852) );
  NAND2_X1 U944 ( .A1(G124), .A2(n989), .ZN(n847) );
  XOR2_X1 U945 ( .A(KEYINPUT44), .B(n847), .Z(n848) );
  XNOR2_X1 U946 ( .A(n848), .B(KEYINPUT113), .ZN(n850) );
  NAND2_X1 U947 ( .A1(G100), .A2(n993), .ZN(n849) );
  NAND2_X1 U948 ( .A1(n850), .A2(n849), .ZN(n851) );
  NOR2_X1 U949 ( .A1(n852), .A2(n851), .ZN(G162) );
  INV_X1 U950 ( .A(n853), .ZN(n855) );
  NOR2_X1 U951 ( .A1(n855), .A2(n854), .ZN(n862) );
  XOR2_X1 U952 ( .A(G2084), .B(G160), .Z(n856) );
  NOR2_X1 U953 ( .A1(n1005), .A2(n856), .ZN(n858) );
  NAND2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U955 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n862), .A2(n861), .ZN(n881) );
  XOR2_X1 U957 ( .A(G164), .B(G2078), .Z(n873) );
  NAND2_X1 U958 ( .A1(G127), .A2(n989), .ZN(n864) );
  NAND2_X1 U959 ( .A1(G115), .A2(n990), .ZN(n863) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n865), .B(KEYINPUT47), .ZN(n867) );
  NAND2_X1 U962 ( .A1(G103), .A2(n993), .ZN(n866) );
  NAND2_X1 U963 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n994), .A2(G139), .ZN(n868) );
  XOR2_X1 U965 ( .A(KEYINPUT114), .B(n868), .Z(n869) );
  NOR2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n1013) );
  XNOR2_X1 U967 ( .A(n871), .B(n1013), .ZN(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U969 ( .A(KEYINPUT50), .B(n874), .ZN(n879) );
  XOR2_X1 U970 ( .A(G2090), .B(G162), .Z(n875) );
  NOR2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U972 ( .A(KEYINPUT51), .B(n877), .Z(n878) );
  NAND2_X1 U973 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U974 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U975 ( .A(KEYINPUT52), .B(n882), .ZN(n883) );
  INV_X1 U976 ( .A(KEYINPUT55), .ZN(n956) );
  NAND2_X1 U977 ( .A1(n883), .A2(n956), .ZN(n884) );
  NAND2_X1 U978 ( .A1(n884), .A2(G29), .ZN(n965) );
  XNOR2_X1 U979 ( .A(G2090), .B(G35), .ZN(n899) );
  XOR2_X1 U980 ( .A(G1991), .B(G25), .Z(n885) );
  NAND2_X1 U981 ( .A1(n885), .A2(G28), .ZN(n896) );
  XNOR2_X1 U982 ( .A(G2067), .B(G26), .ZN(n887) );
  XNOR2_X1 U983 ( .A(G2072), .B(G33), .ZN(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(KEYINPUT118), .B(n888), .ZN(n894) );
  XOR2_X1 U986 ( .A(n889), .B(G27), .Z(n892) );
  XOR2_X1 U987 ( .A(n890), .B(G32), .Z(n891) );
  NOR2_X1 U988 ( .A1(n892), .A2(n891), .ZN(n893) );
  NAND2_X1 U989 ( .A1(n894), .A2(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT53), .B(n897), .ZN(n898) );
  NOR2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n902) );
  XOR2_X1 U993 ( .A(G2084), .B(G34), .Z(n900) );
  XNOR2_X1 U994 ( .A(KEYINPUT54), .B(n900), .ZN(n901) );
  NAND2_X1 U995 ( .A1(n902), .A2(n901), .ZN(n957) );
  NOR2_X1 U996 ( .A1(G29), .A2(KEYINPUT55), .ZN(n903) );
  NAND2_X1 U997 ( .A1(n957), .A2(n903), .ZN(n904) );
  NAND2_X1 U998 ( .A1(G11), .A2(n904), .ZN(n963) );
  XNOR2_X1 U999 ( .A(G16), .B(KEYINPUT56), .ZN(n929) );
  XOR2_X1 U1000 ( .A(G168), .B(G1966), .Z(n905) );
  XNOR2_X1 U1001 ( .A(KEYINPUT119), .B(n905), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n908), .B(KEYINPUT57), .ZN(n927) );
  XNOR2_X1 U1004 ( .A(n1018), .B(G1341), .ZN(n925) );
  XOR2_X1 U1005 ( .A(n909), .B(G1956), .Z(n910) );
  NOR2_X1 U1006 ( .A1(n911), .A2(n910), .ZN(n918) );
  AND2_X1 U1007 ( .A1(G303), .A2(G1971), .ZN(n915) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(n916), .B(KEYINPUT120), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n922) );
  XNOR2_X1 U1012 ( .A(G171), .B(G1961), .ZN(n920) );
  XOR2_X1 U1013 ( .A(G1348), .B(n1021), .Z(n919) );
  NAND2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1016 ( .A(KEYINPUT121), .B(n923), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1018 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1019 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1020 ( .A(n930), .B(KEYINPUT122), .ZN(n961) );
  XNOR2_X1 U1021 ( .A(G5), .B(G1961), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(n931), .B(KEYINPUT123), .ZN(n945) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G21), .ZN(n943) );
  XOR2_X1 U1024 ( .A(G1348), .B(KEYINPUT59), .Z(n932) );
  XNOR2_X1 U1025 ( .A(G4), .B(n932), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(G1981), .B(G6), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(G1341), .B(G19), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1029 ( .A(n935), .B(KEYINPUT125), .ZN(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n940) );
  XOR2_X1 U1031 ( .A(G1956), .B(G20), .Z(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT124), .B(n938), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT60), .B(n941), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n952) );
  XNOR2_X1 U1037 ( .A(G1976), .B(G23), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G1971), .B(G22), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G1986), .B(G24), .Z(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(KEYINPUT58), .B(n950), .ZN(n951) );
  NOR2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1044 ( .A(n953), .B(KEYINPUT61), .Z(n954) );
  XNOR2_X1 U1045 ( .A(KEYINPUT126), .B(n954), .ZN(n955) );
  NOR2_X1 U1046 ( .A1(G16), .A2(n955), .ZN(n959) );
  NOR2_X1 U1047 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1048 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1049 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1050 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1052 ( .A(KEYINPUT62), .B(n966), .Z(G311) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1054 ( .A(G108), .ZN(G238) );
  INV_X1 U1055 ( .A(G96), .ZN(G221) );
  INV_X1 U1056 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(n969), .B(KEYINPUT111), .ZN(G261) );
  INV_X1 U1059 ( .A(G261), .ZN(G325) );
  XOR2_X1 U1060 ( .A(G2100), .B(G2096), .Z(n971) );
  XNOR2_X1 U1061 ( .A(G2090), .B(KEYINPUT43), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(n972) );
  XOR2_X1 U1063 ( .A(n972), .B(KEYINPUT42), .Z(n974) );
  XNOR2_X1 U1064 ( .A(G2072), .B(G2678), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n978) );
  XOR2_X1 U1066 ( .A(KEYINPUT112), .B(G2084), .Z(n976) );
  XNOR2_X1 U1067 ( .A(G2067), .B(G2078), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n978), .B(n977), .ZN(G227) );
  XOR2_X1 U1070 ( .A(G1961), .B(G1971), .Z(n980) );
  XNOR2_X1 U1071 ( .A(G1996), .B(G1986), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1073 ( .A(n981), .B(KEYINPUT41), .Z(n983) );
  XNOR2_X1 U1074 ( .A(G1976), .B(G1956), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G2474), .B(G1966), .Z(n985) );
  XNOR2_X1 U1077 ( .A(G1991), .B(G1981), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n985), .B(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(n987), .B(n986), .ZN(G229) );
  INV_X1 U1080 ( .A(n988), .ZN(G319) );
  NAND2_X1 U1081 ( .A1(G130), .A2(n989), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(G118), .A2(n990), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n999) );
  NAND2_X1 U1084 ( .A1(n993), .A2(G106), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n994), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1087 ( .A(n997), .B(KEYINPUT45), .Z(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(KEYINPUT115), .B(n1000), .Z(n1001) );
  XOR2_X1 U1090 ( .A(n1001), .B(KEYINPUT48), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(G164), .B(KEYINPUT46), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1003), .B(n1002), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(n1005), .B(n1004), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1009), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1010), .B(G162), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1012), .B(n1011), .ZN(n1015) );
  XOR2_X1 U1098 ( .A(G160), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1099 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(G37), .A2(n1016), .ZN(G395) );
  XNOR2_X1 U1101 ( .A(n1018), .B(n1017), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G286), .B(G301), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(n1020), .B(n1019), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NOR2_X1 U1105 ( .A1(G37), .A2(n1023), .ZN(G397) );
  NOR2_X1 U1106 ( .A1(G227), .A2(G229), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT116), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT49), .B(n1025), .ZN(n1030) );
  NOR2_X1 U1109 ( .A1(G395), .A2(G397), .ZN(n1026) );
  XOR2_X1 U1110 ( .A(KEYINPUT117), .B(n1026), .Z(n1027) );
  NAND2_X1 U1111 ( .A1(G319), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1112 ( .A1(G401), .A2(n1028), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(G225) );
  INV_X1 U1114 ( .A(G225), .ZN(G308) );
endmodule

