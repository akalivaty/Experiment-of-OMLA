//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G116), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G116), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(KEYINPUT67), .A3(G119), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT2), .A2(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT2), .A2(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT2), .A3(G113), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n194), .A2(new_n200), .A3(KEYINPUT68), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n194), .B2(new_n200), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(new_n211), .B2(G101), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n206), .A2(new_n209), .A3(new_n217), .A4(new_n210), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n216), .A2(KEYINPUT77), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT77), .B1(new_n216), .B2(new_n218), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n204), .B(new_n214), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n194), .A2(new_n200), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n194), .A2(new_n200), .A3(KEYINPUT68), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n205), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n208), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n218), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(new_n189), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n232), .B(G113), .C1(KEYINPUT5), .C2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n221), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT6), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n221), .A2(KEYINPUT79), .A3(new_n235), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(new_n239), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G125), .ZN(new_n244));
  INV_X1    g058(.A(G128), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n247), .B2(KEYINPUT1), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n246), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n246), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n248), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n250), .A2(new_n252), .A3(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n247), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n244), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n247), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n255), .B1(new_n253), .B2(new_n246), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n262), .B1(new_n244), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G224), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n221), .A2(KEYINPUT79), .A3(new_n235), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT79), .B1(new_n221), .B2(new_n235), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n274), .A2(new_n275), .A3(new_n241), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n221), .A2(new_n235), .A3(new_n241), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT6), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n243), .B(new_n273), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G210), .B1(G237), .B2(G902), .ZN(new_n280));
  XOR2_X1   g094(.A(new_n241), .B(KEYINPUT8), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n226), .A2(new_n234), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n230), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n235), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n272), .A2(KEYINPUT7), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT80), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n270), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n285), .A2(KEYINPUT80), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n270), .A2(new_n287), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n284), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G902), .B1(new_n292), .B2(new_n277), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n279), .A2(new_n280), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n280), .B1(new_n279), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G237), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(new_n271), .A3(G143), .A4(G214), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n298), .A2(KEYINPUT82), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(KEYINPUT82), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT64), .B(G143), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(new_n271), .A3(G214), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n303), .B1(new_n302), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n301), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT17), .A3(G131), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n244), .A2(G140), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(KEYINPUT74), .A3(G125), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n311), .A2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n316), .A2(new_n246), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n246), .B1(new_n316), .B2(new_n318), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n308), .A2(G131), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n302), .A2(new_n304), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT81), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n326), .A2(new_n305), .B1(new_n300), .B2(new_n299), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n308), .A2(KEYINPUT18), .A3(G131), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT18), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n311), .A2(new_n312), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n246), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n314), .A2(G146), .A3(new_n315), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n327), .A2(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n323), .A2(new_n331), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G113), .B(G122), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(new_n205), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT83), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n332), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n324), .A2(new_n329), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n316), .A2(new_n318), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G146), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n335), .A2(KEYINPUT19), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n314), .A2(new_n315), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(KEYINPUT19), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n346), .B1(new_n349), .B2(G146), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n343), .B1(new_n344), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n341), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n339), .A2(new_n342), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(G475), .A2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT20), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n352), .ZN(new_n357));
  INV_X1    g171(.A(new_n331), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n343), .B(new_n342), .C1(new_n358), .C2(new_n322), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n354), .ZN(new_n362));
  INV_X1    g176(.A(G902), .ZN(new_n363));
  INV_X1    g177(.A(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n323), .A2(new_n331), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n341), .B1(new_n365), .B2(new_n343), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n363), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n356), .A2(new_n362), .B1(new_n367), .B2(G475), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n250), .A2(new_n252), .A3(G128), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n245), .A2(G143), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(G134), .ZN(new_n372));
  INV_X1    g186(.A(G134), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n369), .B2(new_n370), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G122), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G116), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n208), .B1(new_n377), .B2(KEYINPUT14), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n188), .A2(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n378), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT86), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n372), .A2(new_n374), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n384), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n370), .B1(new_n369), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n369), .A2(new_n387), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT85), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n369), .A2(KEYINPUT85), .A3(new_n387), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(new_n373), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n380), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n397), .A3(new_n208), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n399), .B(new_n400), .C1(G134), .C2(new_n371), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n383), .A2(new_n386), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT9), .B(G234), .ZN(new_n403));
  INV_X1    g217(.A(G217), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n403), .A2(new_n404), .A3(G953), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n405), .ZN(new_n407));
  OAI221_X1 g221(.A(new_n407), .B1(new_n394), .B2(new_n401), .C1(new_n383), .C2(new_n386), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n363), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n409), .B(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI211_X1 g227(.A(new_n363), .B(new_n271), .C1(G234), .C2(G237), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(KEYINPUT87), .A2(G952), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT87), .A2(G952), .ZN(new_n418));
  AOI21_X1  g232(.A(G953), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n297), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n368), .A2(new_n413), .A3(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n296), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G472), .A2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT32), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n256), .B1(new_n302), .B2(G146), .ZN(new_n430));
  INV_X1    g244(.A(new_n247), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n302), .B2(G146), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n430), .A2(new_n267), .B1(new_n432), .B2(new_n263), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n434));
  INV_X1    g248(.A(G137), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(KEYINPUT11), .A2(G134), .ZN(new_n437));
  NAND2_X1  g251(.A1(KEYINPUT65), .A2(G137), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT11), .A2(G134), .ZN(new_n440));
  NOR2_X1   g254(.A1(KEYINPUT11), .A2(G134), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(G137), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n439), .A2(new_n442), .A3(new_n328), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n436), .A2(new_n373), .A3(new_n438), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n328), .B1(G134), .B2(G137), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n445), .B(new_n450), .C1(new_n257), .C2(new_n261), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n447), .A2(new_n451), .B1(new_n226), .B2(new_n201), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n445), .A2(new_n450), .ZN(new_n453));
  INV_X1    g267(.A(new_n248), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n430), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(new_n260), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n439), .A2(new_n328), .A3(new_n442), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n328), .B1(new_n439), .B2(new_n442), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT69), .B1(new_n459), .B2(new_n269), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n433), .A2(new_n446), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n456), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n204), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n452), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT70), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n204), .B(new_n456), .C1(new_n460), .C2(new_n462), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n468), .B(KEYINPUT28), .C1(new_n469), .C2(new_n452), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n447), .A3(new_n451), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G210), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(G237), .A3(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT27), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G101), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n460), .A2(new_n462), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n480), .B1(new_n481), .B2(new_n451), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n447), .A2(new_n451), .A3(new_n480), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n204), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n469), .ZN(new_n486));
  INV_X1    g300(.A(new_n478), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT31), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n483), .B1(new_n463), .B2(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n469), .B1(new_n490), .B2(new_n204), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n429), .B1(new_n479), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n478), .B1(new_n471), .B2(new_n466), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n496), .A2(KEYINPUT29), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n463), .A2(new_n464), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT28), .B1(new_n498), .B2(new_n469), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n467), .A2(new_n470), .A3(new_n496), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT29), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n491), .B2(new_n487), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n500), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G472), .ZN(new_n505));
  AND4_X1   g319(.A1(new_n492), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n492), .B1(new_n491), .B2(new_n487), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n473), .A2(new_n478), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n427), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n495), .B(new_n505), .C1(new_n510), .C2(KEYINPUT32), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n403), .B2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G140), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n271), .A2(G227), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT78), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n258), .A2(new_n247), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT1), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n253), .B2(new_n246), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(new_n245), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n230), .B1(new_n520), .B2(new_n260), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n521), .B2(KEYINPUT10), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT1), .B1(new_n302), .B2(G146), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n523), .A2(G128), .B1(new_n247), .B2(new_n258), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n231), .B1(new_n524), .B2(new_n261), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT10), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT78), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n218), .A2(new_n229), .A3(KEYINPUT10), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n455), .B2(new_n260), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT77), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n216), .A2(KEYINPUT77), .A3(new_n218), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n269), .A2(new_n213), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n528), .A2(new_n459), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n459), .B1(new_n528), .B2(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n515), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n528), .A2(new_n459), .A3(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(new_n515), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n455), .A2(new_n230), .A3(new_n260), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n446), .B1(new_n521), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(KEYINPUT12), .B(new_n446), .C1(new_n521), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n541), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  AOI211_X1 g363(.A(G469), .B(G902), .C1(new_n540), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n541), .A2(new_n548), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n515), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n521), .A2(new_n516), .A3(KEYINPUT10), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT78), .B1(new_n525), .B2(new_n526), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n537), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n446), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n541), .A3(new_n542), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(new_n557), .A3(G469), .ZN(new_n558));
  NAND2_X1  g372(.A1(G469), .A2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n512), .B1(new_n550), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n245), .A2(G119), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n191), .B2(G128), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n245), .A2(KEYINPUT71), .A3(G119), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n191), .A2(G128), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT72), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n562), .A2(new_n569), .A3(new_n570), .A4(KEYINPUT23), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT72), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n572), .A2(new_n574), .A3(G119), .A4(new_n245), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n568), .B1(new_n576), .B2(G110), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(new_n346), .A3(new_n336), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n575), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n575), .A3(KEYINPUT73), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(G110), .A3(new_n582), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n566), .A2(new_n567), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n578), .B1(new_n585), .B2(new_n321), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT75), .B(new_n578), .C1(new_n585), .C2(new_n321), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n587), .A3(new_n592), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n404), .B1(G234), .B2(new_n363), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT76), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(KEYINPUT76), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n594), .B2(new_n595), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n597), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g419(.A(KEYINPUT25), .B(G902), .C1(new_n594), .C2(new_n595), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n601), .B(new_n602), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n561), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n425), .A2(new_n511), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  OAI21_X1  g424(.A(new_n363), .B1(new_n479), .B2(new_n494), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n509), .A2(new_n489), .A3(new_n493), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n611), .A2(G472), .B1(new_n426), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n406), .A2(new_n615), .A3(new_n408), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT88), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n406), .A2(KEYINPUT88), .A3(new_n408), .A4(new_n615), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n407), .A2(KEYINPUT89), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n615), .B1(new_n402), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n402), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n410), .A2(G902), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n618), .A2(new_n619), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n409), .A2(new_n410), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n361), .B1(new_n360), .B2(new_n354), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT20), .B(new_n355), .C1(new_n357), .C2(new_n359), .ZN(new_n628));
  INV_X1    g442(.A(G475), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n343), .B1(new_n358), .B2(new_n322), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n352), .ZN(new_n631));
  AOI21_X1  g445(.A(G902), .B1(new_n631), .B2(new_n359), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n614), .A2(new_n296), .A3(new_n422), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT34), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  XNOR2_X1  g451(.A(new_n422), .B(KEYINPUT90), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n187), .B(new_n638), .C1(new_n294), .C2(new_n295), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n413), .A2(new_n633), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n614), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(G469), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n542), .B1(new_n556), .B2(new_n541), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n541), .A2(new_n542), .A3(new_n548), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n646), .B(new_n363), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n559), .A3(new_n558), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n593), .A2(KEYINPUT36), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n586), .A2(KEYINPUT91), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n598), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n605), .B2(new_n606), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n650), .A2(new_n657), .A3(new_n512), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n425), .A2(new_n613), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT92), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  NAND2_X1  g476(.A1(new_n612), .A2(new_n426), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n428), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n612), .A2(new_n429), .B1(new_n504), .B2(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n296), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n658), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n368), .A2(new_n412), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n414), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(new_n421), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n279), .A2(new_n293), .ZN(new_n675));
  INV_X1    g489(.A(new_n280), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n279), .A2(new_n280), .A3(new_n293), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n657), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n368), .A2(new_n413), .ZN(new_n683));
  AND4_X1   g497(.A1(new_n187), .A2(new_n681), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n671), .B(KEYINPUT39), .Z(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n561), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT40), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n498), .A2(new_n469), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n478), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n478), .B2(new_n491), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n612), .A2(new_n429), .B1(G472), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n664), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(KEYINPUT94), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n684), .B(new_n688), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n253), .ZN(G45));
  INV_X1    g511(.A(new_n671), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n626), .A2(new_n633), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n667), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  INV_X1    g516(.A(new_n607), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n363), .B1(new_n647), .B2(new_n648), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n512), .A3(new_n649), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT95), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(KEYINPUT95), .A3(new_n512), .A4(new_n649), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n511), .A2(new_n703), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n634), .ZN(new_n711));
  INV_X1    g525(.A(new_n187), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n677), .B2(new_n678), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n713), .A3(new_n423), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT96), .B1(new_n710), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n708), .A2(new_n709), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n607), .B1(new_n664), .B2(new_n665), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT96), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n296), .A2(new_n634), .A3(new_n422), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT41), .B(G113), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n722), .B(new_n724), .ZN(G15));
  NOR2_X1   g539(.A1(new_n710), .A2(new_n642), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n188), .ZN(G18));
  NAND4_X1  g541(.A1(new_n657), .A2(new_n368), .A3(new_n413), .A4(new_n423), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n664), .B2(new_n665), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n705), .A2(new_n512), .A3(new_n649), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT98), .B1(new_n713), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT98), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n296), .A2(new_n706), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n729), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT99), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n729), .B(KEYINPUT99), .C1(new_n731), .C2(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  NAND2_X1  g553(.A1(new_n499), .A2(new_n472), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n478), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n489), .A3(new_n493), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n426), .ZN(new_n743));
  INV_X1    g557(.A(G472), .ZN(new_n744));
  AOI21_X1  g558(.A(G902), .B1(new_n508), .B2(new_n509), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n703), .B(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n427), .B1(new_n508), .B2(new_n741), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(G472), .B2(new_n611), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(KEYINPUT100), .A3(new_n703), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT101), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n713), .A2(new_n683), .ZN(new_n754));
  INV_X1    g568(.A(new_n638), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n716), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n753), .B1(new_n752), .B2(new_n756), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n376), .ZN(G24));
  NOR2_X1   g574(.A1(new_n745), .A2(new_n744), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n761), .A2(new_n682), .A3(new_n749), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n700), .C1(new_n731), .C2(new_n733), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  NOR3_X1   g578(.A1(new_n294), .A2(new_n295), .A3(new_n712), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n511), .A2(new_n608), .A3(new_n700), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n677), .A2(new_n187), .A3(new_n678), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n664), .B2(new_n665), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n770), .A2(KEYINPUT42), .A3(new_n608), .A4(new_n700), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n768), .A2(KEYINPUT102), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT102), .B1(new_n768), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NAND4_X1  g589(.A1(new_n511), .A2(new_n608), .A3(new_n672), .A4(new_n765), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G134), .ZN(G36));
  NAND2_X1  g591(.A1(new_n552), .A2(new_n557), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n646), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n779), .B2(new_n778), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n559), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n550), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n559), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n512), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n686), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n626), .A2(new_n368), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT43), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n790), .B(new_n657), .C1(new_n510), .C2(new_n761), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT44), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n769), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n787), .B(new_n793), .C1(new_n792), .C2(new_n791), .ZN(new_n794));
  XOR2_X1   g608(.A(KEYINPUT103), .B(G137), .Z(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT104), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n794), .B(new_n796), .ZN(G39));
  XNOR2_X1  g611(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n786), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(new_n512), .A3(new_n798), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n511), .A2(new_n703), .A3(new_n699), .A4(new_n769), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT106), .B(G140), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G42));
  INV_X1    g619(.A(new_n421), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n752), .A2(new_n806), .A3(new_n790), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n681), .A2(new_n187), .A3(new_n706), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n769), .A2(new_n706), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT112), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n813), .A2(new_n806), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n814), .A2(new_n815), .A3(new_n790), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n815), .B1(new_n814), .B2(new_n790), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n762), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n800), .A2(new_n801), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n705), .A2(new_n649), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n512), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n765), .B(new_n807), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n811), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n694), .A2(new_n695), .A3(new_n607), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n626), .A2(new_n633), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT114), .B1(new_n827), .B2(new_n828), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(KEYINPUT51), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(new_n831), .A3(KEYINPUT115), .A4(KEYINPUT51), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  INV_X1    g651(.A(new_n831), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n837), .B1(new_n838), .B2(new_n823), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n807), .B1(new_n731), .B2(new_n733), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n419), .C1(new_n826), .C2(new_n634), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n718), .B1(new_n816), .B2(new_n817), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(KEYINPUT48), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n726), .B1(new_n715), .B2(new_n721), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n738), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n759), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n608), .A2(new_n640), .A3(new_n613), .A4(new_n711), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n850), .A2(new_n609), .A3(new_n659), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n495), .A2(new_n505), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT32), .B1(new_n612), .B2(new_n426), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n765), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n633), .A2(new_n412), .A3(new_n671), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n658), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT108), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n368), .A2(new_n413), .A3(new_n698), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n561), .A3(new_n682), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT108), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n770), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n769), .A2(new_n561), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n750), .A3(new_n657), .A4(new_n700), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n776), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT107), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n639), .B2(new_n668), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n713), .A2(KEYINPUT107), .A3(new_n641), .A4(new_n638), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n608), .A4(new_n613), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n851), .A2(new_n862), .A3(new_n865), .A4(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n773), .A3(new_n772), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT109), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n849), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n773), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n869), .A2(new_n609), .A3(new_n659), .A4(new_n850), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n776), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n861), .B2(new_n857), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n768), .A2(KEYINPUT102), .A3(new_n771), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n874), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n847), .B(new_n738), .C1(new_n757), .C2(new_n758), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT109), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n666), .B(new_n658), .C1(new_n672), .C2(new_n700), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n561), .A2(new_n657), .A3(new_n671), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(new_n693), .A3(new_n713), .A4(new_n683), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n763), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(KEYINPUT52), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n763), .A2(new_n883), .A3(new_n888), .A4(new_n885), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n873), .A2(new_n882), .A3(KEYINPUT53), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT110), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n847), .A2(new_n738), .ZN(new_n894));
  INV_X1    g708(.A(new_n758), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n752), .A2(new_n756), .A3(new_n753), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n862), .A2(new_n865), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n875), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n894), .A2(new_n897), .A3(new_n774), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n890), .B1(new_n900), .B2(KEYINPUT109), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT110), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT53), .A4(new_n873), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n873), .A2(new_n891), .A3(new_n882), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT111), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n768), .B2(new_n771), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n899), .A2(new_n887), .A3(new_n889), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n909), .B1(new_n911), .B2(new_n881), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n876), .A2(new_n878), .A3(new_n910), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n849), .A2(new_n891), .A3(KEYINPUT111), .A4(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n904), .A2(new_n905), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n846), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n626), .A2(new_n368), .A3(new_n187), .A4(new_n512), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n681), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n825), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n271), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n901), .B2(new_n873), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n912), .A2(new_n914), .ZN(new_n929));
  OAI211_X1 g743(.A(G210), .B(G902), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n276), .A2(new_n278), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n239), .B2(new_n276), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n273), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n936), .A2(KEYINPUT56), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n927), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n930), .B2(KEYINPUT117), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(KEYINPUT117), .B2(new_n930), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n940), .B2(new_n936), .ZN(G51));
  XOR2_X1   g755(.A(new_n559), .B(KEYINPUT57), .Z(new_n942));
  OAI21_X1  g756(.A(KEYINPUT54), .B1(new_n928), .B2(new_n929), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT118), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n912), .A2(new_n914), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n906), .A2(new_n944), .A3(new_n916), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n944), .B1(new_n915), .B2(new_n916), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n942), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n540), .A2(new_n549), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n915), .A2(new_n363), .A3(new_n781), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n926), .B1(new_n951), .B2(new_n952), .ZN(G54));
  INV_X1    g767(.A(new_n915), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n353), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n927), .B1(new_n955), .B2(new_n353), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n955), .B2(new_n353), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G60));
  AND3_X1   g774(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n961));
  NAND2_X1  g775(.A1(G478), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT59), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n961), .B(new_n963), .C1(new_n947), .C2(new_n948), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n927), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n961), .B1(new_n918), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G63));
  OR2_X1    g781(.A1(new_n654), .A2(new_n655), .ZN(new_n968));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT121), .Z(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  OAI211_X1 g785(.A(new_n968), .B(new_n971), .C1(new_n928), .C2(new_n929), .ZN(new_n972));
  INV_X1    g786(.A(new_n971), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n915), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n927), .B(new_n972), .C1(new_n974), .C2(new_n596), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT120), .ZN(new_n976));
  XNOR2_X1  g790(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n977), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(G66));
  INV_X1    g795(.A(new_n415), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n271), .B1(new_n982), .B2(G224), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n849), .A2(new_n876), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n271), .ZN(new_n985));
  INV_X1    g799(.A(G898), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n933), .B1(new_n986), .B2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n985), .B(new_n987), .ZN(G69));
  AND2_X1   g802(.A1(new_n794), .A2(new_n803), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n763), .A2(new_n883), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n696), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n770), .A2(new_n608), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n686), .B1(new_n634), .B2(new_n668), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n991), .A2(KEYINPUT62), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n989), .B(new_n994), .C1(KEYINPUT62), .C2(new_n991), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(new_n271), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n490), .B(new_n349), .Z(new_n997));
  OR2_X1    g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n271), .A2(G900), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n787), .A2(new_n713), .A3(new_n683), .A4(new_n718), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n990), .A2(new_n776), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n989), .A2(new_n774), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n999), .B1(new_n1002), .B2(new_n271), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n997), .B1(new_n1003), .B2(KEYINPUT123), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(KEYINPUT123), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n998), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n271), .B1(G227), .B2(G900), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(KEYINPUT124), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1007), .A2(KEYINPUT124), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1003), .A2(KEYINPUT123), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1003), .A2(KEYINPUT123), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1011), .A2(new_n997), .A3(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1013), .A2(KEYINPUT124), .A3(new_n1007), .A4(new_n998), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1010), .A2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT125), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1018), .B1(new_n1002), .B2(new_n984), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n491), .A2(new_n478), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n926), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1018), .B1(new_n995), .B2(new_n984), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n491), .A2(new_n478), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1017), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n907), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1029), .A2(KEYINPUT126), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT126), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1025), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(G57));
endmodule


