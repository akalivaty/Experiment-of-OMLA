//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n625, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT69), .B(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n463), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n470), .A2(new_n471), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  INV_X1    g054(.A(new_n463), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n475), .A2(new_n481), .ZN(G160));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n478), .B(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n489), .B2(G136), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n486), .A2(new_n480), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n491), .A2(new_n492), .A3(G124), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n491), .B2(G124), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(new_n490), .C1(new_n493), .C2(new_n494), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n497), .A2(new_n500), .ZN(G162));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n502), .B(G2104), .C1(G114), .C2(new_n487), .ZN(new_n503));
  OAI211_X1 g078(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  AND3_X1   g083(.A1(new_n506), .A2(new_n508), .A3(G138), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n509), .A2(new_n510), .A3(new_n467), .A4(new_n472), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(new_n508), .A3(G138), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n465), .A2(new_n466), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT4), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n511), .B2(new_n514), .ZN(G164));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT74), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G62), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n522), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n531), .A2(G88), .B1(G50), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(G166));
  AND2_X1   g110(.A1(new_n531), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n522), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n537), .B(new_n539), .C1(new_n540), .C2(new_n532), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n530), .A2(new_n545), .B1(new_n532), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n531), .A2(G81), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n533), .A2(G43), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n516), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n549), .A2(new_n550), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT76), .B1(new_n557), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT79), .B1(new_n530), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n522), .A2(new_n529), .A3(new_n569), .A4(G91), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n571), .B(KEYINPUT9), .C1(new_n532), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n529), .A2(G53), .A3(G543), .A4(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n568), .A2(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n520), .A2(KEYINPUT81), .A3(new_n521), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G78), .A2(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT80), .Z(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n584), .ZN(G299));
  INV_X1    g160(.A(G171), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  NAND3_X1  g162(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(G303));
  AOI22_X1  g163(.A1(new_n531), .A2(G87), .B1(G49), .B2(new_n533), .ZN(new_n589));
  INV_X1    g164(.A(new_n522), .ZN(new_n590));
  INV_X1    g165(.A(G74), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n516), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(new_n594), .B2(new_n595), .ZN(G288));
  AOI22_X1  g171(.A1(new_n522), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n597), .A2(new_n516), .B1(new_n532), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n522), .A2(G86), .A3(new_n529), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(G305));
  AND2_X1   g176(.A1(new_n522), .A2(G60), .ZN(new_n602));
  AND2_X1   g177(.A1(G72), .A2(G543), .ZN(new_n603));
  OAI21_X1  g178(.A(G651), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT83), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n531), .A2(G85), .B1(G47), .B2(new_n533), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n604), .A2(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT85), .B(G66), .Z(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n579), .B2(new_n580), .ZN(new_n613));
  AND2_X1   g188(.A1(G79), .A2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G54), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n532), .B2(KEYINPUT84), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(KEYINPUT84), .B2(new_n532), .ZN(new_n618));
  AOI21_X1  g193(.A(KEYINPUT10), .B1(new_n531), .B2(G92), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n615), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT86), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n611), .B1(new_n622), .B2(new_n610), .ZN(G284));
  AOI21_X1  g198(.A(new_n611), .B1(new_n622), .B2(new_n610), .ZN(G321));
  NAND2_X1  g199(.A1(G299), .A2(new_n610), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g201(.A(new_n625), .B1(new_n610), .B2(G168), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n622), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n559), .A2(new_n610), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n628), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g209(.A1(new_n467), .A2(new_n472), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(new_n476), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT87), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n489), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n491), .A2(G123), .ZN(new_n643));
  OAI221_X1 g218(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n463), .C2(G111), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2096), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n639), .B2(new_n638), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT88), .Z(G156));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n655), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(G401));
  INV_X1    g240(.A(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT17), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n639), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(KEYINPUT18), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n682), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  MUX2_X1   g263(.A(new_n688), .B(new_n687), .S(new_n680), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n698), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  NOR2_X1   g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT89), .Z(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n486), .A2(new_n480), .ZN(new_n706));
  INV_X1    g281(.A(G119), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n705), .B1(new_n706), .B2(new_n707), .C1(new_n708), .C2(new_n488), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G25), .B2(G29), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G24), .ZN(new_n720));
  INV_X1    g295(.A(G290), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  INV_X1    g297(.A(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n716), .B2(new_n717), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G6), .B(G305), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT92), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT32), .B(G1981), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n719), .A2(G22), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G166), .B2(new_n719), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(G1971), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G23), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT93), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G288), .B2(new_n719), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT33), .B(G1976), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n734), .A2(G1971), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n731), .A2(new_n735), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n726), .B1(new_n742), .B2(KEYINPUT34), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT36), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n742), .A2(KEYINPUT34), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n726), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT100), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  INV_X1    g329(.A(G139), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n754), .B1(new_n488), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT96), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n635), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(new_n463), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n757), .A2(KEYINPUT97), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT97), .B1(new_n757), .B2(new_n759), .ZN(new_n761));
  OAI21_X1  g336(.A(KEYINPUT98), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(new_n759), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n757), .A2(KEYINPUT97), .A3(new_n759), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n752), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n752), .A2(G33), .ZN(new_n770));
  OR3_X1    g345(.A1(new_n769), .A2(KEYINPUT99), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(KEYINPUT99), .B1(new_n769), .B2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n751), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n771), .A2(KEYINPUT100), .A3(G2072), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n752), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n489), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n491), .A2(G129), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(G105), .B2(new_n476), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n779), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n778), .B1(new_n787), .B2(new_n752), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT101), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n719), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n719), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1966), .ZN(new_n795));
  INV_X1    g370(.A(G34), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(KEYINPUT24), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n752), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G160), .B2(new_n752), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n795), .B1(G2084), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G2084), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n719), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n560), .B2(new_n719), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n719), .A2(G20), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT23), .Z(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G299), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1956), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR4_X1   g385(.A1(new_n792), .A2(new_n802), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G171), .A2(new_n719), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G5), .B2(new_n719), .ZN(new_n813));
  INV_X1    g388(.A(G1961), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  NAND2_X1  g391(.A1(G164), .A2(G29), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G27), .B2(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n815), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n816), .B2(new_n818), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT31), .B(G11), .Z(new_n821));
  INV_X1    g396(.A(G28), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT30), .ZN(new_n823));
  AOI21_X1  g398(.A(G29), .B1(new_n822), .B2(KEYINPUT30), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n825), .B1(new_n752), .B2(new_n645), .C1(new_n813), .C2(new_n814), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n788), .B2(new_n790), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n752), .A2(G26), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT28), .Z(new_n829));
  NOR2_X1   g404(.A1(G104), .A2(G2105), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT95), .Z(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n832));
  INV_X1    g407(.A(G128), .ZN(new_n833));
  INV_X1    g408(.A(G140), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n832), .B1(new_n706), .B2(new_n833), .C1(new_n834), .C2(new_n488), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(G29), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2067), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n820), .A2(new_n827), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G1348), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n622), .A2(new_n719), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G4), .B2(new_n719), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(G29), .A2(G35), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G162), .B2(G29), .ZN(new_n844));
  XNOR2_X1  g419(.A(KEYINPUT29), .B(G2090), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n841), .A2(new_n839), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n811), .A2(new_n842), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n774), .B2(new_n773), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n750), .A2(new_n777), .A3(new_n850), .ZN(G311));
  NAND3_X1  g426(.A1(new_n750), .A2(new_n777), .A3(new_n850), .ZN(G150));
  AOI22_X1  g427(.A1(new_n531), .A2(G93), .B1(G55), .B2(new_n533), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n516), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n559), .A2(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n855), .A2(new_n554), .A3(new_n557), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n621), .B(KEYINPUT86), .Z(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n628), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n859), .B(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n863), .A2(new_n864), .A3(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n855), .A2(G860), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  OR2_X1    g443(.A1(new_n835), .A2(G164), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n835), .A2(G164), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n786), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n787), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n762), .A2(new_n768), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n760), .C2(new_n761), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n711), .A2(new_n637), .A3(new_n712), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n637), .B1(new_n711), .B2(new_n712), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n489), .A2(new_n880), .A3(G142), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n489), .B2(G142), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI221_X1 g458(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n463), .C2(G118), .ZN(new_n884));
  INV_X1    g459(.A(G130), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n706), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n878), .A2(new_n879), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n877), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n876), .A3(new_n875), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n497), .A2(new_n500), .B1(new_n475), .B2(new_n481), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT102), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n496), .A2(G160), .A3(new_n499), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n645), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n900), .ZN(new_n902));
  INV_X1    g477(.A(new_n645), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n903), .A3(new_n898), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n894), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n891), .A3(new_n893), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n906), .B2(new_n908), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(G395));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n632), .A2(new_n858), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n621), .B(G299), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n631), .A2(new_n856), .A3(new_n857), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n914), .A2(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(G299), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n621), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n915), .A2(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n913), .B(new_n917), .C1(new_n918), .C2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n924), .B1(new_n914), .B2(new_n916), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G290), .B(G288), .ZN(new_n930));
  XNOR2_X1  g505(.A(G166), .B(G305), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n928), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(G868), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT105), .B1(new_n855), .B2(new_n610), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n933), .A2(KEYINPUT105), .A3(G868), .A4(new_n935), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  AND2_X1   g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  XNOR2_X1  g517(.A(G168), .B(G171), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n858), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n856), .A2(new_n857), .A3(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n920), .ZN(new_n948));
  INV_X1    g523(.A(new_n924), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n947), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n942), .B1(new_n950), .B2(new_n932), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n915), .B1(new_n945), .B2(new_n946), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n945), .A2(new_n946), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n924), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n934), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT106), .B(KEYINPUT43), .C1(new_n951), .C2(new_n955), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n960), .B2(new_n923), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n948), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n932), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n954), .B2(new_n934), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n958), .A2(new_n959), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n965), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n950), .A2(new_n932), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT43), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT44), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(G397));
  XOR2_X1   g550(.A(new_n835), .B(G2067), .Z(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT110), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n787), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n512), .A2(KEYINPUT4), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n478), .A2(new_n463), .A3(G138), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n635), .A2(new_n982), .B1(new_n983), .B2(KEYINPUT4), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n984), .B2(new_n505), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n473), .A2(new_n474), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n480), .ZN(new_n989));
  INV_X1    g564(.A(new_n481), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(G40), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n978), .A2(new_n980), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n979), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(new_n786), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT109), .Z(new_n996));
  AND2_X1   g571(.A1(new_n714), .A2(new_n717), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n714), .A2(new_n717), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n992), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n721), .A2(new_n723), .A3(new_n992), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT48), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n993), .A2(new_n996), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n978), .A2(new_n992), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n994), .B(KEYINPUT46), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n835), .A2(G2067), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1008), .B1(new_n992), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n1013));
  INV_X1    g588(.A(new_n505), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n467), .A2(new_n472), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n463), .A2(new_n510), .A3(G138), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n510), .B1(new_n509), .B2(new_n478), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1013), .B1(new_n1019), .B2(new_n981), .ZN(new_n1020));
  NOR3_X1   g595(.A1(G164), .A2(KEYINPUT111), .A3(G1384), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n986), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G164), .A2(G1384), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n991), .B1(KEYINPUT45), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1966), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1013), .A3(new_n981), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT111), .B1(G164), .B2(G1384), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n991), .B1(KEYINPUT50), .B2(new_n985), .ZN(new_n1030));
  INV_X1    g605(.A(G2084), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(G8), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(G168), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT51), .B1(new_n1036), .B2(KEYINPUT121), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1019), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1041));
  INV_X1    g616(.A(G40), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n475), .A2(new_n1042), .A3(new_n481), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n986), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1040), .B1(new_n1046), .B2(G1966), .ZN(new_n1047));
  OAI211_X1 g622(.A(G8), .B(new_n1037), .C1(new_n1047), .C2(G286), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1035), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT62), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT126), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1050), .A2(KEYINPUT62), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1026), .A2(new_n1027), .A3(new_n1043), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1055), .A2(new_n1056), .A3(G8), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1055), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  OR2_X1    g635(.A1(G288), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G303), .A2(G8), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1971), .ZN(new_n1067));
  INV_X1    g642(.A(new_n987), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(new_n1044), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(G2090), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1066), .A2(new_n1071), .A3(G8), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT113), .B(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1061), .B(new_n1074), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1075));
  INV_X1    g650(.A(G1981), .ZN(new_n1076));
  INV_X1    g651(.A(new_n599), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT114), .B(G86), .Z(new_n1078));
  NAND2_X1  g653(.A1(new_n531), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n599), .A2(G1981), .A3(new_n600), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT115), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1084), .A2(new_n1085), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1063), .A2(new_n1072), .A3(new_n1075), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT50), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1088));
  INV_X1    g663(.A(G2090), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n991), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1069), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1034), .B1(new_n1092), .B2(KEYINPUT116), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1069), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1066), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n987), .A2(new_n816), .A3(new_n1043), .A4(new_n1041), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1070), .A2(new_n814), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1022), .A2(KEYINPUT122), .A3(new_n816), .A4(new_n1024), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT53), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT122), .B1(new_n1046), .B2(new_n816), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1087), .A2(new_n1096), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1050), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1053), .A2(new_n1054), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1047), .A2(G8), .A3(G168), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1087), .A2(new_n1096), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1066), .B1(new_n1071), .B2(G8), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1110), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1109), .A2(KEYINPUT63), .B1(new_n1087), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1059), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1086), .ZN(new_n1115));
  OR2_X1    g690(.A1(G288), .A2(G1976), .ZN(new_n1116));
  OAI22_X1  g691(.A1(new_n1115), .A2(new_n1116), .B1(G1981), .B2(G305), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1063), .A2(new_n1075), .A3(new_n1086), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1072), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1114), .A2(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1107), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1087), .A2(new_n1096), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(new_n1050), .ZN(new_n1123));
  OAI211_X1 g698(.A(G301), .B(new_n1099), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1070), .A2(new_n814), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n991), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1043), .A2(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1098), .A2(G2078), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n987), .A3(new_n1041), .A4(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1126), .A2(new_n1127), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1125), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT124), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1124), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1103), .A2(G171), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1134), .A2(G171), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1125), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1123), .A2(KEYINPUT125), .A3(new_n1140), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1055), .A2(G2067), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1070), .A2(new_n839), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT118), .B1(new_n1055), .B2(G2067), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(KEYINPUT60), .A4(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n860), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1146), .A2(new_n1145), .B1(new_n1070), .B2(new_n839), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1152), .A2(KEYINPUT60), .A3(new_n622), .A4(new_n1149), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1151), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1028), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1043), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n809), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT57), .ZN(new_n1162));
  AOI211_X1 g737(.A(KEYINPUT117), .B(new_n1162), .C1(new_n576), .C2(new_n584), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(KEYINPUT117), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT117), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT57), .ZN(new_n1166));
  AND4_X1   g741(.A1(new_n584), .A2(new_n576), .A3(new_n1164), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(KEYINPUT56), .B(G2072), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1024), .A2(new_n987), .A3(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1161), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1158), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(KEYINPUT58), .B(G1341), .Z(new_n1174));
  NAND2_X1  g749(.A1(new_n1055), .A2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(KEYINPUT120), .B(G1996), .Z(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n987), .A2(new_n1043), .A3(new_n1041), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n559), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT59), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1179), .B(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1161), .A2(new_n1170), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1168), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1161), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n1185), .A3(KEYINPUT61), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1173), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1157), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1172), .B1(new_n1154), .B2(new_n622), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1189), .B1(new_n1190), .B2(new_n1171), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n860), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1192));
  OAI211_X1 g767(.A(KEYINPUT119), .B(new_n1185), .C1(new_n1192), .C2(new_n1172), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1140), .A2(new_n1143), .A3(new_n1122), .A4(new_n1050), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1121), .B1(new_n1144), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n992), .A2(G290), .A3(G1986), .ZN(new_n1200));
  AND2_X1   g775(.A1(new_n1000), .A2(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT108), .Z(new_n1202));
  NAND4_X1  g777(.A1(new_n993), .A2(new_n996), .A3(new_n999), .A4(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1012), .B1(new_n1199), .B2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(new_n461), .A2(G227), .ZN(new_n1206));
  OAI21_X1  g780(.A(new_n1206), .B1(new_n664), .B2(new_n663), .ZN(new_n1207));
  OAI21_X1  g781(.A(KEYINPUT127), .B1(G229), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n1209));
  INV_X1    g783(.A(new_n1207), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n701), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI22_X1  g785(.A1(new_n906), .A2(new_n908), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  AND2_X1   g786(.A1(new_n1212), .A2(new_n968), .ZN(G308));
  NAND2_X1  g787(.A1(new_n1212), .A2(new_n968), .ZN(G225));
endmodule


