//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n542, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n593, new_n594, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT66), .Z(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n461), .A2(new_n462), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(new_n458), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  NOR2_X1   g046(.A1(new_n463), .A2(new_n458), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G124), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n477), .B1(new_n464), .B2(G136), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  NAND2_X1  g055(.A1(new_n468), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G126), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n458), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n464), .A2(G138), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n464), .A2(new_n488), .A3(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n487), .B2(new_n489), .ZN(G164));
  OR2_X1    g065(.A1(KEYINPUT5), .A2(G543), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT5), .A2(G543), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n493), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G50), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AND2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G88), .ZN(new_n505));
  OAI22_X1  g080(.A1(new_n498), .A2(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n496), .A2(new_n506), .ZN(G166));
  NAND3_X1  g082(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT7), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(G51), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n498), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n501), .A2(new_n500), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n497), .A2(G89), .ZN(new_n513));
  NAND2_X1  g088(.A1(G63), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n511), .A2(new_n515), .ZN(G168));
  INV_X1    g091(.A(G64), .ZN(new_n517));
  INV_X1    g092(.A(G77), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n512), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n522), .B1(new_n518), .B2(new_n519), .C1(new_n512), .C2(new_n517), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n521), .A2(G651), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(new_n504), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n525), .A2(G90), .B1(G52), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  AOI22_X1  g106(.A1(new_n493), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n495), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n498), .A2(new_n534), .B1(new_n504), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g114(.A(KEYINPUT70), .B(KEYINPUT8), .Z(new_n540));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  AND3_X1   g118(.A1(KEYINPUT71), .A2(G53), .A3(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(new_n502), .B2(new_n503), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT9), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT9), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n497), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  OAI21_X1  g123(.A(G65), .B1(new_n501), .B2(new_n500), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n546), .A2(new_n548), .B1(new_n551), .B2(G651), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n504), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n493), .A2(new_n497), .A3(KEYINPUT72), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G91), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  INV_X1    g133(.A(G166), .ZN(G303));
  AND2_X1   g134(.A1(new_n554), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G87), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n493), .A2(G74), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n528), .B2(G49), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(G288));
  NAND2_X1  g139(.A1(new_n560), .A2(G86), .ZN(new_n565));
  NAND2_X1  g140(.A1(G73), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n512), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(G48), .B2(new_n528), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n493), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n495), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n528), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G290));
  NAND2_X1  g149(.A1(G301), .A2(G868), .ZN(new_n575));
  INV_X1    g150(.A(G66), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n491), .B2(new_n492), .ZN(new_n577));
  NAND2_X1  g152(.A1(G79), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(KEYINPUT73), .A2(G79), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n577), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n528), .A2(G54), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n554), .A2(G92), .A3(new_n555), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n554), .A2(KEYINPUT10), .A3(G92), .A4(new_n555), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n575), .B1(G868), .B2(new_n590), .ZN(G284));
  OAI21_X1  g166(.A(new_n575), .B1(G868), .B2(new_n590), .ZN(G321));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(G299), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(new_n593), .B2(G168), .ZN(G297));
  XNOR2_X1  g170(.A(G297), .B(KEYINPUT74), .ZN(G280));
  INV_X1    g171(.A(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(G860), .ZN(G148));
  OR2_X1    g173(.A1(new_n533), .A2(new_n536), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(new_n593), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n588), .A2(new_n589), .ZN(new_n601));
  INV_X1    g176(.A(new_n585), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n600), .B1(new_n604), .B2(new_n593), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g181(.A1(new_n458), .A2(G2104), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n468), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT12), .Z(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT13), .Z(new_n610));
  INV_X1    g185(.A(G2100), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n473), .A2(G123), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n458), .A2(G111), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT75), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n614), .B2(KEYINPUT75), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n615), .A2(new_n617), .B1(new_n464), .B2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n610), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(G2096), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n612), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n634), .B(new_n635), .Z(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  AND3_X1   g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(G401));
  INV_X1    g214(.A(KEYINPUT18), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT77), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT17), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2100), .ZN(new_n648));
  NOR2_X1   g223(.A1(G2072), .A2(G2078), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n442), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n644), .B2(KEYINPUT18), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n660), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT79), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT78), .ZN(new_n667));
  XOR2_X1   g242(.A(G1981), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n665), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G288), .ZN(new_n673));
  INV_X1    g248(.A(G16), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(G23), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT33), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT81), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT32), .B(G1981), .Z(new_n679));
  AND2_X1   g254(.A1(new_n674), .A2(G6), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G305), .B2(G16), .ZN(new_n681));
  AOI22_X1  g256(.A1(new_n676), .A2(new_n678), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n678), .B2(new_n676), .ZN(new_n683));
  NOR2_X1   g258(.A1(G166), .A2(new_n674), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n674), .B2(G22), .ZN(new_n685));
  INV_X1    g260(.A(G1971), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(new_n688), .C1(new_n679), .C2(new_n681), .ZN(new_n689));
  OR3_X1    g264(.A1(new_n683), .A2(KEYINPUT34), .A3(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(KEYINPUT34), .B1(new_n683), .B2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(G290), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n674), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n674), .B2(G24), .ZN(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(KEYINPUT80), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(KEYINPUT80), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n473), .A2(G119), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n464), .B2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n700), .B(new_n701), .C1(new_n708), .C2(new_n698), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n696), .B(new_n697), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(new_n709), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n690), .A2(new_n691), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  OR2_X1    g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  NAND2_X1  g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n716), .A2(new_n698), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n619), .B2(new_n698), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n674), .A2(G21), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G168), .B2(new_n674), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n720), .B1(G1966), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  NOR2_X1   g299(.A1(G171), .A2(new_n674), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G5), .B2(new_n674), .ZN(new_n726));
  OAI221_X1 g301(.A(new_n723), .B1(G1966), .B2(new_n722), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT86), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n464), .A2(G139), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT83), .Z(new_n730));
  NAND3_X1  g305(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT82), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n468), .A2(G127), .ZN(new_n734));
  AND2_X1   g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(G2105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(G33), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  AND2_X1   g314(.A1(new_n698), .A2(G32), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n473), .A2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n464), .A2(G141), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT84), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT26), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n747), .A2(new_n748), .B1(G105), .B2(new_n607), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n741), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT85), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n744), .A2(new_n741), .A3(new_n752), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n740), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT87), .B(KEYINPUT23), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n674), .A2(G20), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1956), .Z(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n726), .B2(new_n724), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n739), .A2(new_n757), .A3(new_n758), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n698), .A2(G26), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT28), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n473), .A2(G128), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(G116), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G2105), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n464), .B2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G2067), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n674), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n537), .B2(new_n674), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n780), .A2(KEYINPUT24), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(KEYINPUT24), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n698), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G160), .B2(new_n698), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2084), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n776), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G27), .A2(G29), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G164), .B2(G29), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G35), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G162), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT29), .B(G2090), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n786), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n674), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n590), .B2(new_n674), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1348), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n728), .A2(new_n765), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n715), .A2(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  INV_X1    g376(.A(KEYINPUT88), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n525), .A2(G93), .B1(G55), .B2(new_n528), .ZN(new_n803));
  OAI21_X1  g378(.A(G67), .B1(new_n501), .B2(new_n500), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n495), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n802), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n498), .A2(new_n809), .B1(new_n504), .B2(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n811), .A2(KEYINPUT88), .A3(new_n806), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n599), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n803), .A2(new_n802), .A3(new_n807), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT88), .B1(new_n811), .B2(new_n806), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n814), .A2(new_n537), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT38), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n590), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  INV_X1    g396(.A(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n811), .A2(new_n806), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n822), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(G145));
  XOR2_X1   g403(.A(new_n479), .B(new_n619), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G160), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n473), .A2(G130), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  INV_X1    g407(.A(G118), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(G2105), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n464), .B2(G142), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n751), .A2(new_n753), .A3(new_n773), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n773), .B1(new_n751), .B2(new_n753), .ZN(new_n839));
  OAI21_X1  g414(.A(G164), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n839), .ZN(new_n841));
  INV_X1    g416(.A(G164), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n837), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT90), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n737), .B2(KEYINPUT89), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n840), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n737), .A2(new_n844), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n840), .A2(new_n843), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n836), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n836), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n840), .A2(new_n843), .A3(new_n845), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n840), .A2(new_n843), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n847), .A2(new_n845), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n707), .B(new_n609), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT91), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n849), .B2(new_n854), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n830), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n849), .A2(new_n854), .ZN(new_n861));
  INV_X1    g436(.A(new_n855), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n830), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n863), .A2(KEYINPUT91), .A3(new_n864), .A4(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g442(.A(G299), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n603), .A2(KEYINPUT93), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT93), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n590), .B2(G299), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n585), .B1(new_n552), .B2(new_n556), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n601), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(KEYINPUT94), .A3(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT92), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n601), .A2(new_n872), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n601), .B2(new_n872), .ZN(new_n883));
  OAI21_X1  g458(.A(KEYINPUT41), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n869), .A2(new_n871), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT93), .B1(new_n603), .B2(new_n868), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n590), .A2(new_n870), .A3(G299), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n873), .A2(KEYINPUT92), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n875), .B1(new_n891), .B2(new_n881), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT95), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n878), .B(new_n879), .C1(new_n887), .C2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n604), .B(new_n817), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(KEYINPUT97), .A2(KEYINPUT42), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n869), .B(new_n871), .C1(new_n882), .C2(new_n883), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  OR3_X1    g475(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n692), .ZN(new_n902));
  NAND2_X1  g477(.A1(G288), .A2(G290), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT96), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT96), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G305), .B(G303), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n909), .B1(new_n904), .B2(KEYINPUT96), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(KEYINPUT97), .B2(KEYINPUT42), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n897), .B1(new_n896), .B2(new_n900), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n901), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n914), .B1(new_n901), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g492(.A(G868), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g494(.A(new_n918), .B1(G868), .B2(new_n825), .ZN(G331));
  NAND2_X1  g495(.A1(G301), .A2(G286), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n524), .A2(G168), .A3(new_n529), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n813), .A2(new_n921), .A3(new_n816), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT100), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n524), .A2(G168), .A3(new_n529), .ZN(new_n925));
  AOI21_X1  g500(.A(G168), .B1(new_n524), .B2(new_n529), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n816), .A4(new_n813), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n817), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT99), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n817), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  AND4_X1   g510(.A1(new_n898), .A2(new_n930), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n923), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n894), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT43), .B1(new_n938), .B2(new_n913), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n910), .B2(new_n912), .ZN(new_n941));
  INV_X1    g516(.A(new_n909), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n905), .B2(new_n907), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n943), .A2(new_n911), .A3(KEYINPUT102), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n938), .B2(new_n946), .ZN(new_n947));
  AOI211_X1 g522(.A(KEYINPUT101), .B(new_n936), .C1(new_n894), .C2(new_n937), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n860), .B(new_n939), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n930), .A2(new_n933), .A3(new_n935), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n950), .B(new_n951), .C1(KEYINPUT41), .C2(new_n898), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n952), .B1(new_n899), .B2(new_n937), .ZN(new_n953));
  AOI21_X1  g528(.A(G37), .B1(new_n953), .B2(new_n945), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n938), .A2(new_n913), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  OAI211_X1 g534(.A(KEYINPUT44), .B(new_n949), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n860), .B(new_n956), .C1(new_n947), .C2(new_n948), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n961), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT103), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n954), .A2(new_n939), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT98), .B(KEYINPUT44), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(G397));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(G164), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(G160), .A2(G40), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G1996), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT46), .Z(new_n974));
  INV_X1    g549(.A(new_n972), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n773), .A2(G2067), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n768), .A2(new_n775), .A3(new_n772), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n978), .B2(new_n754), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT124), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT47), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n972), .A2(G1986), .A3(G290), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(G1996), .A3(new_n754), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT106), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n975), .B2(new_n978), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n973), .A2(new_n751), .A3(new_n753), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT105), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n707), .A2(new_n711), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n708), .A2(new_n710), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n975), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT125), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT125), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n988), .A2(new_n996), .A3(new_n990), .A4(new_n993), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n985), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n972), .B1(new_n999), .B2(new_n977), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n983), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(G164), .A2(G1384), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1003), .A2(new_n971), .A3(new_n969), .ZN(new_n1004));
  INV_X1    g579(.A(G1966), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n971), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1002), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1006), .B(G168), .C1(G2084), .C2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(G8), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1012), .A2(new_n1016), .A3(G8), .A4(new_n1013), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1012), .A2(G8), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1015), .B(new_n1017), .C1(KEYINPUT51), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1011), .A2(G2084), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n1021), .B2(new_n1006), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G286), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1025));
  INV_X1    g600(.A(G2090), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1008), .A2(new_n1026), .A3(new_n1010), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT108), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1008), .A2(new_n1029), .A3(new_n1026), .A4(new_n1010), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1004), .A2(new_n686), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n1033), .B(KEYINPUT55), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(G8), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(G305), .A2(G1981), .ZN(new_n1039));
  INV_X1    g614(.A(G86), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n569), .B1(new_n1040), .B2(new_n504), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G1981), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(KEYINPUT49), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1039), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1020), .B1(new_n971), .B2(new_n1002), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1045), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1976), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1047), .B1(new_n1054), .B2(G288), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(KEYINPUT110), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(KEYINPUT110), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1047), .B(new_n1058), .C1(new_n1054), .C2(G288), .ZN(new_n1059));
  NAND3_X1  g634(.A1(G288), .A2(new_n1056), .A3(new_n1054), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1053), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n971), .A2(new_n1007), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1010), .A2(KEYINPUT114), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1002), .A2(new_n1065), .A3(new_n1009), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1067), .A2(new_n1026), .B1(new_n686), .B2(new_n1004), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1034), .B1(new_n1068), .B2(new_n1020), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(KEYINPUT115), .B(new_n1034), .C1(new_n1068), .C2(new_n1020), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1062), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1038), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1019), .A2(new_n1075), .A3(new_n1023), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1011), .A2(new_n724), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1003), .A2(new_n969), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n789), .A4(new_n971), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1004), .B2(G2078), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(KEYINPUT122), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(KEYINPUT122), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1077), .B(new_n1079), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(G171), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1025), .A2(new_n1074), .A3(new_n1076), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1067), .A2(G1956), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT56), .B(G2072), .Z(new_n1089));
  NOR2_X1   g664(.A1(new_n1004), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(G299), .B(KEYINPUT57), .Z(new_n1092));
  OAI21_X1  g667(.A(new_n1087), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1092), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT117), .B(new_n1094), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1095));
  INV_X1    g670(.A(G1348), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n971), .A2(new_n1002), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1011), .A2(new_n1096), .B1(new_n775), .B2(new_n1098), .ZN(new_n1099));
  OR3_X1    g674(.A1(new_n1099), .A2(KEYINPUT116), .A3(new_n603), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT116), .B1(new_n1099), .B2(new_n603), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1093), .A2(new_n1095), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT61), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1103), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n1099), .A2(new_n603), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1099), .A2(new_n603), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1099), .A2(new_n1111), .A3(new_n590), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT58), .B(G1341), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1004), .A2(G1996), .B1(new_n1098), .B2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n537), .A2(KEYINPUT118), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(KEYINPUT59), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT59), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1091), .A2(new_n1105), .A3(new_n1092), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1107), .A2(new_n1110), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1104), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(G301), .B(KEYINPUT54), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1084), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT53), .B(new_n789), .C1(new_n971), .C2(KEYINPUT123), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(KEYINPUT123), .B2(new_n971), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1123), .B1(new_n1126), .B2(new_n1078), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(new_n1077), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1023), .B2(new_n1019), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1122), .A2(new_n1074), .A3(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1053), .A2(new_n1022), .A3(G168), .A4(new_n1061), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1035), .B1(new_n1032), .B2(G8), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT63), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n673), .A2(new_n1054), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT113), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1136), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1039), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1047), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1022), .A2(G168), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(KEYINPUT63), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1038), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1062), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1086), .A2(new_n1131), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G290), .B(G1986), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n975), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n988), .A2(new_n990), .A3(new_n993), .A4(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT107), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1001), .B1(new_n1147), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g727(.A1(new_n653), .A2(G319), .ZN(new_n1154));
  XNOR2_X1  g728(.A(new_n1154), .B(KEYINPUT126), .ZN(new_n1155));
  NOR3_X1   g729(.A1(G229), .A2(new_n1155), .A3(G401), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n866), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g731(.A1(new_n965), .A2(new_n1157), .ZN(G308));
  OR2_X1    g732(.A1(new_n963), .A2(new_n964), .ZN(new_n1159));
  OAI211_X1 g733(.A(new_n866), .B(new_n1156), .C1(new_n1159), .C2(new_n962), .ZN(G225));
endmodule


