//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT67), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(new_n190), .B2(G116), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n187), .A2(KEYINPUT68), .A3(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n197), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n199), .A2(new_n192), .A3(new_n194), .A4(new_n195), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT65), .A3(G143), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(new_n202), .B2(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n205), .A3(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n212), .A3(new_n204), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G128), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n207), .A2(new_n209), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G137), .ZN(new_n219));
  INV_X1    g033(.A(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(G137), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n218), .A2(G137), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n220), .A2(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n198), .B(new_n200), .C1(new_n216), .C2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n213), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n203), .A2(new_n206), .A3(new_n204), .A4(new_n230), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT69), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n224), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n229), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT74), .B1(new_n241), .B2(KEYINPUT28), .ZN(new_n242));
  INV_X1    g056(.A(new_n229), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n234), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n234), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n240), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n242), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n246), .A2(KEYINPUT70), .A3(new_n240), .A4(new_n247), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(new_n243), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n213), .A2(new_n215), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n203), .A2(new_n206), .A3(new_n209), .A4(new_n204), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n224), .A2(new_n227), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT66), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n233), .A2(new_n234), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n240), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n198), .A2(new_n200), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n257), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT28), .ZN(new_n272));
  XOR2_X1   g086(.A(KEYINPUT26), .B(G101), .Z(new_n273));
  INV_X1    g087(.A(G237), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(G210), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n273), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT73), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n253), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n269), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n268), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n255), .A2(KEYINPUT30), .A3(new_n262), .A4(new_n256), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n257), .ZN(new_n287));
  INV_X1    g101(.A(new_n279), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n288), .A2(new_n290), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n255), .A2(new_n256), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n255), .A2(new_n262), .A3(new_n256), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n293), .A2(new_n243), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n253), .B(new_n292), .C1(new_n295), .C2(new_n251), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G472), .B1(new_n291), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n284), .A2(new_n285), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n257), .A2(new_n279), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT31), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n280), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n242), .A2(new_n252), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n251), .B1(new_n257), .B2(new_n270), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n307));
  NAND4_X1  g121(.A1(new_n286), .A2(new_n279), .A3(new_n257), .A4(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n302), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(KEYINPUT32), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(KEYINPUT32), .A3(new_n310), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n299), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n190), .A2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n208), .A2(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT77), .A2(KEYINPUT23), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT77), .B(KEYINPUT23), .Z(new_n322));
  OAI211_X1 g136(.A(new_n318), .B(new_n321), .C1(new_n322), .C2(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G110), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT78), .ZN(new_n325));
  OR2_X1    g139(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n318), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  OR2_X1    g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT16), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n333), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  AOI21_X1  g150(.A(G146), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n335), .A2(new_n336), .A3(G146), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n323), .A2(new_n341), .A3(G110), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n325), .A2(new_n330), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n328), .A2(new_n329), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n344), .B1(new_n323), .B2(G110), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n205), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n339), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n348), .A3(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n297), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n317), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n357), .B2(new_n356), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n317), .A3(new_n357), .ZN(new_n360));
  INV_X1    g174(.A(G217), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(G234), .B2(new_n297), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n354), .A2(new_n355), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n362), .A2(G902), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n359), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n316), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G478), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT15), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT93), .B1(new_n187), .B2(G122), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT93), .ZN(new_n372));
  INV_X1    g186(.A(G122), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G116), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT94), .B1(new_n373), .B2(G116), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT94), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n187), .A3(G122), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n376), .B2(new_n378), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT96), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n375), .B(new_n380), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AOI211_X1 g197(.A(KEYINPUT96), .B(new_n379), .C1(new_n376), .C2(new_n378), .ZN(new_n384));
  OAI21_X1  g198(.A(G107), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT97), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT97), .B(G107), .C1(new_n383), .C2(new_n384), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(new_n378), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n375), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT95), .B1(new_n208), .B2(G143), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n202), .A3(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n208), .A2(G143), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n218), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n218), .B1(new_n395), .B2(new_n396), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n391), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n387), .A2(new_n388), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n375), .A2(new_n389), .A3(new_n390), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n390), .B1(new_n375), .B2(new_n389), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT13), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n395), .A2(new_n406), .B1(new_n208), .B2(G143), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT13), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n218), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n402), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT9), .B(G234), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n413), .A2(new_n361), .A3(G953), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n402), .A2(new_n411), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT98), .B1(new_n418), .B2(new_n297), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n400), .B1(new_n385), .B2(new_n386), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n415), .B(new_n410), .C1(new_n420), .C2(new_n388), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n402), .B2(new_n411), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT98), .B(new_n297), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n370), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n369), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G113), .B(G122), .ZN(new_n428));
  INV_X1    g242(.A(G104), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n274), .A2(new_n275), .A3(G214), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(G143), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n222), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n432), .B(new_n202), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(KEYINPUT18), .A3(G131), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n346), .B(new_n205), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n441));
  INV_X1    g255(.A(new_n339), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n337), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT90), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(KEYINPUT17), .A3(G131), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT17), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n433), .B(G131), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n446), .A2(KEYINPUT91), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT91), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n443), .A2(new_n444), .A3(new_n450), .A4(new_n445), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n431), .B(new_n440), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n446), .A2(KEYINPUT91), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n447), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n430), .B1(new_n455), .B2(new_n439), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n297), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G475), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n275), .A2(G952), .ZN(new_n459));
  INV_X1    g273(.A(G234), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n274), .ZN(new_n461));
  XOR2_X1   g275(.A(new_n461), .B(KEYINPUT99), .Z(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(G902), .B(G953), .C1(new_n460), .C2(new_n274), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT100), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT21), .B(G898), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT101), .Z(new_n468));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n430), .A3(new_n439), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n346), .B(KEYINPUT19), .Z(new_n471));
  OAI21_X1  g285(.A(new_n339), .B1(new_n471), .B2(G146), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n472), .A2(new_n448), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n430), .B1(new_n473), .B2(new_n439), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(G475), .A2(G902), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT92), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n469), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g294(.A(KEYINPUT20), .B(new_n478), .C1(new_n470), .C2(new_n475), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n458), .B(new_n468), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n427), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G113), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n187), .A2(G119), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT5), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n196), .B2(new_n488), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n200), .ZN(new_n491));
  OR2_X1    g305(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n390), .A2(G104), .ZN(new_n493));
  AND2_X1   g307(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G101), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n429), .A2(G107), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n429), .A2(G107), .ZN(new_n498));
  NOR2_X1   g312(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n390), .A2(G104), .ZN(new_n502));
  OAI21_X1  g316(.A(G101), .B1(new_n502), .B2(new_n498), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n491), .A2(KEYINPUT86), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT86), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n490), .B(new_n200), .C1(new_n504), .C2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G110), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT8), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G224), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT7), .B1(new_n512), .B2(G953), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n258), .A2(new_n333), .A3(new_n259), .ZN(new_n514));
  OR2_X1    g328(.A1(new_n514), .A2(KEYINPUT87), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n266), .B2(new_n333), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n513), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n516), .A2(new_n513), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n497), .B1(new_n492), .B2(new_n493), .ZN(new_n520));
  NAND2_X1  g334(.A1(KEYINPUT81), .A2(KEYINPUT3), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n499), .B1(new_n498), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G101), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT4), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n525), .B(G101), .C1(new_n520), .C2(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n269), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n505), .A2(new_n200), .A3(new_n490), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n509), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n511), .A2(new_n518), .A3(new_n519), .A4(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n530), .A2(new_n297), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n528), .ZN(new_n532));
  INV_X1    g346(.A(new_n509), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT6), .A3(new_n529), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n512), .A2(G953), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n516), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G210), .B1(G237), .B2(G902), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT89), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n531), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n545), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n548), .A3(new_n540), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n485), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G221), .B1(new_n413), .B2(G902), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT80), .ZN(new_n552));
  INV_X1    g366(.A(G469), .ZN(new_n553));
  XNOR2_X1  g367(.A(G110), .B(G140), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n275), .A2(G227), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n557));
  NAND3_X1  g371(.A1(new_n203), .A2(new_n204), .A3(new_n206), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n215), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n559), .A2(new_n259), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n560), .B2(new_n504), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n259), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n503), .A3(new_n501), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n557), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n504), .A2(new_n216), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n502), .B1(new_n498), .B2(new_n499), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT4), .B(new_n496), .C1(new_n570), .C2(new_n495), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n523), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n573), .B2(new_n237), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n240), .B(KEYINPUT84), .Z(new_n575));
  AND3_X1   g389(.A1(new_n567), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n240), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n567), .B2(new_n574), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT85), .B(new_n556), .C1(new_n576), .C2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n564), .B1(new_n505), .B2(new_n260), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n240), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(KEYINPUT12), .A3(new_n240), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n567), .A2(new_n574), .A3(new_n575), .ZN(new_n586));
  INV_X1    g400(.A(new_n556), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n564), .A2(new_n565), .A3(new_n557), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n565), .B1(new_n564), .B2(new_n557), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n505), .A2(KEYINPUT10), .A3(new_n260), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n246), .A2(new_n247), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n524), .A2(new_n526), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n240), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n586), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT85), .B1(new_n598), .B2(new_n556), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n553), .B(new_n297), .C1(new_n589), .C2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n576), .A2(new_n556), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n585), .A2(new_n586), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n601), .A2(new_n597), .B1(new_n602), .B2(new_n556), .ZN(new_n603));
  OAI21_X1  g417(.A(G469), .B1(new_n603), .B2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n552), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n483), .A2(new_n550), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n367), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(new_n496), .ZN(G3));
  NAND2_X1  g422(.A1(new_n600), .A2(new_n604), .ZN(new_n609));
  INV_X1    g423(.A(new_n552), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n366), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n309), .B2(new_n297), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n311), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(KEYINPUT102), .B(new_n612), .C1(new_n309), .C2(new_n297), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n549), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n548), .B1(new_n531), .B2(new_n540), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n484), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n416), .A2(KEYINPUT103), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n418), .A2(new_n621), .A3(KEYINPUT33), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n416), .B(new_n417), .C1(KEYINPUT103), .C2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(G478), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n297), .B1(new_n421), .B2(new_n422), .ZN(new_n626));
  MUX2_X1   g440(.A(new_n297), .B(new_n626), .S(new_n368), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n440), .B1(new_n449), .B2(new_n451), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n474), .B1(new_n629), .B2(new_n430), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT20), .B1(new_n630), .B2(new_n478), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n476), .A2(new_n469), .A3(new_n479), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n631), .A2(new_n632), .B1(G475), .B2(new_n457), .ZN(new_n633));
  INV_X1    g447(.A(new_n468), .ZN(new_n634));
  NOR4_X1   g448(.A1(new_n620), .A2(new_n628), .A3(new_n633), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n617), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT104), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT34), .B(G104), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G6));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n626), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n369), .B1(new_n641), .B2(new_n423), .ZN(new_n642));
  INV_X1    g456(.A(new_n426), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n458), .B1(new_n480), .B2(new_n481), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n644), .A2(new_n620), .A3(new_n645), .A4(new_n634), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n617), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n349), .A2(KEYINPUT105), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n349), .A2(KEYINPUT105), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n656), .A2(new_n365), .B1(new_n359), .B2(new_n363), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n483), .A2(new_n658), .A3(new_n550), .A4(new_n605), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n309), .A2(new_n297), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G472), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n613), .A2(new_n614), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n311), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n465), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT106), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n462), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n644), .A2(new_n620), .A3(new_n645), .A4(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(new_n316), .A3(new_n605), .A4(new_n658), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XNOR2_X1  g489(.A(new_n671), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n605), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  AOI21_X1  g492(.A(new_n548), .B1(new_n541), .B2(new_n542), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n618), .B1(new_n679), .B2(new_n546), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n681), .A2(new_n485), .A3(new_n644), .A4(new_n633), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n300), .A2(new_n301), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n294), .A2(new_n269), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n257), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n683), .B1(new_n303), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n314), .A2(new_n315), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n678), .A2(new_n682), .A3(new_n657), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  AND3_X1   g504(.A1(new_n316), .A2(new_n605), .A3(new_n658), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n628), .A2(new_n633), .A3(new_n672), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n541), .A2(new_n545), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n485), .B1(new_n694), .B2(new_n549), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n645), .A2(new_n625), .A3(new_n627), .A4(new_n671), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT107), .B1(new_n697), .B2(new_n620), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n691), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  OAI21_X1  g514(.A(new_n297), .B1(new_n589), .B2(new_n599), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n600), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n367), .A2(new_n552), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n635), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n646), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  AND2_X1   g523(.A1(new_n702), .A2(new_n600), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n483), .A3(new_n610), .A4(new_n695), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n316), .A2(new_n658), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT108), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n304), .B1(new_n685), .B2(KEYINPUT28), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n292), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n281), .A2(new_n289), .A3(new_n290), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n612), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND3_X1   g531(.A1(new_n309), .A2(KEYINPUT32), .A3(new_n310), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n657), .B1(new_n719), .B2(new_n314), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n702), .A2(new_n610), .A3(new_n600), .A4(new_n695), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n644), .A2(new_n633), .A3(new_n468), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n713), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR2_X1   g541(.A1(new_n714), .A2(new_n280), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n302), .A2(new_n308), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n310), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n661), .A2(new_n366), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n427), .A2(new_n645), .A3(new_n468), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n721), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n373), .ZN(G24));
  NAND2_X1  g548(.A1(new_n661), .A2(new_n730), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n735), .A2(new_n697), .A3(new_n657), .ZN(new_n736));
  INV_X1    g550(.A(new_n721), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(new_n366), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n719), .B2(new_n314), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n552), .A2(new_n485), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n600), .B2(new_n604), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n680), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT109), .B1(new_n745), .B2(new_n680), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n741), .B(new_n742), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT32), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n311), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n299), .A2(new_n750), .A3(new_n315), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n366), .A3(new_n692), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n745), .A2(new_n680), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n680), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n748), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n222), .ZN(G33));
  NOR3_X1   g574(.A1(new_n644), .A2(new_n645), .A3(new_n672), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n741), .B(new_n761), .C1(new_n746), .C2(new_n747), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n603), .A2(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n603), .A2(KEYINPUT45), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(G469), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(G469), .A2(G902), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT46), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n768), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n600), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n610), .ZN(new_n774));
  INV_X1    g588(.A(new_n676), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n764), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(KEYINPUT110), .A3(new_n610), .A4(new_n676), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n680), .A2(new_n484), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n664), .A2(new_n658), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT112), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n628), .A2(new_n645), .A3(KEYINPUT43), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n645), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n633), .A2(KEYINPUT111), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n625), .A4(new_n627), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n782), .B1(new_n786), .B2(KEYINPUT43), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n781), .A2(KEYINPUT44), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n787), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT44), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n779), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(KEYINPUT113), .B(G137), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G39));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n774), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n773), .A2(KEYINPUT47), .A3(new_n610), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n778), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n799), .A2(new_n316), .A3(new_n366), .A4(new_n697), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  AND2_X1   g616(.A1(new_n787), .A2(new_n463), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n740), .B1(new_n719), .B2(new_n750), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n703), .A2(new_n552), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n805), .A2(new_n778), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT48), .ZN(new_n808));
  INV_X1    g622(.A(new_n731), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(new_n737), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n628), .A2(new_n633), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n688), .A2(new_n740), .A3(new_n462), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n806), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n808), .A2(new_n459), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT118), .Z(new_n815));
  NOR2_X1   g629(.A1(new_n735), .A2(new_n657), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n803), .A2(new_n816), .A3(new_n806), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n806), .A2(new_n812), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n628), .A2(new_n633), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n796), .B(new_n797), .C1(new_n610), .C2(new_n703), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n803), .A2(new_n809), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n799), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n820), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n681), .A2(new_n485), .A3(new_n805), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n822), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(KEYINPUT50), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT50), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n830), .A3(new_n822), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n824), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT51), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n815), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n665), .A2(new_n607), .A3(new_n733), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n741), .B(new_n805), .C1(new_n635), .C2(new_n646), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n680), .A2(new_n485), .A3(new_n634), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n425), .B2(new_n426), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT114), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n839), .B(new_n633), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n811), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n425), .A2(new_n840), .A3(new_n426), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT114), .B1(new_n642), .B2(new_n643), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n839), .B1(new_n848), .B2(new_n633), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n617), .B(new_n838), .C1(new_n845), .C2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n836), .A2(new_n726), .A3(new_n837), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n755), .A2(new_n756), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n680), .A2(new_n484), .A3(new_n633), .A4(new_n671), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n848), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n852), .A2(new_n736), .B1(new_n691), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n746), .A2(new_n747), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT42), .B1(new_n856), .B2(new_n752), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n857), .A3(new_n748), .A4(new_n762), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n738), .A2(new_n674), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n688), .A2(new_n657), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n644), .A2(new_n620), .A3(new_n633), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n605), .A3(new_n671), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n699), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n696), .A2(new_n698), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n316), .A2(new_n605), .A3(new_n658), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n738), .B(new_n674), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n863), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT52), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  NOR4_X1   g685(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n722), .A4(new_n721), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n850), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n483), .A2(new_n550), .A3(new_n605), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n741), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n615), .A2(new_n616), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n877), .A3(new_n658), .ZN(new_n878));
  INV_X1    g692(.A(new_n733), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n837), .A2(new_n876), .A3(new_n878), .A4(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n691), .A2(new_n854), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n736), .B1(new_n746), .B2(new_n747), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n762), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n759), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n881), .A2(new_n885), .A3(new_n865), .A4(new_n870), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT53), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n871), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT54), .B1(new_n871), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n835), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n886), .A2(new_n887), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n886), .A2(new_n887), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n871), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(KEYINPUT116), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  OAI22_X1  g712(.A1(new_n834), .A2(new_n898), .B1(G952), .B2(G953), .ZN(new_n899));
  INV_X1    g713(.A(new_n681), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n786), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n710), .B(KEYINPUT49), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n688), .A2(new_n740), .A3(new_n744), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n904), .ZN(G75));
  NAND2_X1  g719(.A1(new_n871), .A2(new_n888), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(G902), .A3(new_n545), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n535), .A2(new_n537), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(new_n539), .Z(new_n909));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n907), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n907), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n275), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  NOR2_X1   g732(.A1(new_n889), .A2(new_n890), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n768), .B(KEYINPUT57), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n599), .B2(new_n589), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n906), .A2(G902), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(new_n767), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n917), .B1(new_n922), .B2(new_n924), .ZN(G54));
  NAND4_X1  g739(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n630), .ZN(new_n927));
  INV_X1    g741(.A(new_n917), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n926), .B2(new_n630), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT121), .B1(new_n926), .B2(new_n630), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(G60));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n622), .A2(new_n624), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n368), .A2(new_n297), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  AND2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n932), .B1(new_n919), .B2(new_n936), .ZN(new_n937));
  AND4_X1   g751(.A1(new_n932), .A2(new_n895), .A3(new_n896), .A4(new_n936), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n928), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n898), .B2(new_n935), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(G63));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n361), .A2(new_n297), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n906), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n656), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n928), .B1(new_n946), .B2(new_n364), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n946), .A2(new_n364), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n947), .A3(KEYINPUT61), .A4(new_n928), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n466), .B2(new_n512), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n881), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n908), .B1(G898), .B2(new_n275), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  INV_X1    g771(.A(new_n268), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n285), .B1(KEYINPUT30), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n471), .Z(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(G900), .B2(G953), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n801), .A2(new_n762), .ZN(new_n963));
  INV_X1    g777(.A(new_n759), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n868), .B(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n776), .A2(new_n804), .A3(new_n777), .A4(new_n862), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n963), .A2(new_n964), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n792), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n962), .B1(new_n970), .B2(new_n275), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n367), .A2(new_n799), .A3(new_n677), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n849), .B2(new_n845), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n792), .A2(new_n801), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n966), .A2(new_n689), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(KEYINPUT62), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT126), .ZN(new_n982));
  AOI21_X1  g796(.A(G953), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n960), .B(KEYINPUT124), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n972), .B(new_n974), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n978), .B2(KEYINPUT62), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n977), .B(new_n979), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n984), .B1(new_n989), .B2(new_n275), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n973), .B1(new_n990), .B2(new_n971), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n985), .A2(new_n991), .ZN(G72));
  XNOR2_X1  g806(.A(new_n287), .B(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n279), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n980), .A2(new_n982), .A3(new_n881), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n993), .A2(new_n279), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n968), .A2(new_n969), .A3(new_n851), .ZN(new_n1000));
  INV_X1    g814(.A(new_n997), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n683), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1003), .B2(new_n289), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n917), .B1(new_n906), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n998), .A2(new_n1006), .ZN(G57));
endmodule


