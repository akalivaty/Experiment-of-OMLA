

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576;

  XNOR2_X1 U321 ( .A(n373), .B(n372), .ZN(n569) );
  NOR2_X1 U322 ( .A1(n448), .A2(n376), .ZN(n377) );
  XNOR2_X1 U323 ( .A(n429), .B(n367), .ZN(n368) );
  XNOR2_X1 U324 ( .A(n369), .B(n368), .ZN(n370) );
  INV_X1 U325 ( .A(G211GAT), .ZN(n445) );
  XNOR2_X1 U326 ( .A(n444), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U327 ( .A(n569), .B(n374), .ZN(n553) );
  XNOR2_X1 U328 ( .A(n445), .B(KEYINPUT126), .ZN(n446) );
  XNOR2_X1 U329 ( .A(n447), .B(n446), .ZN(G1354GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n290) );
  XNOR2_X1 U331 ( .A(G57GAT), .B(G64GAT), .ZN(n289) );
  XNOR2_X1 U332 ( .A(n290), .B(n289), .ZN(n306) );
  XOR2_X1 U333 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n292) );
  NAND2_X1 U334 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U336 ( .A(n293), .B(KEYINPUT14), .Z(n298) );
  XNOR2_X1 U337 ( .A(G15GAT), .B(G22GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n294), .B(KEYINPUT72), .ZN(n358) );
  XOR2_X1 U339 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n296) );
  XNOR2_X1 U340 ( .A(G71GAT), .B(KEYINPUT73), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n365) );
  XNOR2_X1 U342 ( .A(n358), .B(n365), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U344 ( .A(G8GAT), .B(KEYINPUT82), .Z(n330) );
  XOR2_X1 U345 ( .A(G1GAT), .B(G127GAT), .Z(n311) );
  XOR2_X1 U346 ( .A(n330), .B(n311), .Z(n300) );
  XNOR2_X1 U347 ( .A(G155GAT), .B(G78GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U349 ( .A(n302), .B(n301), .Z(n304) );
  XNOR2_X1 U350 ( .A(G183GAT), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U352 ( .A(n306), .B(n305), .Z(n448) );
  INV_X1 U353 ( .A(n448), .ZN(n558) );
  XOR2_X1 U354 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n308) );
  XNOR2_X1 U355 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n320) );
  XOR2_X1 U357 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n310) );
  XNOR2_X1 U358 ( .A(G85GAT), .B(KEYINPUT4), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n312) );
  XOR2_X1 U360 ( .A(n312), .B(n311), .Z(n318) );
  XOR2_X1 U361 ( .A(G113GAT), .B(KEYINPUT0), .Z(n412) );
  XNOR2_X1 U362 ( .A(G120GAT), .B(G148GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n313), .B(G57GAT), .ZN(n366) );
  XOR2_X1 U364 ( .A(G29GAT), .B(G134GAT), .Z(n382) );
  XOR2_X1 U365 ( .A(n366), .B(n382), .Z(n315) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U368 ( .A(n412), .B(n316), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT3), .B(KEYINPUT89), .Z(n322) );
  XNOR2_X1 U372 ( .A(G141GAT), .B(G155GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT2), .Z(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n440) );
  XNOR2_X1 U376 ( .A(n325), .B(n440), .ZN(n455) );
  XNOR2_X1 U377 ( .A(KEYINPUT95), .B(n455), .ZN(n504) );
  XOR2_X1 U378 ( .A(G211GAT), .B(KEYINPUT21), .Z(n327) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n431) );
  XOR2_X1 U381 ( .A(n431), .B(KEYINPUT96), .Z(n329) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n331) );
  XOR2_X1 U384 ( .A(n331), .B(n330), .Z(n336) );
  XOR2_X1 U385 ( .A(G92GAT), .B(G64GAT), .Z(n333) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(G204GAT), .B(n334), .Z(n364) );
  XOR2_X1 U389 ( .A(G36GAT), .B(G190GAT), .Z(n391) );
  XNOR2_X1 U390 ( .A(n364), .B(n391), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n341) );
  XNOR2_X1 U392 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n337), .B(KEYINPUT18), .ZN(n338) );
  XOR2_X1 U394 ( .A(n338), .B(KEYINPUT87), .Z(n340) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(G183GAT), .ZN(n339) );
  XOR2_X1 U396 ( .A(n340), .B(n339), .Z(n422) );
  XNOR2_X1 U397 ( .A(n341), .B(n422), .ZN(n452) );
  XOR2_X1 U398 ( .A(G113GAT), .B(G29GAT), .Z(n343) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G36GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U401 ( .A(G1GAT), .B(G141GAT), .Z(n345) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G197GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n347), .B(n346), .Z(n352) );
  XOR2_X1 U405 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n349) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U408 ( .A(KEYINPUT68), .B(n350), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U410 ( .A(KEYINPUT71), .B(KEYINPUT69), .Z(n354) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(KEYINPUT70), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U413 ( .A(n356), .B(n355), .Z(n360) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n357) );
  XNOR2_X1 U415 ( .A(n357), .B(KEYINPUT7), .ZN(n393) );
  XNOR2_X1 U416 ( .A(n393), .B(n358), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n565) );
  XOR2_X1 U418 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n362) );
  XNOR2_X1 U419 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n373) );
  XOR2_X1 U422 ( .A(G99GAT), .B(G85GAT), .Z(n381) );
  XOR2_X1 U423 ( .A(n365), .B(n381), .Z(n371) );
  XOR2_X1 U424 ( .A(n366), .B(KEYINPUT77), .Z(n369) );
  XOR2_X1 U425 ( .A(G106GAT), .B(G78GAT), .Z(n429) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n374) );
  NOR2_X1 U429 ( .A1(n565), .A2(n553), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  XNOR2_X1 U431 ( .A(KEYINPUT112), .B(n377), .ZN(n398) );
  XOR2_X1 U432 ( .A(G92GAT), .B(G106GAT), .Z(n379) );
  NAND2_X1 U433 ( .A1(G232GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U435 ( .A(G162GAT), .B(n380), .ZN(n397) );
  XOR2_X1 U436 ( .A(KEYINPUT9), .B(KEYINPUT80), .Z(n384) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U439 ( .A(n385), .B(KEYINPUT11), .Z(n390) );
  XOR2_X1 U440 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n387) );
  XNOR2_X1 U441 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U443 ( .A(G218GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U445 ( .A(n392), .B(n391), .Z(n395) );
  XOR2_X1 U446 ( .A(G50GAT), .B(KEYINPUT78), .Z(n434) );
  XNOR2_X1 U447 ( .A(n393), .B(n434), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n561) );
  NAND2_X1 U450 ( .A1(n398), .A2(n561), .ZN(n399) );
  XNOR2_X1 U451 ( .A(KEYINPUT47), .B(n399), .ZN(n405) );
  XNOR2_X1 U452 ( .A(KEYINPUT36), .B(n561), .ZN(n573) );
  NOR2_X1 U453 ( .A1(n573), .A2(n558), .ZN(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n403) );
  NAND2_X1 U456 ( .A1(n569), .A2(n565), .ZN(n402) );
  NOR2_X1 U457 ( .A1(n403), .A2(n402), .ZN(n404) );
  NOR2_X1 U458 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U459 ( .A(KEYINPUT48), .B(n406), .ZN(n517) );
  NOR2_X1 U460 ( .A1(n452), .A2(n517), .ZN(n407) );
  XOR2_X1 U461 ( .A(n407), .B(KEYINPUT54), .Z(n408) );
  NOR2_X1 U462 ( .A1(n504), .A2(n408), .ZN(n548) );
  XOR2_X1 U463 ( .A(G99GAT), .B(G134GAT), .Z(n410) );
  XNOR2_X1 U464 ( .A(G43GAT), .B(G190GAT), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U467 ( .A1(G227GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U469 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n416) );
  XNOR2_X1 U470 ( .A(G176GAT), .B(KEYINPUT86), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U472 ( .A(n418), .B(n417), .Z(n424) );
  XOR2_X1 U473 ( .A(G71GAT), .B(G127GAT), .Z(n420) );
  XNOR2_X1 U474 ( .A(G15GAT), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U476 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n550) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U479 ( .A(G22GAT), .B(G204GAT), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n439) );
  XOR2_X1 U481 ( .A(KEYINPUT91), .B(G148GAT), .Z(n428) );
  XNOR2_X1 U482 ( .A(KEYINPUT88), .B(KEYINPUT90), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U484 ( .A(n430), .B(n429), .Z(n437) );
  XOR2_X1 U485 ( .A(KEYINPUT24), .B(n431), .Z(n433) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n547) );
  NOR2_X1 U492 ( .A1(n550), .A2(n547), .ZN(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT26), .B(n442), .Z(n443) );
  XNOR2_X1 U494 ( .A(KEYINPUT97), .B(n443), .ZN(n535) );
  AND2_X1 U495 ( .A1(n548), .A2(n535), .ZN(n444) );
  NOR2_X1 U496 ( .A1(n558), .A2(n572), .ZN(n447) );
  NAND2_X1 U497 ( .A1(n561), .A2(n448), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT16), .B(n449), .Z(n463) );
  INV_X1 U499 ( .A(n452), .ZN(n506) );
  NAND2_X1 U500 ( .A1(n550), .A2(n506), .ZN(n450) );
  NAND2_X1 U501 ( .A1(n547), .A2(n450), .ZN(n451) );
  XOR2_X1 U502 ( .A(KEYINPUT25), .B(n451), .Z(n454) );
  XOR2_X1 U503 ( .A(n452), .B(KEYINPUT27), .Z(n457) );
  NAND2_X1 U504 ( .A1(n457), .A2(n535), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n454), .A2(n453), .ZN(n456) );
  NAND2_X1 U506 ( .A1(n456), .A2(n455), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n504), .A2(n457), .ZN(n516) );
  XNOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(n547), .ZN(n519) );
  NOR2_X1 U510 ( .A1(n516), .A2(n519), .ZN(n460) );
  INV_X1 U511 ( .A(n550), .ZN(n459) );
  NAND2_X1 U512 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n462), .A2(n461), .ZN(n475) );
  NAND2_X1 U514 ( .A1(n463), .A2(n475), .ZN(n492) );
  INV_X1 U515 ( .A(n565), .ZN(n491) );
  NAND2_X1 U516 ( .A1(n569), .A2(n491), .ZN(n478) );
  NOR2_X1 U517 ( .A1(n492), .A2(n478), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n464), .B(KEYINPUT98), .ZN(n473) );
  NAND2_X1 U519 ( .A1(n473), .A2(n504), .ZN(n468) );
  XOR2_X1 U520 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n466) );
  XNOR2_X1 U521 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U522 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(G1324GAT) );
  NAND2_X1 U524 ( .A1(n473), .A2(n506), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n471) );
  NAND2_X1 U527 ( .A1(n550), .A2(n473), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U529 ( .A(G15GAT), .B(n472), .Z(G1326GAT) );
  NAND2_X1 U530 ( .A1(n473), .A2(n519), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n481) );
  NAND2_X1 U533 ( .A1(n558), .A2(n475), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n476), .A2(n573), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(KEYINPUT37), .ZN(n503) );
  NOR2_X1 U536 ( .A1(n503), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT38), .B(n479), .ZN(n489) );
  NAND2_X1 U538 ( .A1(n504), .A2(n489), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G29GAT), .B(n482), .ZN(G1328GAT) );
  XOR2_X1 U541 ( .A(G36GAT), .B(KEYINPUT103), .Z(n484) );
  NAND2_X1 U542 ( .A1(n489), .A2(n506), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1329GAT) );
  XNOR2_X1 U544 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n486) );
  NAND2_X1 U546 ( .A1(n550), .A2(n489), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1330GAT) );
  NAND2_X1 U549 ( .A1(n489), .A2(n519), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(G50GAT), .ZN(G1331GAT) );
  OR2_X1 U551 ( .A1(n491), .A2(n553), .ZN(n502) );
  NOR2_X1 U552 ( .A1(n502), .A2(n492), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT106), .ZN(n499) );
  NAND2_X1 U554 ( .A1(n504), .A2(n499), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT42), .B(n494), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(n495), .ZN(G1332GAT) );
  XOR2_X1 U557 ( .A(G64GAT), .B(KEYINPUT107), .Z(n497) );
  NAND2_X1 U558 ( .A1(n499), .A2(n506), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n550), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U562 ( .A(G78GAT), .B(KEYINPUT43), .Z(n501) );
  NAND2_X1 U563 ( .A1(n499), .A2(n519), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1335GAT) );
  NOR2_X1 U565 ( .A1(n503), .A2(n502), .ZN(n511) );
  NAND2_X1 U566 ( .A1(n504), .A2(n511), .ZN(n505) );
  XNOR2_X1 U567 ( .A(G85GAT), .B(n505), .ZN(G1336GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n511), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(KEYINPUT108), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G92GAT), .B(n508), .ZN(G1337GAT) );
  XOR2_X1 U571 ( .A(G99GAT), .B(KEYINPUT109), .Z(n510) );
  NAND2_X1 U572 ( .A1(n511), .A2(n550), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1338GAT) );
  XNOR2_X1 U574 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n515) );
  XOR2_X1 U575 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n513) );
  NAND2_X1 U576 ( .A1(n511), .A2(n519), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1339GAT) );
  NOR2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n550), .A2(n534), .ZN(n518) );
  NOR2_X1 U581 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(KEYINPUT113), .B(n520), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n565), .A2(n530), .ZN(n522) );
  XNOR2_X1 U584 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  NOR2_X1 U587 ( .A1(n553), .A2(n530), .ZN(n525) );
  XNOR2_X1 U588 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G120GAT), .B(n526), .ZN(G1341GAT) );
  NOR2_X1 U591 ( .A1(n558), .A2(n530), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(n529), .ZN(G1342GAT) );
  NOR2_X1 U595 ( .A1(n561), .A2(n530), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT118), .B(KEYINPUT51), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G134GAT), .B(n533), .ZN(G1343GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(n536), .Z(n545) );
  NOR2_X1 U601 ( .A1(n565), .A2(n545), .ZN(n537) );
  XOR2_X1 U602 ( .A(G141GAT), .B(n537), .Z(n538) );
  XNOR2_X1 U603 ( .A(KEYINPUT120), .B(n538), .ZN(G1344GAT) );
  NOR2_X1 U604 ( .A1(n553), .A2(n545), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n540) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT121), .B(n541), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U610 ( .A1(n558), .A2(n545), .ZN(n544) );
  XOR2_X1 U611 ( .A(G155GAT), .B(n544), .Z(G1346GAT) );
  NOR2_X1 U612 ( .A1(n561), .A2(n545), .ZN(n546) );
  XOR2_X1 U613 ( .A(G162GAT), .B(n546), .Z(G1347GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT55), .B(n549), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n551), .A2(n550), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n560), .A2(n565), .ZN(n552) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U619 ( .A1(n560), .A2(n553), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n558), .A2(n560), .ZN(n559) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n559), .Z(G1350GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U627 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G190GAT), .B(n564), .Z(G1351GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n572), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n572), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(n576), .ZN(G1355GAT) );
endmodule

