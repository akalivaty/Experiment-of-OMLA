//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XOR2_X1   g000(.A(G116), .B(G119), .Z(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(new_n198), .B2(G146), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n196), .A2(KEYINPUT64), .A3(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n197), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n201), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G137), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  AOI21_X1  g030(.A(G131), .B1(new_n210), .B2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n217), .A3(new_n213), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n195), .B1(new_n208), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n211), .A2(new_n217), .A3(new_n213), .ZN(new_n221));
  INV_X1    g035(.A(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n212), .A2(G134), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(new_n214), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n197), .A3(new_n199), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n198), .A2(G146), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT64), .B1(new_n196), .B2(G143), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n202), .A2(new_n198), .A3(G146), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n226), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT28), .B1(new_n220), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n237), .B1(new_n221), .B2(new_n224), .ZN(new_n238));
  INV_X1    g052(.A(new_n224), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(new_n218), .A3(KEYINPUT65), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n208), .A2(new_n219), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n195), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n227), .A2(new_n197), .A3(new_n199), .ZN(new_n245));
  INV_X1    g059(.A(new_n233), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(new_n205), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n218), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n225), .A2(new_n234), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n220), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n236), .B1(new_n253), .B2(KEYINPUT28), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT27), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT30), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n262), .B1(new_n243), .B2(new_n263), .ZN(new_n264));
  AOI211_X1 g078(.A(KEYINPUT66), .B(KEYINPUT30), .C1(new_n241), .C2(new_n242), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n249), .A2(KEYINPUT30), .A3(new_n242), .A4(new_n251), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n195), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT68), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n267), .A2(new_n195), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n270), .B(new_n271), .C1(new_n265), .C2(new_n264), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n252), .B2(new_n259), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT31), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n279), .B(new_n276), .C1(new_n269), .C2(new_n272), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n261), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT29), .B1(new_n254), .B2(new_n259), .ZN(new_n286));
  INV_X1    g100(.A(new_n252), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n269), .B2(new_n272), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n288), .B2(new_n259), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n249), .A2(new_n242), .A3(new_n251), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n195), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n252), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n236), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n281), .A2(new_n285), .B1(new_n296), .B2(G472), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n273), .A2(new_n277), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n279), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n276), .B1(new_n269), .B2(new_n272), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT31), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n260), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n284), .B1(new_n302), .B2(new_n283), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT16), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n307), .A2(KEYINPUT16), .A3(G140), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n196), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n310), .A3(G146), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G128), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(G128), .ZN(new_n318));
  OAI211_X1 g132(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(KEYINPUT23), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  XNOR2_X1  g134(.A(G119), .B(G128), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n314), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT70), .B(G110), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n319), .A2(new_n324), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n196), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n313), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G137), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n329), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT71), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n336));
  AOI21_X1  g150(.A(G902), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT71), .A3(KEYINPUT25), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n334), .B(new_n337), .C1(new_n335), .C2(new_n336), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  INV_X1    g155(.A(G902), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(G234), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n334), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n344), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT72), .Z(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n331), .A2(G227), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G107), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n359), .A2(KEYINPUT3), .A3(G104), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT3), .B1(new_n359), .B2(G104), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(G101), .ZN(new_n364));
  INV_X1    g178(.A(G101), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n359), .A2(G104), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n359), .A2(KEYINPUT3), .A3(G104), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n370), .B2(new_n358), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n365), .B(new_n358), .C1(new_n360), .C2(new_n361), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n208), .B(new_n364), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT73), .B1(new_n359), .B2(G104), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n357), .A3(G107), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n377), .A3(new_n366), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G101), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n372), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G143), .B(G146), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n228), .B1(new_n233), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n379), .A3(new_n372), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n380), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n219), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT75), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n389), .A3(new_n219), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n219), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n374), .A2(new_n392), .A3(new_n385), .A4(new_n380), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n356), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n379), .A2(new_n372), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n383), .B1(new_n395), .B2(new_n234), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n392), .A2(KEYINPUT74), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT12), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n393), .A2(new_n356), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n353), .B(new_n342), .C1(new_n394), .C2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n386), .A2(new_n389), .A3(new_n219), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n389), .B1(new_n386), .B2(new_n219), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n393), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n356), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n404), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT76), .A3(new_n353), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n403), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n391), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n393), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n411), .B1(new_n402), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n353), .B1(new_n421), .B2(new_n342), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n352), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G210), .B1(G237), .B2(G902), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT83), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n373), .A2(new_n371), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n364), .A2(new_n195), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT77), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n362), .A2(G101), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(KEYINPUT4), .A3(new_n372), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT77), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n195), .A4(new_n364), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n315), .A3(G116), .ZN(new_n435));
  OAI211_X1 g249(.A(G113), .B(new_n435), .C1(new_n187), .C2(new_n434), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n395), .A2(new_n194), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n429), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT78), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n429), .A2(new_n440), .A3(new_n433), .A4(new_n437), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(KEYINPUT6), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n307), .B(new_n228), .C1(new_n232), .C2(new_n233), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT79), .B(new_n447), .C1(new_n208), .C2(new_n307), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT79), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n232), .A2(new_n206), .A3(new_n200), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n449), .B(G125), .C1(new_n450), .C2(new_n201), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT80), .B(G224), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n331), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT81), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n452), .B(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n444), .A2(new_n446), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n448), .B2(new_n451), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT82), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n440), .B(KEYINPUT8), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n436), .A2(new_n194), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n379), .A2(new_n372), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n437), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n448), .A2(new_n458), .A3(new_n451), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n443), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n342), .B1(new_n461), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n426), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n459), .B(KEYINPUT82), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n443), .A2(new_n467), .A3(new_n468), .ZN(new_n473));
  AOI21_X1  g287(.A(G902), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n444), .A2(new_n446), .A3(new_n456), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(new_n475), .A3(new_n425), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G214), .B1(G237), .B2(G902), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n331), .A2(G952), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n477), .A2(new_n478), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(G475), .A2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT89), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n491));
  INV_X1    g305(.A(G237), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n331), .A3(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n198), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n491), .B1(new_n496), .B2(G131), .ZN(new_n497));
  AOI211_X1 g311(.A(KEYINPUT86), .B(new_n222), .C1(new_n494), .C2(new_n495), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT17), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n500));
  AOI21_X1  g314(.A(G143), .B1(new_n255), .B2(G214), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT86), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n496), .A2(new_n491), .A3(G131), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n222), .A3(new_n495), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n314), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n357), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n500), .A2(new_n501), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT18), .A4(G131), .ZN(new_n514));
  NAND2_X1  g328(.A1(KEYINPUT18), .A2(G131), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n496), .B2(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n196), .B1(new_n306), .B2(new_n308), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT84), .B1(new_n519), .B2(new_n327), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n306), .A2(new_n308), .A3(new_n196), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n521), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n509), .A2(new_n511), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n309), .A2(G146), .A3(new_n310), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n306), .A2(new_n308), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT19), .ZN(new_n532));
  AOI21_X1  g346(.A(G146), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n528), .B1(new_n533), .B2(KEYINPUT87), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n326), .A2(KEYINPUT19), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n196), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n527), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n511), .B1(new_n540), .B2(new_n525), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n526), .B1(new_n541), .B2(KEYINPUT88), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n543), .B(new_n511), .C1(new_n540), .C2(new_n525), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n490), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT20), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n490), .C1(new_n542), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G122), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n550), .A2(G116), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(G116), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(new_n359), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(G128), .A3(new_n198), .ZN(new_n556));
  XOR2_X1   g370(.A(G128), .B(G143), .Z(new_n557));
  OAI211_X1 g371(.A(new_n556), .B(G134), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n554), .B(new_n558), .C1(G134), .C2(new_n557), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT14), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n551), .B1(new_n560), .B2(new_n552), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n560), .B2(new_n552), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G107), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n557), .B(G134), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n553), .A2(new_n359), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n350), .A2(new_n341), .A3(G953), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n559), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n342), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n572));
  NOR2_X1   g386(.A1(KEYINPUT92), .A2(KEYINPUT15), .ZN(new_n573));
  OAI21_X1  g387(.A(G478), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n571), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n503), .A2(new_n504), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n314), .B1(new_n576), .B2(KEYINPUT17), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n577), .A2(new_n507), .B1(new_n517), .B2(new_n524), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT90), .B1(new_n578), .B2(new_n511), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n509), .A2(new_n525), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  INV_X1    g395(.A(new_n511), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n579), .A2(new_n583), .B1(new_n511), .B2(new_n578), .ZN(new_n584));
  OAI21_X1  g398(.A(G475), .B1(new_n584), .B2(G902), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n549), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n488), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n304), .A2(new_n349), .A3(new_n424), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT93), .B(G101), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(G3));
  NOR2_X1   g404(.A1(new_n302), .A2(new_n283), .ZN(new_n591));
  INV_X1    g405(.A(G472), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n281), .B2(new_n342), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n349), .A3(new_n424), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n549), .A2(new_n585), .ZN(new_n596));
  INV_X1    g410(.A(new_n570), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n597), .B2(new_n568), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT95), .B1(new_n598), .B2(G478), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n571), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT94), .B1(new_n569), .B2(new_n570), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n559), .B2(new_n566), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n601), .A2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n603), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n596), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n478), .ZN(new_n614));
  INV_X1    g428(.A(new_n425), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n457), .B2(new_n470), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n616), .B2(new_n476), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n487), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n595), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT34), .B(G104), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  XNOR2_X1  g435(.A(new_n598), .B(new_n574), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n549), .A2(new_n622), .A3(new_n585), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n595), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n333), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT96), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT97), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT96), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n628), .B(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n329), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n630), .A2(new_n634), .A3(new_n323), .A4(new_n328), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n346), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n344), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n594), .A2(new_n587), .A3(new_n424), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  AOI21_X1  g457(.A(KEYINPUT76), .B1(new_n414), .B2(new_n353), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n404), .B1(new_n411), .B2(new_n410), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n645), .A2(new_n406), .A3(G469), .A4(G902), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n423), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n352), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n474), .A2(new_n475), .A3(new_n425), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n425), .B1(new_n474), .B2(new_n475), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n478), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n481), .B1(G900), .B2(new_n483), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n549), .A2(new_n585), .A3(new_n622), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(KEYINPUT98), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n654), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n617), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n649), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n640), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n297), .B2(new_n303), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT99), .B(G128), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G30));
  INV_X1    g478(.A(new_n259), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n292), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n342), .B1(new_n667), .B2(new_n300), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  INV_X1    g483(.A(new_n285), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n669), .B1(new_n302), .B2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT32), .B1(new_n281), .B2(new_n282), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n477), .B(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n575), .B1(new_n549), .B2(new_n585), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(new_n478), .A3(new_n660), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n653), .B(KEYINPUT39), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n424), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT102), .B(G143), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G45));
  NAND3_X1  g499(.A1(new_n596), .A2(new_n612), .A3(new_n653), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n640), .B(new_n478), .C1(new_n650), .C2(new_n651), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n281), .A2(new_n285), .ZN(new_n689));
  INV_X1    g503(.A(new_n286), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT30), .B1(new_n241), .B2(new_n242), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n262), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n271), .B1(new_n692), .B2(new_n270), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n266), .A2(KEYINPUT68), .A3(new_n268), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n252), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n690), .B1(new_n695), .B2(new_n665), .ZN(new_n696));
  INV_X1    g510(.A(new_n295), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n424), .B(new_n688), .C1(new_n699), .C2(new_n672), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  OAI21_X1  g515(.A(G469), .B1(new_n645), .B2(G902), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n648), .B(new_n702), .C1(new_n644), .C2(new_n646), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n618), .A2(new_n613), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n304), .A2(new_n704), .A3(new_n349), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NOR2_X1   g522(.A1(new_n618), .A2(new_n623), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n304), .A2(new_n704), .A3(new_n349), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT103), .B(G116), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G18));
  NOR3_X1   g526(.A1(new_n703), .A2(new_n486), .A3(new_n652), .ZN(new_n713));
  INV_X1    g527(.A(new_n586), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n304), .A3(new_n714), .A4(new_n640), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  NAND2_X1  g530(.A1(new_n299), .A2(new_n301), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n293), .A2(KEYINPUT104), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n293), .A2(KEYINPUT104), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n665), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n283), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n593), .A2(new_n721), .A3(new_n348), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n676), .A3(new_n713), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G122), .ZN(G24));
  NOR3_X1   g538(.A1(new_n593), .A2(new_n721), .A3(new_n660), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n703), .A2(new_n652), .A3(new_n686), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  AOI21_X1  g542(.A(new_n422), .B1(new_n407), .B2(new_n415), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n471), .A2(new_n476), .A3(new_n478), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n729), .A2(new_n352), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n686), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n304), .A2(new_n349), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n348), .B1(new_n297), .B2(new_n303), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT42), .A3(new_n732), .A4(new_n731), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G131), .ZN(G33));
  AND4_X1   g553(.A1(new_n304), .A2(new_n349), .A3(new_n656), .A4(new_n731), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n210), .ZN(G36));
  XNOR2_X1  g555(.A(new_n604), .B(new_n607), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n742), .A2(new_n610), .B1(new_n599), .B2(new_n602), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n596), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n594), .A2(new_n660), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n748), .A2(KEYINPUT106), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n756), .B1(new_n421), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n353), .B1(new_n421), .B2(new_n757), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n418), .A2(KEYINPUT105), .A3(KEYINPUT45), .A4(new_n420), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n416), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n648), .A3(new_n679), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n730), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n754), .A2(new_n755), .A3(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  NOR4_X1   g585(.A1(new_n304), .A2(new_n349), .A3(new_n686), .A4(new_n730), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT108), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n767), .A2(new_n648), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n779));
  NOR2_X1   g593(.A1(G952), .A2(G953), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n746), .A2(new_n481), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n703), .A2(new_n730), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(G472), .B1(new_n302), .B2(G902), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n720), .B1(new_n278), .B2(new_n280), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(new_n282), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(new_n640), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n348), .A2(new_n481), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n673), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n743), .A2(new_n585), .A3(new_n549), .ZN(new_n790));
  OAI22_X1  g604(.A1(new_n783), .A2(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n675), .A2(new_n704), .A3(new_n614), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n781), .A2(new_n722), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(KEYINPUT113), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n791), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n416), .A2(new_n702), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n648), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT112), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n776), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n801), .B2(new_n776), .ZN(new_n803));
  INV_X1    g617(.A(new_n730), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n781), .A2(new_n722), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n736), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n783), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n781), .A2(new_n617), .A3(new_n704), .A4(new_n722), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n811), .B(new_n479), .C1(new_n613), .C2(new_n789), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n791), .A2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n795), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n805), .B1(new_n776), .B2(new_n800), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n817), .A2(new_n821), .A3(new_n795), .A4(new_n819), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n816), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n807), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n344), .A2(new_n639), .A3(new_n653), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n617), .A2(new_n676), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n829), .B(new_n424), .C1(new_n671), .C2(new_n672), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n700), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n659), .A2(new_n661), .B1(new_n725), .B2(new_n726), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT111), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT111), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n657), .B1(new_n656), .B2(new_n617), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n652), .A2(new_n654), .A3(KEYINPUT98), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n424), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n640), .B1(new_n699), .B2(new_n672), .ZN(new_n838));
  INV_X1    g652(.A(new_n702), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n407), .B2(new_n415), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n732), .A2(new_n840), .A3(new_n648), .A4(new_n617), .ZN(new_n841));
  OAI22_X1  g655(.A1(new_n837), .A2(new_n838), .B1(new_n787), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n700), .A2(new_n830), .A3(KEYINPUT52), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n834), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n700), .A2(new_n830), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n833), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n488), .B1(new_n613), .B2(new_n623), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n594), .A2(new_n849), .A3(new_n349), .A4(new_n424), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n710), .A2(new_n715), .A3(new_n723), .A4(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n588), .A2(new_n706), .A3(new_n641), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n640), .A2(new_n653), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n647), .A2(new_n804), .A3(new_n648), .A4(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n714), .B1(new_n699), .B2(new_n672), .ZN(new_n855));
  INV_X1    g669(.A(new_n613), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n784), .A2(new_n856), .A3(new_n786), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n740), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n851), .A2(new_n738), .A3(new_n852), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n827), .B1(new_n848), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n715), .A2(new_n710), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n723), .A2(new_n850), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n852), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n738), .A2(new_n859), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n847), .B1(new_n842), .B2(new_n843), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n826), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT53), .B1(new_n848), .B2(new_n860), .ZN(new_n870));
  INV_X1    g684(.A(new_n864), .ZN(new_n871));
  INV_X1    g685(.A(new_n865), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n872), .A3(new_n867), .A4(new_n827), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT54), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n780), .B1(new_n825), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT109), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n348), .A2(new_n352), .A3(new_n614), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n675), .A2(new_n744), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n878), .A2(new_n673), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT110), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n779), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n883), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n807), .A2(new_n824), .A3(new_n869), .A4(new_n874), .ZN(new_n886));
  OAI211_X1 g700(.A(KEYINPUT116), .B(new_n885), .C1(new_n886), .C2(new_n780), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(G75));
  NAND3_X1  g702(.A1(new_n833), .A2(new_n844), .A3(new_n847), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n827), .B1(new_n866), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n662), .A2(new_n727), .A3(new_n700), .A4(new_n830), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n891), .A2(new_n845), .B1(new_n831), .B2(new_n832), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n860), .A2(new_n892), .A3(KEYINPUT53), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G902), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n444), .A2(new_n446), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n456), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n331), .A2(G952), .ZN(new_n902));
  NOR2_X1   g716(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n903));
  AND2_X1   g717(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n896), .B2(new_n426), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n901), .A2(new_n902), .A3(new_n906), .ZN(G51));
  OAI21_X1  g721(.A(new_n826), .B1(new_n890), .B2(new_n893), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n874), .A2(KEYINPUT118), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n873), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n762), .B(KEYINPUT57), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n394), .B2(new_n404), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n895), .A2(new_n761), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n902), .B1(new_n916), .B2(new_n917), .ZN(G54));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n870), .A2(G902), .A3(new_n873), .A4(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n542), .A2(new_n544), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n919), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n902), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n922), .A2(KEYINPUT119), .A3(new_n924), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT120), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n866), .B2(new_n889), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n860), .A2(new_n892), .A3(new_n827), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n935), .B2(new_n908), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT121), .B1(new_n936), .B2(new_n742), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n609), .A2(new_n932), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n912), .B1(new_n874), .B2(KEYINPUT118), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n909), .B(KEYINPUT54), .C1(new_n870), .C2(new_n873), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n932), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n869), .B2(new_n874), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n609), .ZN(new_n945));
  INV_X1    g759(.A(new_n902), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n937), .A2(new_n941), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n902), .B1(new_n913), .B2(new_n938), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(KEYINPUT122), .A3(new_n937), .A4(new_n945), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n894), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n902), .B1(new_n955), .B2(new_n345), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n638), .B(KEYINPUT123), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n956), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(G66));
  INV_X1    g774(.A(new_n453), .ZN(new_n961));
  OAI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n485), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n871), .B2(G953), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n898), .B1(G898), .B2(new_n331), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT124), .Z(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT125), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n963), .B(new_n966), .ZN(G69));
  NAND2_X1  g781(.A1(new_n692), .A2(new_n267), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT126), .Z(new_n969));
  NOR2_X1   g783(.A1(new_n535), .A2(new_n536), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n331), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n770), .A2(new_n777), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n730), .B1(new_n613), .B2(new_n623), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n680), .A2(new_n736), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n832), .A2(new_n700), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n683), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT62), .Z(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n740), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n736), .A2(new_n617), .A3(new_n676), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n984), .A2(new_n768), .ZN(new_n985));
  AND4_X1   g799(.A1(new_n738), .A2(new_n979), .A3(new_n983), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n974), .A2(new_n331), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n972), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n982), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n988), .ZN(new_n992));
  NAND2_X1  g806(.A1(G227), .A2(G900), .ZN(new_n993));
  AND4_X1   g807(.A1(G953), .A2(new_n992), .A3(new_n993), .A4(new_n971), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n991), .A2(new_n994), .ZN(G72));
  NAND4_X1  g809(.A1(new_n974), .A2(new_n871), .A3(new_n981), .A4(new_n976), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  AOI211_X1 g812(.A(new_n665), .B(new_n288), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n288), .A2(new_n665), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n974), .A2(new_n871), .A3(new_n986), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n998), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n288), .A2(new_n259), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n998), .B1(new_n1004), .B2(new_n300), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n861), .B2(new_n868), .ZN(new_n1006));
  NOR4_X1   g820(.A1(new_n999), .A2(new_n1003), .A3(new_n902), .A4(new_n1006), .ZN(G57));
endmodule


