//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n188), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n191));
  XNOR2_X1  g005(.A(G143), .B(G146), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT82), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n190), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n193), .A2(new_n195), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT3), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT79), .A2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT79), .A2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n208), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(G104), .B2(G107), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n206), .A2(new_n207), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT83), .B1(new_n203), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n215), .A2(new_n218), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT83), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n193), .A2(new_n195), .A3(new_n202), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT10), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n215), .A2(KEYINPUT84), .A3(new_n218), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n196), .A2(G146), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n189), .B2(G143), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n196), .A2(KEYINPUT65), .A3(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n195), .B1(new_n235), .B2(new_n191), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n196), .A2(KEYINPUT65), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n196), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n190), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n198), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n195), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n238), .A2(new_n243), .A3(KEYINPUT10), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n225), .A2(new_n226), .B1(new_n230), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT11), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT67), .A2(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT67), .A2(G134), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(G137), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G137), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G134), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n248), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT11), .B1(new_n253), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(G131), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT67), .A2(G134), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT67), .A2(G134), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n246), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(new_n251), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n259), .B2(G137), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n256), .B(new_n260), .C1(new_n262), .C2(new_n246), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT81), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n201), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT66), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT0), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n188), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n241), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n188), .ZN(new_n276));
  AND3_X1   g090(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(new_n235), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n268), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT79), .A2(G107), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT79), .A2(G107), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n212), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G107), .B1(new_n204), .B2(KEYINPUT3), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(new_n205), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n282), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n208), .A2(new_n213), .A3(KEYINPUT80), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(G101), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n215), .A2(KEYINPUT4), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n208), .A2(new_n213), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n214), .B1(new_n294), .B2(new_n282), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n293), .B1(new_n295), .B2(new_n290), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n266), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(G101), .A3(new_n290), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT4), .A3(new_n215), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT81), .A3(new_n281), .A4(new_n291), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n245), .A2(new_n265), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n244), .A2(new_n230), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n226), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n301), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n265), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n245), .A2(KEYINPUT87), .A3(new_n301), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n303), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(G110), .B(G140), .ZN(new_n313));
  INV_X1    g127(.A(G227), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G953), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n313), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n187), .B1(new_n312), .B2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n297), .A2(new_n300), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n304), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n309), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n264), .A3(new_n311), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n302), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT88), .A3(new_n316), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n302), .A2(new_n317), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT85), .B1(new_n221), .B2(new_n236), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n219), .A2(new_n327), .A3(new_n242), .A4(new_n195), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n326), .B(new_n328), .C1(new_n305), .C2(new_n306), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT12), .A3(new_n264), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n305), .A2(new_n306), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n328), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n264), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n325), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n318), .A2(new_n324), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G469), .ZN(new_n339));
  INV_X1    g153(.A(G902), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n339), .A2(new_n340), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n325), .B1(new_n310), .B2(new_n311), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n329), .A2(KEYINPUT12), .A3(new_n264), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n329), .B2(new_n264), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n302), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT86), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n302), .B(new_n348), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n350), .B2(new_n316), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n342), .B1(new_n351), .B2(G469), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  INV_X1    g168(.A(G953), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G214), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n196), .ZN(new_n357));
  NOR2_X1   g171(.A1(G237), .A2(G953), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(G143), .A3(G214), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT18), .A2(G131), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G125), .ZN(new_n364));
  INV_X1    g178(.A(G125), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G140), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G146), .ZN(new_n368));
  XNOR2_X1  g182(.A(G125), .B(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n189), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n371), .A2(KEYINPUT94), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(KEYINPUT94), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n362), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT95), .B(G104), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n256), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n360), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n357), .A2(new_n256), .A3(new_n359), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n364), .A2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT76), .B1(new_n369), .B2(KEYINPUT16), .ZN(new_n385));
  OAI211_X1 g199(.A(G146), .B(new_n384), .C1(new_n385), .C2(new_n382), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n367), .B(KEYINPUT19), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n381), .B(new_n386), .C1(G146), .C2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n374), .A2(new_n377), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n377), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT16), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n383), .B1(new_n367), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(KEYINPUT16), .B2(new_n364), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n394), .A2(KEYINPUT77), .A3(G146), .A4(new_n384), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n385), .A2(new_n382), .ZN(new_n398));
  INV_X1    g212(.A(new_n384), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n189), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n378), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n381), .B2(KEYINPUT17), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n374), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n390), .B1(new_n391), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n391), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n409), .A2(new_n389), .A3(new_n407), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n377), .A2(KEYINPUT96), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n340), .B1(new_n404), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(G475), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n196), .A2(G128), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n196), .A2(G128), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n259), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G122), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G116), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT70), .B(G116), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G122), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n217), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n425), .A2(new_n427), .A3(new_n206), .A4(new_n207), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT13), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n420), .B1(new_n418), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT98), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n435), .B(new_n420), .C1(new_n418), .C2(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n196), .A2(KEYINPUT13), .A3(G128), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT99), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(G134), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n438), .B2(G134), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n421), .B(new_n431), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n419), .A2(new_n420), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n253), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n430), .A2(new_n443), .B1(new_n421), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n425), .B1(KEYINPUT14), .B2(new_n427), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n427), .A2(KEYINPUT14), .ZN(new_n448));
  OAI21_X1  g262(.A(G107), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n446), .B(new_n449), .C1(new_n443), .C2(new_n430), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  INV_X1    g265(.A(G217), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n451), .A2(new_n452), .A3(G953), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n442), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n442), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n340), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G478), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT15), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n456), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n355), .A2(G952), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n460), .B1(G234), .B2(G237), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n340), .B(new_n355), .C1(G234), .C2(G237), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(G898), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n417), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT91), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n195), .B(new_n365), .C1(new_n235), .C2(new_n191), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT89), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n355), .A2(G224), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n471), .B(new_n475), .C1(new_n365), .C2(new_n281), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n469), .B(KEYINPUT89), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n281), .A2(new_n365), .ZN(new_n478));
  OAI22_X1  g292(.A1(new_n477), .A2(new_n478), .B1(new_n474), .B2(new_n473), .ZN(new_n479));
  XNOR2_X1  g293(.A(G110), .B(G122), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n480), .B(KEYINPUT8), .Z(new_n481));
  INV_X1    g295(.A(G119), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n482), .A2(G116), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n426), .B2(G119), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT5), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G113), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  XOR2_X1   g303(.A(KEYINPUT2), .B(G113), .Z(new_n490));
  AOI22_X1  g304(.A1(new_n485), .A2(new_n489), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n481), .B1(new_n491), .B2(new_n219), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n484), .A2(KEYINPUT90), .A3(KEYINPUT5), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n494), .A2(new_n495), .B1(new_n484), .B2(new_n490), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n496), .B2(new_n219), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n491), .A2(new_n228), .A3(new_n229), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n484), .B(new_n490), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n291), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n498), .B(new_n480), .C1(new_n500), .C2(new_n296), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n476), .A2(new_n479), .A3(new_n497), .A4(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n502), .A2(new_n340), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n498), .B1(new_n500), .B2(new_n296), .ZN(new_n504));
  INV_X1    g318(.A(new_n480), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n471), .B(new_n472), .C1(new_n365), .C2(new_n281), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n511), .A3(new_n505), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n468), .B1(new_n514), .B2(KEYINPUT92), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT92), .ZN(new_n516));
  INV_X1    g330(.A(new_n468), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n503), .A2(new_n513), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n503), .A2(new_n513), .A3(new_n467), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT92), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G214), .B1(G237), .B2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n353), .A2(new_n465), .A3(new_n466), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n264), .A2(new_n281), .ZN(new_n527));
  INV_X1    g341(.A(new_n499), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n259), .A2(G137), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n250), .A2(G134), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n238), .A2(new_n243), .A3(new_n531), .A4(new_n263), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT72), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n263), .A2(new_n531), .A3(new_n236), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n281), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n536), .B1(new_n541), .B2(new_n499), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n535), .B1(new_n542), .B2(new_n534), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n358), .A2(G210), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT27), .Z(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT26), .B(G101), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n545), .B(new_n546), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n539), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT69), .B1(new_n264), .B2(new_n281), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n499), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n533), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n543), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT30), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n527), .A2(KEYINPUT30), .A3(new_n532), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n499), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n547), .A3(new_n533), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT31), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT31), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n558), .A2(new_n561), .A3(new_n547), .A4(new_n533), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G472), .A2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT32), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n563), .A2(KEYINPUT32), .A3(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT74), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT73), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n558), .A2(new_n533), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n548), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n548), .B1(new_n543), .B2(new_n553), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n533), .A2(new_n534), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n527), .A2(new_n532), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n499), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n533), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n584), .B2(KEYINPUT28), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n548), .A2(new_n576), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n340), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n573), .B(G472), .C1(new_n579), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT72), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n542), .A2(new_n590), .A3(new_n534), .ZN(new_n591));
  INV_X1    g405(.A(new_n535), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n552), .B2(KEYINPUT28), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n547), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT29), .B1(new_n574), .B2(new_n548), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G472), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT73), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n570), .A2(new_n572), .B1(new_n589), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n452), .B1(G234), .B2(new_n340), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT24), .B(G110), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(KEYINPUT75), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n482), .A2(G128), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n188), .A2(G119), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n482), .A2(G128), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n604), .B(new_n608), .C1(new_n609), .C2(KEYINPUT23), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(G110), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n401), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT78), .B(G110), .Z(new_n614));
  OAI21_X1  g428(.A(new_n613), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n386), .A3(new_n370), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT22), .B(G137), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n355), .A2(G221), .A3(G234), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n617), .B(new_n618), .Z(new_n619));
  AND3_X1   g433(.A1(new_n612), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n612), .B2(new_n616), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT25), .B1(new_n622), .B2(new_n340), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT25), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n620), .A2(new_n621), .A3(new_n624), .A4(G902), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n600), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n600), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n622), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n526), .A2(new_n599), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(new_n214), .ZN(G3));
  INV_X1    g445(.A(new_n466), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n341), .B2(new_n352), .ZN(new_n633));
  INV_X1    g447(.A(new_n565), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n597), .B1(new_n563), .B2(new_n340), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(new_n635), .A3(new_n629), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n467), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n514), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n524), .B1(new_n639), .B2(new_n519), .ZN(new_n640));
  INV_X1    g454(.A(new_n464), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n457), .A2(new_n340), .ZN(new_n643));
  INV_X1    g457(.A(new_n456), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(new_n457), .ZN(new_n645));
  OR3_X1    g459(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT33), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT33), .B1(new_n454), .B2(new_n455), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(G478), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n417), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n642), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n637), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  AND3_X1   g469(.A1(new_n405), .A2(new_n411), .A3(new_n407), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n411), .B1(new_n405), .B2(new_n407), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n416), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n659), .A2(new_n640), .A3(new_n641), .A4(new_n459), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n637), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n612), .A2(new_n616), .ZN(new_n665));
  INV_X1    g479(.A(new_n619), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n665), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n627), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n626), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n465), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n671), .A2(new_n634), .A3(new_n635), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n633), .A2(new_n525), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  XOR2_X1   g489(.A(KEYINPUT101), .B(G900), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n462), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n461), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n416), .B(new_n679), .C1(new_n656), .C2(new_n657), .ZN(new_n680));
  INV_X1    g494(.A(new_n458), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n456), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n640), .A2(new_n683), .A3(new_n670), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n317), .B1(new_n322), .B2(new_n302), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n336), .B1(new_n686), .B2(KEYINPUT88), .ZN(new_n687));
  AOI211_X1 g501(.A(G469), .B(G902), .C1(new_n687), .C2(new_n318), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n351), .A2(G469), .ZN(new_n689));
  INV_X1    g503(.A(new_n342), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n466), .B(new_n685), .C1(new_n688), .C2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT102), .B1(new_n599), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n598), .A2(new_n589), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT32), .B1(new_n563), .B2(new_n564), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n571), .A2(new_n695), .A3(KEYINPUT74), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n569), .A2(new_n568), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n632), .B(new_n684), .C1(new_n341), .C2(new_n352), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n693), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(new_n679), .B(KEYINPUT39), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n633), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n570), .A2(new_n572), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n548), .B1(new_n558), .B2(new_n533), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n340), .B1(new_n584), .B2(new_n547), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n521), .B(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n412), .A2(new_n416), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n682), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n714), .A2(new_n524), .A3(new_n670), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n706), .A2(new_n707), .A3(new_n712), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  INV_X1    g534(.A(new_n633), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n599), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n650), .A2(new_n417), .A3(new_n679), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n724), .A2(new_n640), .A3(new_n670), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  AOI21_X1  g541(.A(new_n339), .B1(new_n338), .B2(new_n340), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n688), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n729), .B2(new_n466), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n338), .A2(new_n340), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n466), .A4(new_n341), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n730), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n629), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n698), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n732), .A2(new_n466), .A3(new_n341), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT105), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n733), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n735), .A2(new_n738), .A3(new_n652), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(KEYINPUT41), .B(G113), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G15));
  AND2_X1   g560(.A1(new_n735), .A2(new_n743), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n737), .A2(new_n660), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G116), .ZN(G18));
  NOR2_X1   g564(.A1(new_n730), .A2(new_n734), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n599), .A2(new_n671), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n640), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  OAI211_X1 g568(.A(new_n560), .B(new_n562), .C1(new_n547), .C2(new_n585), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n564), .B(KEYINPUT106), .Z(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n635), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n736), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n759), .A2(new_n642), .A3(new_n717), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n747), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G122), .ZN(G24));
  NAND2_X1  g576(.A1(new_n758), .A2(new_n670), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n723), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n741), .A2(new_n640), .A3(new_n733), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  AOI21_X1  g580(.A(new_n317), .B1(new_n347), .B2(new_n349), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n339), .A3(new_n343), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n342), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(new_n341), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n632), .A2(new_n524), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n521), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n772), .A2(new_n724), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT108), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n571), .A2(new_n695), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n694), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n777), .B1(new_n779), .B2(new_n736), .ZN(new_n780));
  AOI211_X1 g594(.A(KEYINPUT108), .B(new_n629), .C1(new_n694), .C2(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n775), .ZN(new_n783));
  INV_X1    g597(.A(new_n349), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n335), .A2(new_n330), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n348), .B1(new_n785), .B2(new_n302), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n316), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n343), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n769), .A3(G469), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n690), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n769), .B1(new_n351), .B2(G469), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n783), .B1(new_n792), .B2(new_n341), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(new_n698), .A3(new_n736), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n782), .A2(KEYINPUT42), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NAND4_X1  g611(.A1(new_n793), .A2(new_n698), .A3(new_n736), .A4(new_n683), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  NOR3_X1   g613(.A1(new_n649), .A2(new_n417), .A3(KEYINPUT43), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n715), .A2(KEYINPUT111), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n650), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n803), .B2(KEYINPUT43), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n634), .A2(new_n635), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n670), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT44), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n522), .A2(new_n523), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n806), .B2(new_n807), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT113), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n351), .A2(KEYINPUT45), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n351), .A2(KEYINPUT45), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(G469), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n342), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n341), .B1(new_n820), .B2(KEYINPUT46), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT46), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT110), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(KEYINPUT110), .A3(KEYINPUT46), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n466), .A3(new_n704), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n814), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(new_n250), .ZN(G39));
  XNOR2_X1  g644(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(new_n466), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n826), .A2(new_n632), .B1(new_n834), .B2(KEYINPUT47), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n698), .A2(new_n736), .A3(new_n723), .A4(new_n811), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g651(.A(KEYINPUT115), .B(G140), .Z(new_n838));
  XNOR2_X1  g652(.A(new_n837), .B(new_n838), .ZN(G42));
  NAND2_X1  g653(.A1(new_n833), .A2(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n729), .A2(new_n632), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n804), .A2(new_n461), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n843), .A2(new_n759), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n811), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n833), .A2(new_n835), .B1(new_n632), .B2(new_n729), .ZN(new_n848));
  INV_X1    g662(.A(new_n845), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n714), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n844), .A2(new_n523), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n751), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT50), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n730), .A2(new_n734), .A3(new_n811), .ZN(new_n855));
  INV_X1    g669(.A(new_n712), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n736), .A3(new_n461), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n715), .A2(new_n649), .ZN(new_n858));
  INV_X1    g672(.A(new_n843), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n763), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n854), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n846), .A2(new_n850), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT51), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n735), .B(new_n743), .C1(new_n748), .C2(new_n760), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n649), .A2(new_n417), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n682), .A2(new_n412), .A3(new_n416), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n641), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n522), .A3(new_n524), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n633), .A2(new_n636), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n673), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n630), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n866), .A2(new_n744), .A3(new_n753), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n793), .A2(new_n764), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n670), .A2(new_n682), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n811), .A2(new_n680), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n698), .A2(new_n633), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n798), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT116), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n798), .A2(new_n883), .A3(new_n877), .A4(new_n880), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n796), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n875), .A2(new_n876), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n796), .A2(new_n882), .A3(new_n884), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT117), .B1(new_n874), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n717), .A2(new_n670), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n640), .A2(new_n466), .A3(new_n679), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n712), .A2(new_n889), .A3(new_n772), .A4(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n702), .A2(new_n726), .A3(new_n765), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n693), .A2(new_n701), .B1(new_n722), .B2(new_n725), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(KEYINPUT52), .A3(new_n765), .A4(new_n891), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n886), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  XOR2_X1   g715(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n630), .A2(new_n872), .A3(new_n899), .ZN(new_n904));
  AND4_X1   g718(.A1(new_n744), .A2(new_n866), .A3(new_n753), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(new_n897), .A3(new_n885), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT118), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n866), .A2(new_n744), .A3(new_n753), .A4(new_n904), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n908), .A2(new_n887), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT118), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(new_n897), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n903), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n900), .A2(KEYINPUT54), .B1(new_n901), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(KEYINPUT51), .B(new_n862), .C1(new_n848), .C2(new_n849), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n780), .A2(new_n781), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n855), .A2(new_n915), .A3(new_n859), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT48), .Z(new_n917));
  NOR2_X1   g731(.A1(new_n857), .A2(new_n651), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n460), .B(KEYINPUT121), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n751), .A2(new_n640), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n844), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT122), .Z(new_n923));
  NAND4_X1  g737(.A1(new_n865), .A2(new_n913), .A3(new_n914), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(G952), .B2(G953), .ZN(new_n925));
  INV_X1    g739(.A(new_n729), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n926), .A2(KEYINPUT49), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n851), .A2(new_n629), .A3(new_n774), .A4(new_n803), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(KEYINPUT49), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(new_n856), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G75));
  NOR2_X1   g745(.A1(new_n355), .A2(G952), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n907), .A2(new_n911), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n340), .B1(new_n901), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(G210), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n507), .A2(new_n512), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(new_n510), .Z(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT55), .Z(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n932), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n938), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT56), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n935), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT124), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n945), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n948), .A3(new_n941), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(G51));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n910), .A2(new_n905), .A3(new_n885), .A4(new_n897), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n910), .B1(new_n909), .B2(new_n897), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n902), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n894), .A2(new_n896), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n874), .A2(new_n887), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n876), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT53), .B1(new_n957), .B2(new_n888), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n951), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n952), .A2(new_n953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n903), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n912), .A2(new_n901), .A3(KEYINPUT125), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n342), .B(KEYINPUT57), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n338), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n934), .A2(new_n818), .A3(new_n819), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n932), .B1(new_n966), .B2(new_n967), .ZN(G54));
  NAND3_X1  g782(.A1(new_n934), .A2(KEYINPUT58), .A3(G475), .ZN(new_n969));
  INV_X1    g783(.A(new_n405), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n932), .ZN(G60));
  AND2_X1   g787(.A1(new_n646), .A2(new_n647), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n643), .B(KEYINPUT59), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n913), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n932), .B1(new_n963), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g794(.A(KEYINPUT126), .B(new_n932), .C1(new_n963), .C2(new_n977), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G63));
  INV_X1    g796(.A(new_n932), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n901), .A2(new_n933), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n452), .A2(new_n340), .A3(KEYINPUT60), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT60), .B1(new_n452), .B2(new_n340), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n668), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n984), .A2(new_n985), .A3(new_n986), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n983), .B(new_n987), .C1(new_n988), .C2(new_n622), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT61), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(G66));
  INV_X1    g806(.A(new_n463), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n355), .B1(new_n993), .B2(G224), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n874), .B2(new_n355), .ZN(new_n995));
  INV_X1    g809(.A(G898), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n936), .B1(new_n996), .B2(G953), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n995), .B(new_n997), .ZN(G69));
  NAND2_X1  g812(.A1(new_n556), .A2(new_n557), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n387), .ZN(new_n1000));
  INV_X1    g814(.A(G900), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(new_n355), .ZN(new_n1002));
  INV_X1    g816(.A(new_n829), .ZN(new_n1003));
  AND4_X1   g817(.A1(new_n765), .A2(new_n796), .A3(new_n798), .A4(new_n895), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n915), .A2(new_n640), .A3(new_n716), .ZN(new_n1005));
  OR2_X1    g819(.A1(new_n828), .A2(new_n1005), .ZN(new_n1006));
  AND4_X1   g820(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n837), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1002), .B1(new_n1007), .B2(new_n355), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n867), .A2(new_n868), .ZN(new_n1009));
  OR4_X1    g823(.A1(new_n737), .A2(new_n705), .A3(new_n811), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n719), .A2(new_n895), .A3(new_n765), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT62), .Z(new_n1012));
  NAND4_X1  g826(.A1(new_n1003), .A2(new_n837), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1000), .B1(new_n1013), .B2(new_n355), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n355), .B1(G227), .B2(G900), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1008), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1015), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1013), .B2(new_n874), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n932), .B1(new_n1021), .B2(new_n709), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1003), .A2(new_n1006), .A3(new_n837), .A4(new_n1004), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1020), .B1(new_n1023), .B2(new_n874), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(new_n548), .A3(new_n533), .A4(new_n558), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n575), .A2(new_n559), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n900), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  AND3_X1   g841(.A1(new_n1022), .A2(new_n1025), .A3(new_n1027), .ZN(G57));
endmodule


