//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT65), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n471), .B1(new_n479), .B2(G2105), .ZN(G160));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  INV_X1    g056(.A(G136), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n469), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n474), .A2(G2105), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT66), .A3(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n474), .A2(new_n468), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n483), .A2(new_n485), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n467), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT4), .B1(new_n469), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n484), .A2(new_n499), .A3(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  NAND2_X1  g076(.A1(G75), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT67), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT68), .B(G88), .Z(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(new_n518), .B1(G50), .B2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n511), .B1(new_n516), .B2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(KEYINPUT67), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT67), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n515), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n529), .A2(new_n507), .A3(new_n513), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT70), .B(G89), .Z(new_n531));
  AOI21_X1  g106(.A(new_n525), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT69), .B1(new_n529), .B2(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT69), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n534), .B(new_n514), .C1(new_n510), .C2(new_n515), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G51), .A3(G543), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n507), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(new_n510), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n533), .A2(G52), .A3(G543), .A4(new_n535), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n530), .A2(G90), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT71), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT71), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n543), .B1(new_n547), .B2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n507), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n530), .A2(G81), .B1(new_n510), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n533), .A2(G43), .A3(G543), .A4(new_n535), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n533), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n503), .B1(new_n516), .B2(KEYINPUT69), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n565), .A2(new_n566), .A3(G53), .A4(new_n535), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n507), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n530), .A2(G91), .B1(G651), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  AND3_X1   g148(.A1(new_n544), .A2(new_n548), .A3(new_n545), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n548), .B1(new_n544), .B2(new_n545), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n542), .B1(new_n574), .B2(new_n575), .ZN(G301));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n537), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n532), .A2(KEYINPUT72), .A3(new_n536), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G286));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n512), .B1(new_n507), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n530), .B2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n565), .A2(new_n535), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(G288));
  AOI22_X1  g161(.A1(new_n518), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(new_n510), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n516), .A2(new_n587), .B1(new_n588), .B2(new_n589), .ZN(G305));
  NAND3_X1  g165(.A1(new_n565), .A2(G47), .A3(new_n535), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n518), .B(new_n514), .C1(new_n510), .C2(new_n515), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT73), .B(G85), .Z(new_n594));
  OAI221_X1 g169(.A(new_n591), .B1(new_n589), .B2(new_n592), .C1(new_n593), .C2(new_n594), .ZN(G290));
  NAND3_X1  g170(.A1(new_n530), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n593), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n565), .A2(G54), .A3(new_n535), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(new_n512), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G284));
  OAI21_X1  g182(.A(new_n606), .B1(G171), .B2(new_n605), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(G299), .B(KEYINPUT74), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  AND3_X1   g187(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g194(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n486), .A2(G123), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n484), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n468), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT75), .B(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(G2100), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n623), .A2(new_n630), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n645));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR3_X1    g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n645), .B1(new_n644), .B2(new_n647), .ZN(new_n649));
  INV_X1    g224(.A(G14), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n644), .B2(new_n647), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT78), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n654));
  NAND4_X1  g229(.A1(new_n648), .A2(new_n654), .A3(new_n649), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT79), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  INV_X1    g238(.A(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(new_n660), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n659), .B(KEYINPUT17), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n660), .A3(new_n664), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(KEYINPUT80), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(KEYINPUT80), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n663), .B(new_n667), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n677), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n675), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n683), .B2(new_n682), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT21), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n688), .B(new_n689), .Z(new_n690));
  OR2_X1    g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT22), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(new_n690), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n693), .B1(new_n691), .B2(new_n694), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G32), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n486), .A2(G129), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n484), .A2(G141), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n462), .A2(G105), .ZN(new_n702));
  NAND3_X1  g277(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT26), .Z(new_n704));
  NAND4_X1  g279(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n699), .B1(new_n706), .B2(new_n698), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT88), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT27), .B(G1996), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT89), .Z(new_n711));
  AND2_X1   g286(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n698), .A2(G27), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G164), .B2(new_n698), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2078), .ZN(new_n715));
  NOR2_X1   g290(.A1(G29), .A2(G33), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT86), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G139), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n462), .A2(G103), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT25), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(KEYINPUT25), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(G115), .A2(G2104), .ZN(new_n723));
  INV_X1    g298(.A(G127), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n474), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n722), .B1(G2105), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n717), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2072), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT30), .B(G28), .ZN(new_n729));
  OR2_X1    g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  NAND2_X1  g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n729), .A2(new_n698), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n628), .B2(new_n698), .ZN(new_n733));
  NOR4_X1   g308(.A1(new_n712), .A2(new_n715), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n556), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1341), .Z(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n698), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT87), .ZN(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g321(.A1(new_n711), .A2(new_n734), .A3(new_n738), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n698), .A2(G35), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n698), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G2090), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n698), .A2(G26), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n486), .A2(G128), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n484), .A2(G140), .ZN(new_n755));
  OR2_X1    g330(.A1(G104), .A2(G2105), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n756), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(new_n698), .ZN(new_n760));
  MUX2_X1   g335(.A(new_n753), .B(new_n760), .S(KEYINPUT28), .Z(new_n761));
  XOR2_X1   g336(.A(KEYINPUT85), .B(G2067), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G168), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT90), .B(G1966), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n745), .B2(new_n744), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n735), .A2(G5), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G171), .B2(new_n735), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT91), .B(G1961), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n735), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n613), .B2(new_n735), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1348), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n770), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT93), .B(KEYINPUT23), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n735), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G299), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n735), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT94), .B(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n772), .B2(new_n774), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n747), .A2(new_n764), .A3(new_n779), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n486), .A2(G119), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n484), .A2(G131), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n468), .A2(G107), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT83), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n735), .A2(G24), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G290), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G1986), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(G1986), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n797), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n735), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n735), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(G16), .A2(G23), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G288), .B2(new_n735), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT33), .B(G1976), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  MUX2_X1   g387(.A(G6), .B(G305), .S(G16), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n807), .A2(new_n811), .A3(new_n812), .A4(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n803), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(KEYINPUT84), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n803), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n816), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n826), .A3(new_n823), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n788), .B1(new_n825), .B2(new_n827), .ZN(G311));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n827), .ZN(new_n829));
  INV_X1    g404(.A(new_n788), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(G150));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n507), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n530), .A2(G93), .B1(new_n510), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n533), .A2(G55), .A3(G543), .A4(new_n535), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(KEYINPUT96), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n554), .A2(new_n555), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n835), .A2(new_n842), .A3(new_n836), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n556), .A2(new_n842), .A3(new_n836), .A4(new_n835), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G559), .B2(new_n613), .ZN(new_n847));
  AOI211_X1 g422(.A(new_n614), .B(new_n604), .C1(new_n844), .C2(new_n845), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  OR3_X1    g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n850), .B1(new_n847), .B2(new_n848), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(KEYINPUT39), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT97), .Z(new_n854));
  AOI21_X1  g429(.A(KEYINPUT39), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n854), .A2(KEYINPUT98), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(KEYINPUT98), .B1(new_n854), .B2(new_n856), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n839), .B1(new_n857), .B2(new_n858), .ZN(G145));
  AOI22_X1  g434(.A1(G130), .A2(new_n486), .B1(new_n484), .B2(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  OR3_X1    g438(.A1(new_n863), .A2(new_n468), .A3(G118), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(KEYINPUT101), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n468), .B2(G118), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n860), .B1(new_n862), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n758), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n621), .B(KEYINPUT102), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n726), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n793), .B(new_n705), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n484), .A2(G137), .B1(G101), .B2(new_n462), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n473), .A2(new_n476), .B1(G113), .B2(G2104), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n875), .B2(new_n468), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n490), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n873), .A2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  INV_X1    g457(.A(new_n869), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n878), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n628), .B(KEYINPUT99), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n498), .A2(new_n500), .ZN(new_n887));
  INV_X1    g462(.A(new_n496), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n886), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n881), .A2(new_n884), .A3(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g471(.A(G290), .B(G288), .Z(new_n897));
  XNOR2_X1  g472(.A(G303), .B(G305), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n897), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT42), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n604), .A2(new_n568), .A3(new_n572), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n604), .B1(new_n572), .B2(new_n568), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G299), .A2(new_n613), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n907), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(KEYINPUT103), .A3(KEYINPUT41), .A4(new_n907), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n846), .B(new_n616), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n911), .A2(new_n907), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n905), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n902), .A2(new_n904), .A3(new_n918), .A4(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n924), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n837), .A2(new_n605), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  AND2_X1   g505(.A1(new_n844), .A2(new_n845), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(G168), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n932), .A2(new_n933), .B1(G171), .B2(G286), .ZN(new_n934));
  NAND3_X1  g509(.A1(G301), .A2(KEYINPUT105), .A3(G168), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n933), .B1(G171), .B2(new_n537), .ZN(new_n937));
  NAND2_X1  g512(.A1(G286), .A2(G171), .ZN(new_n938));
  AND4_X1   g513(.A1(new_n931), .A2(new_n937), .A3(new_n935), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n919), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n935), .A3(new_n938), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n846), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n931), .A2(new_n937), .A3(new_n935), .A4(new_n938), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n914), .A3(new_n915), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n944), .A3(new_n900), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n893), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n910), .A2(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n912), .A2(KEYINPUT108), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n911), .A2(new_n949), .A3(KEYINPUT41), .A4(new_n907), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n919), .A2(new_n951), .A3(new_n906), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n943), .A3(new_n942), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n900), .B1(new_n954), .B2(new_n940), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n940), .A2(new_n944), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n901), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(KEYINPUT106), .A3(new_n893), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n900), .B1(new_n940), .B2(new_n944), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(G37), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n961), .A2(new_n964), .A3(new_n965), .A4(new_n945), .ZN(new_n966));
  OAI211_X1 g541(.A(KEYINPUT109), .B(KEYINPUT43), .C1(new_n946), .C2(new_n955), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n958), .A2(new_n966), .A3(KEYINPUT44), .A4(new_n967), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n946), .A2(new_n955), .A3(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n961), .A2(new_n964), .A3(new_n945), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n970), .B2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(KEYINPUT44), .B2(new_n971), .ZN(G397));
  XOR2_X1   g547(.A(KEYINPUT110), .B(G1384), .Z(new_n973));
  AOI21_X1  g548(.A(new_n973), .B1(new_n887), .B2(new_n888), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT111), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G164), .B2(new_n973), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n876), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n975), .A2(new_n977), .A3(new_n978), .A4(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(KEYINPUT112), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n706), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n983), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n758), .B(G2067), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n793), .A2(new_n796), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n981), .A2(G1996), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n706), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n759), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n992), .A2(new_n994), .B1(new_n983), .B2(new_n982), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n793), .A2(new_n796), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n986), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n988), .A2(new_n991), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT48), .Z(new_n1000));
  AND4_X1   g575(.A1(new_n997), .A2(new_n998), .A3(new_n985), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT127), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n990), .B(KEYINPUT46), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n984), .ZN(new_n1005));
  AND4_X1   g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n988), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n984), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n1007), .B2(new_n988), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT47), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1004), .A2(new_n1005), .A3(new_n988), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT127), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1007), .A2(new_n1002), .A3(new_n988), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n995), .B(new_n1001), .C1(new_n1009), .C2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g590(.A(G1976), .B(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n1016));
  NAND2_X1  g591(.A1(G160), .A2(G40), .ZN(new_n1017));
  AOI21_X1  g592(.A(G1384), .B1(new_n887), .B2(new_n888), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(G8), .B(new_n1016), .C1(new_n1017), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT52), .ZN(new_n1021));
  AND2_X1   g596(.A1(G305), .A2(G1981), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G305), .A2(G1981), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n980), .A2(new_n1018), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(G8), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1026), .A2(new_n1030), .A3(G8), .A4(new_n1016), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1021), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n974), .A2(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n978), .B1(G164), .B2(G1384), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n980), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n806), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(G1384), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n889), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1037), .A2(new_n1040), .A3(new_n980), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n1046));
  OAI22_X1  g621(.A1(G166), .A2(new_n1045), .B1(KEYINPUT114), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(KEYINPUT114), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1032), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1037), .A2(new_n1040), .A3(new_n980), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT113), .A3(new_n1041), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1042), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1055), .A3(new_n1036), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(G8), .A3(new_n1049), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1018), .A2(KEYINPUT45), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n980), .A3(new_n1034), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1052), .A2(new_n745), .B1(new_n1059), .B2(new_n768), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1060), .A2(new_n1045), .A3(G286), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1051), .A2(new_n1057), .A3(KEYINPUT116), .A4(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1051), .A2(new_n1057), .A3(new_n1061), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1057), .A2(new_n1061), .A3(KEYINPUT63), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1032), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1054), .A2(new_n1042), .B1(new_n1035), .B2(new_n806), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1045), .B1(new_n1070), .B2(new_n1053), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1069), .B1(new_n1071), .B2(new_n1049), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1068), .B1(KEYINPUT118), .B2(new_n1072), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1072), .A2(KEYINPUT118), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1064), .A2(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n537), .A2(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n1076), .B(KEYINPUT51), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1058), .A2(new_n980), .A3(new_n1034), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1037), .A2(new_n1040), .A3(new_n980), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1080), .A2(new_n767), .B1(G2084), .B2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(G8), .B(new_n1079), .C1(new_n1082), .C2(new_n537), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1078), .A2(KEYINPUT51), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1077), .B(new_n1084), .C1(new_n1060), .C2(new_n1045), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1077), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1082), .A2(new_n1086), .B1(new_n1076), .B2(KEYINPUT51), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT62), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1033), .A2(new_n1034), .A3(new_n1093), .A4(new_n980), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  INV_X1    g670(.A(G1961), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1094), .A2(new_n1095), .B1(new_n1081), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n1093), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .A4(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(G288), .A2(G1976), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1028), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(G8), .B(new_n1026), .C1(new_n1102), .C2(new_n1023), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1057), .B2(new_n1032), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT115), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1103), .B(new_n1106), .C1(new_n1057), .C2(new_n1032), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1100), .A2(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(G171), .B(KEYINPUT54), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n975), .A2(new_n978), .A3(new_n977), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n468), .B1(new_n479), .B2(KEYINPUT126), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(KEYINPUT126), .B2(new_n479), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n471), .A2(new_n1095), .A3(new_n979), .A4(G2078), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1112), .A2(new_n1033), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1097), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1111), .B1(new_n1110), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(new_n1088), .A3(new_n1057), .A4(new_n1051), .ZN(new_n1119));
  INV_X1    g694(.A(G1956), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1081), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(G2072), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1033), .A2(new_n1034), .A3(new_n980), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n572), .B2(KEYINPUT119), .ZN(new_n1127));
  XNOR2_X1  g702(.A(G299), .B(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1121), .A2(KEYINPUT121), .A3(new_n1124), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(KEYINPUT122), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1026), .ZN(new_n1134));
  INV_X1    g709(.A(G1348), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n993), .A2(new_n1134), .B1(new_n1081), .B2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n604), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT122), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1129), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1052), .A2(G1348), .B1(G2067), .B2(new_n1026), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n1026), .A2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G1996), .Z(new_n1146));
  NAND4_X1  g721(.A1(new_n1033), .A2(new_n1034), .A3(new_n980), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n841), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  OAI22_X1  g723(.A1(new_n1142), .A2(new_n1143), .B1(new_n1148), .B2(KEYINPUT59), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(KEYINPUT59), .B2(new_n1148), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1129), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1142), .A2(new_n613), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT60), .B1(new_n1154), .B2(new_n1137), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1126), .A2(new_n1151), .A3(new_n1128), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1150), .A2(new_n1153), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1119), .B1(new_n1141), .B2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1075), .A2(new_n1109), .A3(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(G290), .B(G1986), .Z(new_n1160));
  OR2_X1    g735(.A1(new_n1160), .A2(new_n981), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n998), .A2(new_n997), .A3(new_n985), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1015), .B1(new_n1159), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g738(.A1(G229), .A2(new_n459), .A3(G227), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n895), .A2(new_n656), .A3(new_n1165), .ZN(new_n1166));
  NOR2_X1   g740(.A1(new_n971), .A2(new_n1166), .ZN(G308));
  OR2_X1    g741(.A1(new_n971), .A2(new_n1166), .ZN(G225));
endmodule


