

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  NAND2_X1 U323 ( .A1(n471), .A2(n470), .ZN(n489) );
  XNOR2_X1 U324 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U325 ( .A(n475), .B(n474), .ZN(n505) );
  XOR2_X1 U326 ( .A(n467), .B(KEYINPUT28), .Z(n537) );
  NAND2_X1 U327 ( .A1(n571), .A2(n570), .ZN(n291) );
  AND2_X1 U328 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U329 ( .A(n350), .B(n292), .ZN(n330) );
  XNOR2_X1 U330 ( .A(n427), .B(KEYINPUT119), .ZN(n428) );
  XNOR2_X1 U331 ( .A(n422), .B(n345), .ZN(n346) );
  INV_X1 U332 ( .A(KEYINPUT75), .ZN(n390) );
  XNOR2_X1 U333 ( .A(n430), .B(n330), .ZN(n331) );
  XNOR2_X1 U334 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U335 ( .A(n391), .B(n390), .ZN(n392) );
  INV_X1 U336 ( .A(KEYINPUT24), .ZN(n335) );
  XNOR2_X1 U337 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U338 ( .A(n393), .B(n392), .ZN(n397) );
  NOR2_X1 U339 ( .A1(n472), .A2(n589), .ZN(n473) );
  XNOR2_X1 U340 ( .A(n356), .B(n355), .ZN(n361) );
  XNOR2_X1 U341 ( .A(n338), .B(n337), .ZN(n342) );
  XNOR2_X1 U342 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n482) );
  XOR2_X1 U343 ( .A(KEYINPUT41), .B(n580), .Z(n570) );
  INV_X1 U344 ( .A(G43GAT), .ZN(n476) );
  XNOR2_X1 U345 ( .A(n483), .B(n482), .ZN(n485) );
  XNOR2_X1 U346 ( .A(n476), .B(KEYINPUT40), .ZN(n477) );
  XNOR2_X1 U347 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XNOR2_X1 U348 ( .A(n478), .B(n477), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n294) );
  XNOR2_X1 U350 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n301) );
  XOR2_X1 U352 ( .A(G155GAT), .B(G78GAT), .Z(n296) );
  XNOR2_X1 U353 ( .A(G183GAT), .B(G71GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(n297), .B(G211GAT), .Z(n299) );
  XOR2_X1 U356 ( .A(G15GAT), .B(G127GAT), .Z(n322) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(n322), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U359 ( .A(n301), .B(n300), .ZN(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n303) );
  NAND2_X1 U361 ( .A1(G231GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U363 ( .A(n304), .B(KEYINPUT12), .Z(n308) );
  XNOR2_X1 U364 ( .A(G8GAT), .B(G1GAT), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n305), .B(KEYINPUT70), .ZN(n363) );
  XNOR2_X1 U366 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n306), .B(KEYINPUT72), .ZN(n381) );
  XNOR2_X1 U368 ( .A(n363), .B(n381), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(n310), .B(n309), .Z(n585) );
  XOR2_X1 U371 ( .A(KEYINPUT20), .B(G176GAT), .Z(n312) );
  NAND2_X1 U372 ( .A1(G227GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U374 ( .A(n313), .B(KEYINPUT86), .Z(n321) );
  XOR2_X1 U375 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n315) );
  XNOR2_X1 U376 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U378 ( .A(G169GAT), .B(n316), .ZN(n425) );
  XOR2_X1 U379 ( .A(G190GAT), .B(G134GAT), .Z(n318) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G99GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U382 ( .A(n425), .B(n319), .Z(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n323) );
  XOR2_X1 U384 ( .A(n323), .B(n322), .Z(n327) );
  XOR2_X1 U385 ( .A(KEYINPUT0), .B(KEYINPUT84), .Z(n325) );
  XNOR2_X1 U386 ( .A(G113GAT), .B(KEYINPUT85), .ZN(n324) );
  XNOR2_X1 U387 ( .A(n325), .B(n324), .ZN(n431) );
  XOR2_X1 U388 ( .A(G120GAT), .B(G71GAT), .Z(n382) );
  XNOR2_X1 U389 ( .A(n431), .B(n382), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n569) );
  XOR2_X1 U391 ( .A(G155GAT), .B(KEYINPUT2), .Z(n329) );
  XNOR2_X1 U392 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n430) );
  XOR2_X1 U394 ( .A(G50GAT), .B(G162GAT), .Z(n350) );
  XOR2_X1 U395 ( .A(n331), .B(KEYINPUT22), .Z(n334) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(G78GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n332), .B(G148GAT), .ZN(n399) );
  XNOR2_X1 U398 ( .A(n399), .B(KEYINPUT87), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G22GAT), .Z(n362) );
  XNOR2_X1 U401 ( .A(n362), .B(KEYINPUT23), .ZN(n336) );
  XOR2_X1 U402 ( .A(G211GAT), .B(G218GAT), .Z(n340) );
  XNOR2_X1 U403 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U405 ( .A(G197GAT), .B(n341), .Z(n418) );
  XOR2_X1 U406 ( .A(n342), .B(n418), .Z(n467) );
  XOR2_X1 U407 ( .A(G134GAT), .B(KEYINPUT77), .Z(n443) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n344) );
  XNOR2_X1 U409 ( .A(G92GAT), .B(KEYINPUT64), .ZN(n343) );
  XOR2_X1 U410 ( .A(n344), .B(n343), .Z(n347) );
  XOR2_X1 U411 ( .A(G36GAT), .B(G190GAT), .Z(n422) );
  XNOR2_X1 U412 ( .A(G218GAT), .B(G106GAT), .ZN(n345) );
  XOR2_X1 U413 ( .A(n443), .B(n348), .Z(n356) );
  XNOR2_X1 U414 ( .A(G99GAT), .B(G85GAT), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n349), .B(KEYINPUT74), .ZN(n389) );
  XNOR2_X1 U416 ( .A(n350), .B(n389), .ZN(n354) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n352) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XOR2_X1 U419 ( .A(n352), .B(n351), .Z(n353) );
  XOR2_X1 U420 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n358) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G29GAT), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U423 ( .A(KEYINPUT7), .B(n359), .ZN(n379) );
  XOR2_X1 U424 ( .A(n379), .B(KEYINPUT9), .Z(n360) );
  XOR2_X1 U425 ( .A(n361), .B(n360), .Z(n562) );
  INV_X1 U426 ( .A(n562), .ZN(n407) );
  XOR2_X1 U427 ( .A(n363), .B(n362), .Z(n365) );
  XNOR2_X1 U428 ( .A(G50GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n378) );
  XOR2_X1 U430 ( .A(G197GAT), .B(G15GAT), .Z(n367) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G113GAT), .ZN(n366) );
  XNOR2_X1 U432 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n369) );
  XNOR2_X1 U434 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n368) );
  XNOR2_X1 U435 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U436 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U437 ( .A(KEYINPUT65), .B(KEYINPUT68), .Z(n373) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U440 ( .A(KEYINPUT71), .B(n374), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U442 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U443 ( .A(n380), .B(n379), .Z(n551) );
  INV_X1 U444 ( .A(n551), .ZN(n566) );
  NAND2_X1 U445 ( .A1(n381), .A2(n382), .ZN(n386) );
  INV_X1 U446 ( .A(n381), .ZN(n384) );
  INV_X1 U447 ( .A(n382), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n384), .A2(n383), .ZN(n385) );
  NAND2_X1 U449 ( .A1(n386), .A2(n385), .ZN(n388) );
  AND2_X1 U450 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n389), .B(KEYINPUT73), .ZN(n391) );
  XOR2_X1 U453 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n395) );
  XNOR2_X1 U454 ( .A(G204GAT), .B(KEYINPUT31), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U456 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U457 ( .A(G176GAT), .B(G92GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n398), .B(G64GAT), .ZN(n417) );
  XNOR2_X1 U459 ( .A(n399), .B(n417), .ZN(n400) );
  XOR2_X1 U460 ( .A(n401), .B(n400), .Z(n580) );
  NAND2_X1 U461 ( .A1(n566), .A2(n570), .ZN(n402) );
  XNOR2_X1 U462 ( .A(n402), .B(KEYINPUT46), .ZN(n403) );
  INV_X1 U463 ( .A(n585), .ZN(n559) );
  NAND2_X1 U464 ( .A1(n403), .A2(n559), .ZN(n404) );
  NOR2_X1 U465 ( .A1(n407), .A2(n404), .ZN(n406) );
  XNOR2_X1 U466 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n415) );
  INV_X1 U468 ( .A(KEYINPUT45), .ZN(n409) );
  XOR2_X1 U469 ( .A(KEYINPUT36), .B(n407), .Z(n589) );
  NOR2_X1 U470 ( .A1(n559), .A2(n589), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n410) );
  NOR2_X1 U472 ( .A1(n410), .A2(n580), .ZN(n412) );
  INV_X1 U473 ( .A(KEYINPUT112), .ZN(n411) );
  XNOR2_X1 U474 ( .A(n412), .B(n411), .ZN(n413) );
  NOR2_X1 U475 ( .A1(n413), .A2(n566), .ZN(n414) );
  NOR2_X1 U476 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U477 ( .A(KEYINPUT48), .B(n416), .ZN(n535) );
  XOR2_X1 U478 ( .A(KEYINPUT92), .B(n417), .Z(n420) );
  XNOR2_X1 U479 ( .A(G8GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U481 ( .A(n422), .B(n421), .Z(n424) );
  NAND2_X1 U482 ( .A1(G226GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U484 ( .A(n426), .B(n425), .Z(n528) );
  NOR2_X1 U485 ( .A1(n535), .A2(n528), .ZN(n429) );
  INV_X1 U486 ( .A(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n452) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n451) );
  XOR2_X1 U489 ( .A(G57GAT), .B(G148GAT), .Z(n433) );
  XNOR2_X1 U490 ( .A(G141GAT), .B(G127GAT), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U492 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n435) );
  XNOR2_X1 U493 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n434) );
  XNOR2_X1 U494 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U495 ( .A(n437), .B(n436), .Z(n449) );
  XOR2_X1 U496 ( .A(KEYINPUT5), .B(KEYINPUT89), .Z(n439) );
  XNOR2_X1 U497 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n447) );
  XOR2_X1 U499 ( .A(G85GAT), .B(G162GAT), .Z(n441) );
  XNOR2_X1 U500 ( .A(G29GAT), .B(G120GAT), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U502 ( .A(n443), .B(n442), .Z(n445) );
  NAND2_X1 U503 ( .A1(G225GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n526) );
  NAND2_X1 U508 ( .A1(n452), .A2(n526), .ZN(n479) );
  NOR2_X1 U509 ( .A1(n467), .A2(n479), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n453), .B(KEYINPUT55), .ZN(n572) );
  NOR2_X1 U511 ( .A1(n569), .A2(n572), .ZN(n577) );
  NAND2_X1 U512 ( .A1(n585), .A2(n577), .ZN(n455) );
  XNOR2_X1 U513 ( .A(G183GAT), .B(KEYINPUT122), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n459) );
  NOR2_X1 U515 ( .A1(n569), .A2(n528), .ZN(n456) );
  NOR2_X1 U516 ( .A1(n467), .A2(n456), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n457), .B(KEYINPUT95), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n459), .B(n458), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n467), .A2(n569), .ZN(n460) );
  XOR2_X1 U520 ( .A(n460), .B(KEYINPUT26), .Z(n549) );
  INV_X1 U521 ( .A(n549), .ZN(n480) );
  XNOR2_X1 U522 ( .A(n528), .B(KEYINPUT27), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n480), .A2(n465), .ZN(n461) );
  XOR2_X1 U524 ( .A(KEYINPUT94), .B(n461), .Z(n462) );
  NAND2_X1 U525 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n526), .ZN(n471) );
  NOR2_X1 U527 ( .A1(n465), .A2(n526), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT93), .ZN(n536) );
  INV_X1 U529 ( .A(n537), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n536), .A2(n468), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n569), .A2(n469), .ZN(n470) );
  NAND2_X1 U532 ( .A1(n559), .A2(n489), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT37), .ZN(n523) );
  OR2_X1 U534 ( .A1(n580), .A2(n551), .ZN(n492) );
  NOR2_X1 U535 ( .A1(n523), .A2(n492), .ZN(n475) );
  XNOR2_X1 U536 ( .A(KEYINPUT99), .B(KEYINPUT38), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n569), .A2(n505), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n481), .B(KEYINPUT123), .ZN(n588) );
  OR2_X1 U540 ( .A1(n588), .A2(n551), .ZN(n483) );
  XOR2_X1 U541 ( .A(G197GAT), .B(KEYINPUT124), .Z(n484) );
  XNOR2_X1 U542 ( .A(n485), .B(n484), .ZN(G1352GAT) );
  NAND2_X1 U543 ( .A1(n562), .A2(n585), .ZN(n488) );
  XNOR2_X1 U544 ( .A(KEYINPUT16), .B(KEYINPUT83), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT82), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n490) );
  NAND2_X1 U547 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U548 ( .A(KEYINPUT97), .B(n491), .Z(n510) );
  OR2_X1 U549 ( .A1(n492), .A2(n510), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n526), .A2(n499), .ZN(n493) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(n493), .Z(n494) );
  XNOR2_X1 U552 ( .A(G1GAT), .B(n494), .ZN(G1324GAT) );
  NOR2_X1 U553 ( .A1(n528), .A2(n499), .ZN(n495) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n569), .A2(n499), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(n498), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n537), .A2(n499), .ZN(n500) );
  XOR2_X1 U560 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U561 ( .A1(n505), .A2(n526), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT100), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT39), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n505), .A2(n528), .ZN(n504) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n504), .Z(G1329GAT) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n507) );
  NOR2_X1 U568 ( .A1(n537), .A2(n505), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1331GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT103), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT102), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n551), .A2(n570), .ZN(n524) );
  OR2_X1 U574 ( .A1(n524), .A2(n510), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n526), .A2(n518), .ZN(n511) );
  XOR2_X1 U576 ( .A(n512), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n528), .A2(n518), .ZN(n514) );
  XNOR2_X1 U578 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n569), .A2(n518), .ZN(n516) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(n516), .Z(n517) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n517), .ZN(G1334GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n537), .ZN(n522) );
  XOR2_X1 U585 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n520) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT108), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1335GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n525), .B(KEYINPUT109), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n526), .A2(n531), .ZN(n527) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n527), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n531), .ZN(n529) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n569), .A2(n531), .ZN(n530) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n537), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U600 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  XOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT113), .Z(n540) );
  NOR2_X1 U602 ( .A1(n535), .A2(n536), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n537), .A2(n550), .ZN(n538) );
  NOR2_X1 U604 ( .A1(n569), .A2(n538), .ZN(n545) );
  NAND2_X1 U605 ( .A1(n545), .A2(n566), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U608 ( .A1(n545), .A2(n570), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n585), .A2(n545), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(KEYINPUT50), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U614 ( .A1(n545), .A2(n407), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n551), .A2(n561), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n558) );
  INV_X1 U624 ( .A(n570), .ZN(n556) );
  NOR2_X1 U625 ( .A1(n556), .A2(n561), .ZN(n557) );
  XOR2_X1 U626 ( .A(n558), .B(n557), .Z(G1345GAT) );
  NOR2_X1 U627 ( .A1(n559), .A2(n561), .ZN(n560) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n577), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n574) );
  INV_X1 U637 ( .A(n569), .ZN(n571) );
  OR2_X1 U638 ( .A1(n291), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(G176GAT), .B(KEYINPUT56), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n407), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT58), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(n579), .ZN(G1351GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n582) );
  INV_X1 U646 ( .A(n588), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n580), .A2(n584), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT126), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G211GAT), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

