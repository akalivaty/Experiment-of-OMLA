

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(n411), .B(KEYINPUT115), .ZN(n412) );
  XNOR2_X1 U323 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U324 ( .A(n413), .B(n412), .ZN(n536) );
  XNOR2_X1 U325 ( .A(n308), .B(n307), .ZN(n405) );
  NOR2_X1 U326 ( .A1(n539), .A2(n452), .ZN(n568) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U328 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  XNOR2_X1 U329 ( .A(G176GAT), .B(G204GAT), .ZN(n290) );
  XNOR2_X1 U330 ( .A(n290), .B(G64GAT), .ZN(n418) );
  INV_X1 U331 ( .A(n418), .ZN(n292) );
  XOR2_X1 U332 ( .A(G92GAT), .B(G85GAT), .Z(n386) );
  INV_X1 U333 ( .A(n386), .ZN(n291) );
  NAND2_X1 U334 ( .A1(n292), .A2(n291), .ZN(n294) );
  NAND2_X1 U335 ( .A1(n418), .A2(n386), .ZN(n293) );
  NAND2_X1 U336 ( .A1(n294), .A2(n293), .ZN(n296) );
  AND2_X1 U337 ( .A1(G230GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n297), .B(KEYINPUT32), .ZN(n298) );
  INV_X1 U340 ( .A(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(KEYINPUT13), .B(G57GAT), .Z(n367) );
  XNOR2_X1 U342 ( .A(n367), .B(KEYINPUT33), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n308) );
  XNOR2_X1 U344 ( .A(G99GAT), .B(G71GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n301), .B(G120GAT), .ZN(n311) );
  XNOR2_X1 U346 ( .A(G106GAT), .B(G78GAT), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n302), .B(G148GAT), .ZN(n326) );
  XOR2_X1 U348 ( .A(n311), .B(n326), .Z(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n304) );
  XNOR2_X1 U350 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT41), .B(n405), .Z(n556) );
  XOR2_X1 U353 ( .A(n556), .B(KEYINPUT107), .Z(n541) );
  XOR2_X1 U354 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n314) );
  XOR2_X1 U355 ( .A(KEYINPUT20), .B(KEYINPUT79), .Z(n310) );
  XNOR2_X1 U356 ( .A(KEYINPUT83), .B(G176GAT), .ZN(n309) );
  XNOR2_X1 U357 ( .A(n310), .B(n309), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U360 ( .A(KEYINPUT0), .B(G127GAT), .Z(n443) );
  XOR2_X1 U361 ( .A(G43GAT), .B(G134GAT), .Z(n396) );
  XOR2_X1 U362 ( .A(n443), .B(n396), .Z(n316) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U365 ( .A(n318), .B(n317), .Z(n325) );
  XOR2_X1 U366 ( .A(G113GAT), .B(G15GAT), .Z(n347) );
  XOR2_X1 U367 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n320) );
  XNOR2_X1 U368 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U370 ( .A(n321), .B(KEYINPUT82), .Z(n323) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G183GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n426) );
  XNOR2_X1 U373 ( .A(n347), .B(n426), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n539) );
  XOR2_X1 U375 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n328) );
  XNOR2_X1 U376 ( .A(n326), .B(KEYINPUT85), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(n329), .ZN(n344) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n330), .B(G162GAT), .ZN(n384) );
  XOR2_X1 U381 ( .A(n384), .B(KEYINPUT86), .Z(n332) );
  NAND2_X1 U382 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n334) );
  XNOR2_X1 U385 ( .A(G204GAT), .B(KEYINPUT87), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U387 ( .A(n336), .B(n335), .Z(n342) );
  XOR2_X1 U388 ( .A(G155GAT), .B(KEYINPUT2), .Z(n338) );
  XNOR2_X1 U389 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n442) );
  XOR2_X1 U391 ( .A(G211GAT), .B(KEYINPUT21), .Z(n340) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n417) );
  XNOR2_X1 U394 ( .A(n442), .B(n417), .ZN(n341) );
  XNOR2_X1 U395 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n472) );
  XOR2_X1 U397 ( .A(G1GAT), .B(G8GAT), .Z(n346) );
  XNOR2_X1 U398 ( .A(G22GAT), .B(KEYINPUT68), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n368) );
  XOR2_X1 U400 ( .A(n368), .B(n347), .Z(n349) );
  XNOR2_X1 U401 ( .A(G50GAT), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n354) );
  XNOR2_X1 U403 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n350), .B(KEYINPUT8), .ZN(n385) );
  XOR2_X1 U405 ( .A(n385), .B(KEYINPUT66), .Z(n352) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U408 ( .A(n354), .B(n353), .Z(n362) );
  XOR2_X1 U409 ( .A(G197GAT), .B(G141GAT), .Z(n356) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(G36GAT), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n358) );
  XNOR2_X1 U413 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n573) );
  NAND2_X1 U417 ( .A1(n573), .A2(n556), .ZN(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n382) );
  XOR2_X1 U420 ( .A(G78GAT), .B(G127GAT), .Z(n366) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(G71GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n381) );
  XOR2_X1 U423 ( .A(n367), .B(G211GAT), .Z(n370) );
  XNOR2_X1 U424 ( .A(n368), .B(G155GAT), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U426 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n372) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n374), .B(n373), .Z(n379) );
  XOR2_X1 U430 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n376) );
  XNOR2_X1 U431 ( .A(G15GAT), .B(G64GAT), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n377), .B(KEYINPUT76), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U435 ( .A(n381), .B(n380), .Z(n581) );
  NOR2_X1 U436 ( .A1(n382), .A2(n581), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n383), .B(KEYINPUT113), .ZN(n401) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n400) );
  XOR2_X1 U439 ( .A(G36GAT), .B(KEYINPUT74), .Z(n422) );
  XOR2_X1 U440 ( .A(n422), .B(n386), .Z(n388) );
  NAND2_X1 U441 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT10), .B(G106GAT), .Z(n390) );
  XNOR2_X1 U444 ( .A(G190GAT), .B(G99GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n398) );
  XOR2_X1 U447 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n394) );
  XNOR2_X1 U448 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U452 ( .A(n400), .B(n399), .ZN(n567) );
  NOR2_X1 U453 ( .A1(n401), .A2(n567), .ZN(n402) );
  XNOR2_X1 U454 ( .A(n402), .B(KEYINPUT47), .ZN(n410) );
  INV_X1 U455 ( .A(n581), .ZN(n499) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n403) );
  INV_X1 U457 ( .A(n567), .ZN(n480) );
  XNOR2_X1 U458 ( .A(n403), .B(n480), .ZN(n497) );
  NOR2_X1 U459 ( .A1(n499), .A2(n497), .ZN(n404) );
  XNOR2_X1 U460 ( .A(KEYINPUT45), .B(n404), .ZN(n407) );
  BUF_X1 U461 ( .A(n405), .Z(n577) );
  NOR2_X1 U462 ( .A1(n573), .A2(n577), .ZN(n406) );
  NAND2_X1 U463 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT114), .B(n408), .ZN(n409) );
  NAND2_X1 U465 ( .A1(n410), .A2(n409), .ZN(n413) );
  XOR2_X1 U466 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n411) );
  XOR2_X1 U467 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n415) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U470 ( .A(n416), .B(KEYINPUT93), .Z(n420) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U473 ( .A(n421), .B(G92GAT), .Z(n424) );
  XNOR2_X1 U474 ( .A(G8GAT), .B(n422), .ZN(n423) );
  XNOR2_X1 U475 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U476 ( .A(n426), .B(n425), .Z(n470) );
  NAND2_X1 U477 ( .A1(n536), .A2(n470), .ZN(n427) );
  XNOR2_X1 U478 ( .A(n427), .B(KEYINPUT121), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n428), .B(KEYINPUT54), .ZN(n450) );
  XOR2_X1 U480 ( .A(G85GAT), .B(G148GAT), .Z(n430) );
  XNOR2_X1 U481 ( .A(G120GAT), .B(G134GAT), .ZN(n429) );
  XNOR2_X1 U482 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT92), .B(G57GAT), .Z(n432) );
  XNOR2_X1 U484 ( .A(G113GAT), .B(G1GAT), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U486 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT90), .Z(n436) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(KEYINPUT6), .B(n437), .ZN(n438) );
  XNOR2_X1 U491 ( .A(n439), .B(n438), .ZN(n449) );
  XOR2_X1 U492 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n441) );
  XNOR2_X1 U493 ( .A(KEYINPUT5), .B(KEYINPUT91), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U495 ( .A(G162GAT), .B(n442), .Z(n445) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U498 ( .A(n447), .B(n446), .Z(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(n553) );
  NAND2_X1 U500 ( .A1(n450), .A2(n553), .ZN(n458) );
  NOR2_X1 U501 ( .A1(n472), .A2(n458), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U503 ( .A1(n541), .A2(n568), .ZN(n456) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .Z(n454) );
  XNOR2_X1 U505 ( .A(KEYINPUT57), .B(KEYINPUT122), .ZN(n453) );
  INV_X1 U506 ( .A(G218GAT), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n472), .A2(n539), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n457), .B(KEYINPUT26), .ZN(n469) );
  NOR2_X1 U509 ( .A1(n458), .A2(n469), .ZN(n582) );
  INV_X1 U510 ( .A(n582), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n497), .A2(n459), .ZN(n460) );
  XNOR2_X1 U512 ( .A(KEYINPUT62), .B(n460), .ZN(n461) );
  XNOR2_X1 U513 ( .A(n462), .B(n461), .ZN(G1355GAT) );
  INV_X1 U514 ( .A(n573), .ZN(n513) );
  NOR2_X1 U515 ( .A1(n577), .A2(n513), .ZN(n503) );
  XOR2_X1 U516 ( .A(n472), .B(KEYINPUT28), .Z(n532) );
  XOR2_X1 U517 ( .A(n470), .B(KEYINPUT27), .Z(n468) );
  INV_X1 U518 ( .A(n468), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n532), .A2(n463), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n553), .A2(n464), .ZN(n537) );
  XNOR2_X1 U521 ( .A(n537), .B(KEYINPUT96), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n539), .B(KEYINPUT84), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(n467), .B(KEYINPUT97), .ZN(n479) );
  INV_X1 U525 ( .A(n553), .ZN(n477) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n551) );
  INV_X1 U527 ( .A(n470), .ZN(n528) );
  NOR2_X1 U528 ( .A1(n539), .A2(n528), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(n473), .B(KEYINPUT25), .Z(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT98), .B(n474), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n551), .A2(n475), .ZN(n476) );
  NOR2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n498) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n482) );
  NAND2_X1 U536 ( .A1(n581), .A2(n480), .ZN(n481) );
  XNOR2_X1 U537 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U538 ( .A(n483), .B(KEYINPUT77), .ZN(n484) );
  NOR2_X1 U539 ( .A1(n498), .A2(n484), .ZN(n485) );
  XOR2_X1 U540 ( .A(KEYINPUT99), .B(n485), .Z(n515) );
  NAND2_X1 U541 ( .A1(n503), .A2(n515), .ZN(n495) );
  NOR2_X1 U542 ( .A1(n553), .A2(n495), .ZN(n487) );
  XNOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U545 ( .A(G1GAT), .B(n488), .Z(G1324GAT) );
  NOR2_X1 U546 ( .A1(n528), .A2(n495), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n495), .A2(n539), .ZN(n494) );
  XOR2_X1 U550 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n492) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U554 ( .A1(n532), .A2(n495), .ZN(n496) );
  XOR2_X1 U555 ( .A(G22GAT), .B(n496), .Z(G1327GAT) );
  NOR2_X1 U556 ( .A1(n498), .A2(n497), .ZN(n500) );
  NAND2_X1 U557 ( .A1(n500), .A2(n499), .ZN(n502) );
  XOR2_X1 U558 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n501) );
  XNOR2_X1 U559 ( .A(n502), .B(n501), .ZN(n525) );
  NAND2_X1 U560 ( .A1(n503), .A2(n525), .ZN(n504) );
  XNOR2_X1 U561 ( .A(n504), .B(KEYINPUT38), .ZN(n511) );
  NOR2_X1 U562 ( .A1(n511), .A2(n553), .ZN(n505) );
  XNOR2_X1 U563 ( .A(n505), .B(KEYINPUT39), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n506), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n511), .A2(n528), .ZN(n507) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(n507), .Z(n508) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n508), .ZN(G1329GAT) );
  NOR2_X1 U568 ( .A1(n539), .A2(n511), .ZN(n509) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(n509), .Z(n510) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NOR2_X1 U571 ( .A1(n532), .A2(n511), .ZN(n512) );
  XOR2_X1 U572 ( .A(G50GAT), .B(n512), .Z(G1331GAT) );
  NAND2_X1 U573 ( .A1(n513), .A2(n541), .ZN(n514) );
  XOR2_X1 U574 ( .A(KEYINPUT108), .B(n514), .Z(n524) );
  NAND2_X1 U575 ( .A1(n515), .A2(n524), .ZN(n521) );
  NOR2_X1 U576 ( .A1(n553), .A2(n521), .ZN(n516) );
  XOR2_X1 U577 ( .A(n516), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U578 ( .A(G57GAT), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n528), .A2(n521), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U582 ( .A1(n539), .A2(n521), .ZN(n520) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n520), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n532), .A2(n521), .ZN(n523) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X1 U588 ( .A1(n553), .A2(n531), .ZN(n526) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n526), .Z(n527) );
  XNOR2_X1 U590 ( .A(KEYINPUT110), .B(n527), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n528), .A2(n531), .ZN(n529) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n529), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n539), .A2(n531), .ZN(n530) );
  XOR2_X1 U594 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n547), .A2(n573), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U604 ( .A1(n547), .A2(n541), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n547), .A2(n581), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n545), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n549) );
  NAND2_X1 U611 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U612 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n536), .ZN(n552) );
  NOR2_X1 U615 ( .A1(n553), .A2(n552), .ZN(n563) );
  NAND2_X1 U616 ( .A1(n563), .A2(n573), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n554), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n558) );
  NAND2_X1 U620 ( .A1(n563), .A2(n556), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT119), .Z(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n563), .A2(n581), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT120), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n562), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n567), .ZN(n564) );
  XNOR2_X1 U628 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n568), .A2(n573), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n568), .A2(n581), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  NAND2_X1 U639 ( .A1(n582), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n582), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n580), .B(G204GAT), .Z(G1353GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n584) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(n585), .ZN(G1354GAT) );
endmodule

