//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n205), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT25), .ZN(new_n220));
  AND3_X1   g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n223), .A2(new_n224), .A3(new_n210), .A4(new_n205), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n212), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n229), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n204), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(new_n230), .A3(new_n208), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT25), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT26), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(new_n206), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT28), .B1(new_n242), .B2(new_n204), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT27), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G183gat), .ZN(new_n246));
  AND4_X1   g045(.A1(KEYINPUT28), .A2(new_n244), .A3(new_n246), .A4(new_n204), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n241), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n234), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n226), .A2(new_n234), .A3(new_n248), .A4(KEYINPUT70), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G211gat), .A2(G218gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259));
  AND2_X1   g058(.A1(G197gat), .A2(G204gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n264));
  XNOR2_X1  g063(.A(G211gat), .B(G218gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n266), .A3(new_n258), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n258), .B2(new_n266), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n249), .A2(new_n276), .A3(new_n252), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n255), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT71), .ZN(new_n280));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n251), .A2(new_n254), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n253), .B1(new_n283), .B2(new_n276), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n242), .A2(new_n204), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n204), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n289), .A2(new_n241), .B1(new_n233), .B2(KEYINPUT25), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n252), .B1(new_n290), .B2(new_n226), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(new_n271), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n278), .B(new_n282), .C1(new_n284), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n291), .A2(new_n271), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT29), .B1(new_n251), .B2(new_n254), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(new_n253), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT72), .A3(new_n278), .A4(new_n282), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n282), .B1(new_n299), .B2(new_n278), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n299), .A2(new_n278), .A3(new_n282), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT30), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(G155gat), .B2(G162gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G155gat), .B(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G120gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G113gat), .ZN(new_n325));
  INV_X1    g124(.A(G113gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G120gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G127gat), .B(G134gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n328), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G127gat), .B(G134gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(KEYINPUT1), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n312), .A3(new_n322), .A4(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G225gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  OR3_X1    g140(.A1(new_n339), .A2(KEYINPUT81), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT81), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(KEYINPUT39), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n336), .A2(KEYINPUT67), .A3(new_n337), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT67), .B1(new_n336), .B2(new_n337), .ZN(new_n347));
  AND3_X1   g146(.A1(new_n312), .A2(new_n322), .A3(KEYINPUT75), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT75), .B1(new_n312), .B2(new_n322), .ZN(new_n349));
  OAI22_X1  g148(.A1(new_n346), .A2(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n350), .B2(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT77), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT73), .B(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n312), .A2(new_n322), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n312), .A2(new_n322), .A3(KEYINPUT74), .A4(new_n353), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n323), .A2(KEYINPUT3), .B1(new_n337), .B2(new_n336), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n323), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n312), .A2(new_n322), .A3(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n331), .B2(new_n332), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n336), .A2(KEYINPUT67), .A3(new_n337), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n345), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n360), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n344), .B1(new_n373), .B2(new_n341), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G1gat), .B(G29gat), .Z(new_n376));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT39), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n381), .A3(new_n341), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n375), .A2(KEYINPUT40), .A3(new_n380), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n380), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n360), .A2(new_n385), .A3(new_n340), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n352), .A3(new_n372), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n368), .A3(KEYINPUT4), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n338), .A2(new_n369), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n389), .A2(new_n360), .A3(new_n340), .A4(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n339), .B2(new_n341), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n380), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT40), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n384), .A2(new_n374), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n305), .A2(new_n383), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n380), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n370), .A2(new_n371), .A3(new_n345), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n371), .B1(new_n370), .B2(new_n345), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n386), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n391), .A2(new_n392), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n380), .A3(new_n393), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT6), .B(new_n400), .C1(new_n403), .C2(new_n404), .ZN(new_n409));
  AND2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n295), .A2(new_n300), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT84), .B(KEYINPUT37), .Z(new_n412));
  NAND3_X1  g211(.A1(new_n299), .A2(new_n278), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n282), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n299), .B2(new_n278), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT38), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n283), .A2(new_n276), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n291), .B1(new_n419), .B2(new_n252), .ZN(new_n420));
  AND2_X1   g219(.A1(new_n268), .A2(new_n270), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n275), .B1(new_n255), .B2(new_n277), .ZN(new_n422));
  OAI22_X1  g221(.A1(new_n420), .A2(new_n421), .B1(KEYINPUT83), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n422), .A2(KEYINPUT83), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT37), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n415), .A2(KEYINPUT38), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n418), .A4(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n305), .A2(new_n396), .A3(KEYINPUT82), .A4(new_n383), .ZN(new_n429));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n353), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n261), .A2(new_n262), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n276), .B1(new_n432), .B2(new_n269), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(new_n433), .B2(KEYINPUT78), .ZN(new_n434));
  AOI211_X1 g233(.A(KEYINPUT78), .B(KEYINPUT29), .C1(new_n263), .C2(new_n267), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n364), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n421), .B1(new_n358), .B2(new_n276), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n268), .A2(new_n270), .A3(new_n276), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT3), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n323), .ZN(new_n443));
  INV_X1    g242(.A(new_n430), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n268), .A2(new_n273), .A3(new_n270), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n273), .B1(new_n268), .B2(new_n270), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n356), .B2(new_n357), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n443), .B(new_n444), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n439), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G22gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT31), .B(G50gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT79), .B(G22gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n449), .A3(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n451), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n457), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT29), .B1(new_n263), .B2(new_n267), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n353), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(new_n435), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n464), .A2(new_n364), .B1(new_n421), .B2(new_n448), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n358), .A2(new_n276), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n430), .B1(new_n275), .B2(new_n466), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n430), .A2(new_n465), .B1(new_n467), .B2(new_n443), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT80), .B1(new_n468), .B2(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470));
  INV_X1    g269(.A(new_n456), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n460), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n459), .B1(new_n473), .B2(new_n455), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n399), .A2(new_n428), .A3(new_n429), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n450), .B2(new_n471), .ZN(new_n476));
  AOI211_X1 g275(.A(KEYINPUT80), .B(new_n456), .C1(new_n439), .C2(new_n449), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n457), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n458), .B1(new_n478), .B2(new_n454), .ZN(new_n479));
  INV_X1    g278(.A(new_n408), .ZN(new_n480));
  INV_X1    g279(.A(new_n409), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n301), .B(new_n304), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n290), .A2(new_n367), .A3(new_n366), .A4(new_n226), .ZN(new_n483));
  INV_X1    g282(.A(G227gat), .ZN(new_n484));
  INV_X1    g283(.A(G233gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n249), .A2(new_n368), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT32), .ZN(new_n489));
  XOR2_X1   g288(.A(G15gat), .B(G43gat), .Z(new_n490));
  XNOR2_X1  g289(.A(G71gat), .B(G99gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n483), .A2(new_n487), .ZN(new_n497));
  INV_X1    g296(.A(new_n486), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g298(.A(KEYINPUT34), .B(new_n486), .C1(new_n483), .C2(new_n487), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n495), .A2(new_n499), .A3(new_n500), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n489), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT34), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n496), .A3(new_n498), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n488), .A2(new_n494), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n493), .ZN(new_n509));
  INV_X1    g308(.A(new_n489), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n501), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n504), .A2(KEYINPUT36), .A3(new_n511), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n479), .A2(new_n482), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n475), .A2(new_n516), .ZN(new_n517));
  NOR3_X1   g316(.A1(new_n502), .A2(new_n503), .A3(new_n489), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n510), .B1(new_n509), .B2(new_n501), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n474), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT35), .B1(new_n521), .B2(new_n482), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n410), .A2(new_n305), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n479), .A2(new_n512), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  INV_X1    g332(.A(G15gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(G22gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n536), .A2(G15gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G8gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT87), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n539), .A2(new_n542), .A3(G8gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT88), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n532), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(G8gat), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n530), .B(KEYINPUT88), .C1(new_n531), .C2(G1gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n538), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NOR3_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(G29gat), .ZN(new_n553));
  INV_X1    g352(.A(G36gat), .ZN(new_n554));
  OAI22_X1  g353(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G43gat), .B(G50gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(KEYINPUT15), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n556), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  XOR2_X1   g357(.A(G43gat), .B(G50gat), .Z(new_n559));
  INV_X1    g358(.A(KEYINPUT15), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT14), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n553), .A3(new_n554), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n552), .A2(KEYINPUT85), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n551), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n557), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n569), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n569), .B2(new_n572), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n547), .A2(new_n546), .A3(new_n538), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n545), .A2(new_n576), .B1(new_n540), .B2(KEYINPUT87), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT17), .B(new_n557), .C1(new_n562), .C2(new_n568), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n543), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n529), .B(new_n570), .C1(new_n575), .C2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT18), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n549), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n583), .B(new_n578), .C1(new_n573), .C2(new_n574), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n570), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT89), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(new_n549), .B2(new_n569), .ZN(new_n587));
  INV_X1    g386(.A(new_n569), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n577), .A2(new_n588), .A3(KEYINPUT89), .A4(new_n543), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n570), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n529), .B(KEYINPUT13), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n585), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G113gat), .B(G141gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G197gat), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT11), .B(G169gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT12), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT90), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n582), .A2(new_n598), .A3(new_n585), .A4(new_n592), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n593), .A2(KEYINPUT90), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(KEYINPUT95), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT93), .B(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(G85gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n611), .A2(new_n612), .B1(KEYINPUT8), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(G99gat), .ZN(new_n615));
  INV_X1    g414(.A(G106gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT7), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n614), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n618), .B1(new_n614), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n610), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n611), .A2(new_n612), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n613), .A2(KEYINPUT8), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n620), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n626), .A2(new_n613), .A3(new_n617), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n614), .A2(new_n618), .A3(new_n620), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(KEYINPUT95), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G71gat), .B(G78gat), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT9), .ZN(new_n632));
  INV_X1    g431(.A(G71gat), .ZN(new_n633));
  INV_X1    g432(.A(G78gat), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G57gat), .B(G64gat), .Z(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n630), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n642), .B(new_n610), .C1(new_n621), .C2(new_n622), .ZN(new_n643));
  INV_X1    g442(.A(G230gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n485), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n609), .B1(new_n646), .B2(KEYINPUT96), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(KEYINPUT96), .B2(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT10), .B1(new_n641), .B2(new_n643), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT94), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n621), .B2(new_n622), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n628), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n654), .A2(new_n655), .A3(new_n640), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n649), .B1(new_n650), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n609), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n643), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n655), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT10), .A3(new_n642), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n645), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n646), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n659), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT21), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n583), .B1(new_n669), .B2(new_n640), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n640), .A2(new_n669), .ZN(new_n671));
  XNOR2_X1  g470(.A(G127gat), .B(G155gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n670), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G231gat), .A2(G233gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT91), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G183gat), .B(G211gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n674), .B(new_n680), .ZN(new_n681));
  AND2_X1   g480(.A1(G232gat), .A2(G233gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT41), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT92), .ZN(new_n684));
  XNOR2_X1  g483(.A(G134gat), .B(G162gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n662), .A2(new_n569), .B1(KEYINPUT41), .B2(new_n682), .ZN(new_n688));
  XOR2_X1   g487(.A(G190gat), .B(G218gat), .Z(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n578), .B(new_n654), .C1(new_n573), .C2(new_n574), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n690), .B1(new_n688), .B2(new_n691), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n686), .A3(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n528), .A2(new_n606), .A3(new_n668), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n410), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g501(.A1(new_n700), .A2(new_n305), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n546), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT97), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT16), .B(G8gat), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(G1325gat));
  NAND3_X1  g508(.A1(new_n700), .A2(new_n534), .A3(new_n520), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n514), .A2(new_n515), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(new_n534), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n700), .A2(new_n479), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT98), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(new_n698), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n517), .B2(new_n527), .ZN(new_n720));
  INV_X1    g519(.A(new_n681), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n605), .A2(new_n667), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n410), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n723), .A2(G29gat), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT45), .Z(new_n726));
  NAND3_X1  g525(.A1(new_n528), .A2(KEYINPUT44), .A3(new_n698), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  AOI22_X1  g527(.A1(new_n475), .A2(new_n516), .B1(new_n522), .B2(new_n526), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g530(.A(new_n722), .B(KEYINPUT99), .Z(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n724), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n726), .A2(new_n734), .ZN(G1328gat));
  INV_X1    g534(.A(new_n305), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n723), .A2(G36gat), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT100), .B1(new_n733), .B2(new_n736), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G36gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n733), .A2(KEYINPUT100), .A3(new_n736), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(G1329gat));
  NAND2_X1  g541(.A1(new_n712), .A2(G43gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n723), .A2(new_n512), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n733), .A2(new_n743), .B1(G43gat), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g545(.A1(new_n479), .A2(G50gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n723), .A2(new_n474), .ZN(new_n748));
  OAI22_X1  g547(.A1(new_n733), .A2(new_n747), .B1(G50gat), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n605), .A2(new_n699), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n729), .A2(new_n668), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n410), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT101), .B(G57gat), .Z(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1332gat));
  AOI21_X1  g554(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT102), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1333gat));
  NAND3_X1  g559(.A1(new_n752), .A2(new_n633), .A3(new_n520), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n752), .A2(new_n712), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n633), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g563(.A1(new_n752), .A2(new_n479), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n606), .A2(new_n721), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n667), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT103), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n731), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n724), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT51), .B1(new_n720), .B2(new_n767), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  INV_X1    g572(.A(new_n767), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n729), .A2(new_n773), .A3(new_n719), .A4(new_n774), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n776), .A2(new_n612), .A3(new_n410), .A4(new_n667), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n771), .A2(new_n777), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n727), .A2(new_n730), .A3(new_n769), .A4(new_n305), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n611), .B1(new_n779), .B2(KEYINPUT107), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(KEYINPUT107), .B2(new_n779), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n736), .A2(new_n668), .A3(G92gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n772), .B2(new_n775), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT52), .B1(new_n783), .B2(KEYINPUT106), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n781), .B(new_n784), .C1(KEYINPUT106), .C2(new_n783), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT105), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT104), .ZN(new_n788));
  INV_X1    g587(.A(new_n611), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n783), .A2(new_n788), .B1(new_n789), .B2(new_n779), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT104), .B(new_n782), .C1(new_n772), .C2(new_n775), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n786), .B(new_n787), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n783), .A2(new_n788), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n779), .A2(new_n789), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT105), .B1(new_n795), .B2(KEYINPUT52), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n785), .B1(new_n792), .B2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n770), .B2(new_n711), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n776), .A2(new_n615), .A3(new_n520), .A4(new_n667), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n776), .A2(new_n616), .A3(new_n479), .A4(new_n667), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n770), .A2(new_n474), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n802), .B2(new_n616), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT53), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n801), .B(new_n805), .C1(new_n802), .C2(new_n616), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(G1339gat));
  NAND3_X1  g606(.A1(new_n605), .A2(new_n668), .A3(new_n699), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n609), .B1(new_n664), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n661), .A2(new_n645), .A3(new_n663), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n814), .A2(new_n815), .B1(new_n657), .B2(new_n648), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n590), .A2(new_n591), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n529), .B1(new_n584), .B2(new_n570), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n597), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n602), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT108), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n602), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n816), .A2(new_n817), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n721), .B1(new_n825), .B2(new_n698), .ZN(new_n826));
  INV_X1    g625(.A(new_n821), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n698), .B1(new_n827), .B2(new_n667), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n812), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n659), .B1(new_n657), .B2(KEYINPUT54), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n815), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n658), .A3(new_n817), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n828), .B1(new_n605), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n809), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT109), .B1(new_n834), .B2(new_n479), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n822), .A2(new_n824), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n698), .B1(new_n836), .B2(new_n832), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n837), .A3(new_n681), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n808), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT109), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(new_n474), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n724), .A2(new_n305), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n520), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n605), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n834), .A2(new_n724), .A3(new_n521), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n736), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n606), .A2(new_n326), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT110), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(G1340gat));
  OAI21_X1  g649(.A(G120gat), .B1(new_n844), .B2(new_n668), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n667), .A2(new_n324), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(KEYINPUT111), .Z(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n847), .B2(new_n853), .ZN(G1341gat));
  INV_X1    g653(.A(G127gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n844), .A2(new_n855), .A3(new_n681), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n847), .A2(KEYINPUT112), .A3(new_n681), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(G127gat), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT112), .B1(new_n847), .B2(new_n681), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n736), .A2(new_n698), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT113), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  XOR2_X1   g664(.A(new_n865), .B(KEYINPUT56), .Z(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n844), .B2(new_n719), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT114), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT114), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n866), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n871), .ZN(G1343gat));
  NOR2_X1   g671(.A1(new_n834), .A2(new_n724), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n712), .A2(new_n474), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n606), .A2(new_n313), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT116), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n873), .A2(new_n736), .A3(new_n874), .A4(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT117), .Z(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n474), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT115), .A4(new_n681), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n808), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT115), .B1(new_n826), .B2(new_n833), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n834), .B2(new_n474), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n843), .A2(new_n711), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n606), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(G141gat), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n878), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n886), .A2(KEYINPUT118), .A3(new_n606), .A4(new_n887), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n892), .A2(G141gat), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n873), .A2(new_n874), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n305), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT58), .B1(new_n897), .B2(new_n876), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n894), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n890), .B1(new_n899), .B2(new_n900), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n315), .A3(new_n667), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n315), .C1(new_n903), .C2(new_n667), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n474), .B1(new_n838), .B2(new_n808), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT120), .B(new_n879), .C1(new_n834), .C2(new_n474), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n839), .A2(new_n880), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n667), .A3(new_n887), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n905), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n902), .B1(new_n904), .B2(new_n913), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n319), .A3(new_n721), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n903), .A2(new_n721), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n915), .B1(new_n916), .B2(new_n319), .ZN(G1346gat));
  AND2_X1   g716(.A1(new_n903), .A2(new_n698), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n864), .A2(new_n320), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n918), .A2(new_n320), .B1(new_n896), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n736), .A2(new_n410), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n839), .A2(new_n524), .A3(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n606), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n736), .A2(new_n410), .A3(new_n512), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n842), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n605), .A2(new_n213), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1348gat));
  NAND3_X1  g727(.A1(new_n926), .A2(G176gat), .A3(new_n667), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n930), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n923), .B2(new_n667), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G1349gat));
  NAND2_X1  g733(.A1(new_n926), .A2(new_n721), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G183gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n923), .A2(new_n242), .A3(new_n721), .ZN(new_n937));
  XNOR2_X1  g736(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n204), .A3(new_n698), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n842), .A2(new_n698), .A3(new_n925), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n943), .A2(new_n944), .A3(G190gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n943), .B2(G190gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT123), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n949), .B(new_n942), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1351gat));
  NAND2_X1  g750(.A1(new_n711), .A2(new_n921), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n834), .A2(new_n474), .A3(new_n952), .ZN(new_n953));
  XOR2_X1   g752(.A(KEYINPUT124), .B(G197gat), .Z(new_n954));
  NAND3_X1  g753(.A1(new_n953), .A2(new_n606), .A3(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n952), .B(KEYINPUT125), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n911), .A2(new_n956), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n957), .A2(new_n606), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n958), .B2(new_n954), .ZN(G1352gat));
  INV_X1    g758(.A(G204gat), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n953), .A2(new_n960), .A3(new_n667), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n962), .A2(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n911), .A2(new_n667), .A3(new_n956), .ZN(new_n966));
  OAI221_X1 g765(.A(new_n965), .B1(new_n963), .B2(new_n961), .C1(new_n966), .C2(new_n960), .ZN(G1353gat));
  INV_X1    g766(.A(G211gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n953), .A2(new_n968), .A3(new_n721), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n952), .A2(new_n681), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n911), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  AOI211_X1 g772(.A(new_n973), .B(new_n968), .C1(new_n911), .C2(new_n970), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT127), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(KEYINPUT127), .B(new_n969), .C1(new_n972), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n953), .B2(new_n698), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n698), .A2(G218gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n980), .B1(new_n957), .B2(new_n981), .ZN(G1355gat));
endmodule


