//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT87), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G141gat), .B(G148gat), .Z(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT2), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G141gat), .B(G148gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n212), .C1(new_n217), .C2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT29), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223));
  INV_X1    g022(.A(G211gat), .ZN(new_n224));
  INV_X1    g023(.A(G218gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n223), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G197gat), .ZN(new_n230));
  INV_X1    g029(.A(G204gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT22), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n232), .A2(new_n233), .B1(new_n234), .B2(new_n227), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(new_n223), .A3(new_n227), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n229), .A2(new_n235), .A3(KEYINPUT78), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n227), .A2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT78), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n236), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(new_n228), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n235), .A2(KEYINPUT78), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n244), .A2(KEYINPUT79), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n235), .A2(KEYINPUT78), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n236), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n240), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n249), .B2(new_n237), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n222), .B1(new_n245), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G228gat), .ZN(new_n252));
  INV_X1    g051(.A(G233gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n219), .B1(new_n244), .B2(KEYINPUT29), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n216), .A2(new_n218), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n251), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n254), .B1(new_n251), .B2(new_n258), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n208), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT88), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n244), .A2(KEYINPUT79), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n246), .A3(new_n237), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n221), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT29), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n268), .A3(new_n237), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n256), .B1(new_n269), .B2(new_n219), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n267), .A2(new_n270), .B1(new_n252), .B2(new_n253), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n254), .A3(new_n258), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n207), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(G22gat), .B1(new_n273), .B2(KEYINPUT88), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n259), .A2(new_n260), .A3(new_n208), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n264), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n264), .B2(new_n274), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n219), .B1(new_n216), .B2(new_n218), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n220), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G113gat), .A2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n282), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(KEYINPUT73), .A3(new_n283), .A4(new_n284), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n289), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n283), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n281), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(KEYINPUT5), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT4), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n294), .A2(new_n256), .A3(new_n301), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n291), .A2(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n307), .B1(new_n310), .B2(new_n256), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n303), .B(new_n306), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT83), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n301), .A3(new_n256), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT4), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n315), .A2(new_n308), .B1(new_n302), .B2(new_n281), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT83), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n306), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n305), .B1(new_n281), .B2(new_n302), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n308), .A2(KEYINPUT82), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n315), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n308), .A2(KEYINPUT82), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n302), .A2(new_n257), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n314), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n325), .B1(new_n327), .B2(new_n305), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT0), .ZN(new_n332));
  XNOR2_X1  g131(.A(G57gat), .B(G85gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n334), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n336), .A3(new_n329), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n338), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT85), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n336), .B1(new_n319), .B2(new_n329), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT85), .A3(new_n340), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G8gat), .B(G36gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT23), .ZN(new_n355));
  NAND2_X1  g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT24), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n359), .B1(new_n367), .B2(KEYINPUT65), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n361), .B2(new_n363), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT65), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n353), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n358), .A4(new_n356), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT66), .B(G183gat), .ZN(new_n374));
  INV_X1    g173(.A(G190gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n364), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(KEYINPUT27), .B(G183gat), .Z(new_n378));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n378), .A2(new_n379), .A3(G190gat), .ZN(new_n380));
  AOI21_X1  g179(.A(G190gat), .B1(new_n374), .B2(KEYINPUT27), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n382));
  NOR2_X1   g181(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n383));
  OAI21_X1  g182(.A(G183gat), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT68), .B(G183gat), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n381), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n380), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n391));
  OR3_X1    g190(.A1(new_n391), .A2(new_n354), .A3(KEYINPUT70), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n354), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT70), .B1(new_n391), .B2(new_n354), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n360), .ZN(new_n397));
  OAI22_X1  g196(.A1(new_n372), .A2(new_n377), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n351), .B1(new_n398), .B2(new_n268), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n388), .A2(new_n389), .ZN(new_n400));
  INV_X1    g199(.A(new_n380), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n397), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(G183gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(KEYINPUT24), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n406), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n360), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT65), .B1(new_n407), .B2(new_n365), .ZN(new_n408));
  INV_X1    g207(.A(new_n359), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n371), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n352), .ZN(new_n411));
  INV_X1    g210(.A(new_n377), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n350), .B1(new_n404), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n245), .A2(new_n250), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n399), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n397), .B1(new_n400), .B2(new_n401), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n377), .B1(new_n410), .B2(new_n352), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n268), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n350), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n351), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(KEYINPUT30), .B(new_n349), .C1(new_n416), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n349), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n415), .B1(new_n399), .B2(new_n414), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n417), .A3(new_n422), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n427), .ZN(new_n433));
  XNOR2_X1  g232(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n426), .A2(new_n431), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n279), .B1(new_n346), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n316), .A2(new_n304), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT39), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n334), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n326), .A2(new_n314), .A3(new_n304), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT39), .B(new_n441), .C1(new_n316), .C2(new_n304), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(KEYINPUT40), .A3(new_n442), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n335), .A3(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n436), .A2(new_n447), .A3(KEYINPUT89), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT89), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n435), .A2(new_n432), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n429), .ZN(new_n451));
  AND4_X1   g250(.A1(KEYINPUT80), .A2(new_n451), .A3(KEYINPUT30), .A4(new_n349), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT80), .B1(new_n430), .B2(KEYINPUT30), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n440), .A2(KEYINPUT40), .A3(new_n442), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT40), .B1(new_n440), .B2(new_n442), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n344), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n449), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n275), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n263), .B1(new_n261), .B2(new_n262), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n273), .A2(KEYINPUT88), .A3(G22gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n276), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT37), .B1(new_n416), .B2(new_n423), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n428), .A2(new_n429), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n349), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n432), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n428), .A2(new_n429), .A3(new_n466), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n466), .B1(new_n428), .B2(new_n429), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n427), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(KEYINPUT38), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n339), .A2(new_n343), .A3(new_n345), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n437), .B1(new_n459), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n398), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n404), .A2(new_n413), .A3(KEYINPUT74), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n302), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n398), .A2(new_n480), .A3(new_n310), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G227gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(new_n253), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n479), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT34), .B(new_n487), .C1(new_n483), .C2(new_n484), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n483), .A2(new_n487), .A3(new_n484), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT32), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G15gat), .B(G43gat), .Z(new_n496));
  XNOR2_X1  g295(.A(G71gat), .B(G99gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n492), .B(KEYINPUT32), .C1(new_n494), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n491), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT76), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(new_n491), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n499), .A3(KEYINPUT76), .A4(new_n501), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT75), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n499), .A2(new_n512), .A3(new_n501), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n499), .B2(new_n501), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n502), .A2(KEYINPUT36), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n502), .A2(new_n276), .A3(new_n463), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n346), .A2(new_n436), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT35), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n509), .ZN(new_n523));
  INV_X1    g322(.A(new_n521), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n478), .A2(new_n518), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  OR2_X1    g328(.A1(G43gat), .A2(G50gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G43gat), .A2(G50gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT91), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT91), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n538), .A3(KEYINPUT14), .ZN(new_n539));
  AND2_X1   g338(.A1(KEYINPUT92), .A2(G36gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(KEYINPUT92), .A2(G36gat), .ZN(new_n541));
  OAI21_X1  g340(.A(G29gat), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n537), .B(new_n543), .C1(G29gat), .C2(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n531), .A2(new_n529), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT93), .B(G43gat), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n203), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n533), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n539), .A2(new_n532), .A3(new_n542), .A4(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G1gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT16), .ZN(new_n553));
  INV_X1    g352(.A(G15gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G22gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n263), .A2(G15gat), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(G1gat), .B1(new_n555), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g357(.A(G8gat), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G8gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n560), .B(new_n561), .C1(new_n562), .C2(G1gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT94), .B1(new_n551), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n549), .A2(new_n564), .A3(new_n567), .A4(new_n550), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n572), .A3(new_n550), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n565), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT95), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n569), .A2(new_n574), .A3(new_n578), .A4(new_n570), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G113gat), .B(G141gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G197gat), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT11), .B(G169gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(new_n584), .B(KEYINPUT12), .Z(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n573), .A2(new_n565), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n588), .A2(new_n571), .B1(new_n566), .B2(new_n568), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n569), .A2(new_n574), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT96), .ZN(new_n593));
  INV_X1    g392(.A(new_n551), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n569), .B1(new_n594), .B2(new_n564), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n570), .B(KEYINPUT13), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n528), .B1(new_n587), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n591), .A2(new_n593), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT18), .B1(new_n575), .B2(KEYINPUT95), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n585), .B1(new_n601), .B2(new_n579), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT97), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n580), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n585), .B(KEYINPUT90), .Z(new_n605));
  AOI22_X1  g404(.A1(new_n599), .A2(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G230gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n607), .A2(new_n253), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G57gat), .B(G64gat), .Z(new_n610));
  INV_X1    g409(.A(G71gat), .ZN(new_n611));
  INV_X1    g410(.A(G78gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G71gat), .A2(G78gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G57gat), .B(G64gat), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n614), .B(new_n613), .C1(new_n619), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT7), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT7), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  INV_X1    g426(.A(G85gat), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n627), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n632), .A2(new_n636), .A3(new_n627), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n635), .A2(new_n637), .A3(new_n626), .A4(new_n630), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n626), .B2(new_n630), .ZN(new_n641));
  INV_X1    g440(.A(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n620), .B(new_n618), .C1(new_n641), .C2(new_n642), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n639), .B(KEYINPUT101), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n621), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n641), .A2(new_n642), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .A4(new_n643), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT10), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n638), .A2(new_n634), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n647), .A3(KEYINPUT10), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n609), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n646), .A2(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n608), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G120gat), .B(G148gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n660), .B(new_n665), .ZN(new_n666));
  AND2_X1   g465(.A1(G232gat), .A2(G233gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT41), .ZN(new_n668));
  XNOR2_X1  g467(.A(G134gat), .B(G162gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n594), .A2(new_n652), .B1(KEYINPUT41), .B2(new_n667), .ZN(new_n671));
  INV_X1    g470(.A(new_n652), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n571), .A2(new_n573), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G190gat), .B(G218gat), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n675), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n671), .A2(new_n673), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n670), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n670), .A3(new_n678), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT21), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n621), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(G127gat), .B(G155gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n684), .B(new_n685), .Z(new_n686));
  OAI21_X1  g485(.A(new_n565), .B1(new_n683), .B2(new_n621), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n687), .ZN(new_n689));
  NAND2_X1  g488(.A1(G231gat), .A2(G233gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT98), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(G183gat), .B(G211gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n688), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n695), .B1(new_n688), .B2(new_n689), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n666), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n527), .A2(new_n606), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n476), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  OAI21_X1  g504(.A(G8gat), .B1(new_n705), .B2(new_n436), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT16), .B(G8gat), .Z(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(new_n454), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n709), .A2(KEYINPUT104), .A3(new_n707), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT104), .B1(new_n709), .B2(new_n707), .ZN(new_n711));
  OAI221_X1 g510(.A(new_n706), .B1(new_n707), .B2(new_n709), .C1(new_n710), .C2(new_n711), .ZN(G1325gat));
  OAI21_X1  g511(.A(G15gat), .B1(new_n705), .B2(new_n518), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n702), .A2(new_n554), .A3(new_n523), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1326gat));
  NAND2_X1  g514(.A1(new_n702), .A2(new_n464), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n527), .B2(new_n682), .ZN(new_n720));
  INV_X1    g519(.A(new_n682), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n521), .A2(new_n464), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT89), .B1(new_n436), .B2(new_n447), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n454), .A2(new_n457), .A3(new_n449), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n468), .A2(new_n469), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n473), .A2(KEYINPUT38), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n727), .A3(new_n432), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n279), .B1(new_n728), .B2(new_n346), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n509), .A2(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n524), .A2(new_n515), .A3(new_n519), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT35), .ZN(new_n734));
  AND4_X1   g533(.A1(new_n734), .A2(new_n279), .A3(new_n346), .A4(new_n436), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n733), .A2(KEYINPUT35), .B1(new_n735), .B2(new_n523), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT44), .B(new_n721), .C1(new_n732), .C2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n720), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n606), .A2(new_n698), .A3(new_n666), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(new_n476), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n534), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n527), .A2(new_n682), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n739), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n534), .A3(new_n476), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n743), .A2(new_n748), .ZN(G1328gat));
  NOR4_X1   g548(.A1(new_n745), .A2(new_n436), .A3(new_n541), .A4(new_n540), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n738), .A2(new_n739), .ZN(new_n752));
  OAI22_X1  g551(.A1(new_n752), .A2(new_n436), .B1(new_n541), .B2(new_n540), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1329gat));
  OAI21_X1  g553(.A(new_n547), .B1(new_n745), .B2(new_n509), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n518), .A2(new_n547), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g558(.A1(new_n720), .A2(new_n464), .A3(new_n737), .A4(new_n739), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G50gat), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n279), .A2(G50gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n763), .A3(KEYINPUT48), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n761), .A2(KEYINPUT106), .B1(new_n746), .B2(new_n762), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n760), .A2(new_n767), .A3(G50gat), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n765), .B(KEYINPUT48), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n761), .A2(KEYINPUT106), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n768), .A3(new_n763), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT107), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n764), .B1(new_n769), .B2(new_n773), .ZN(G1331gat));
  INV_X1    g573(.A(new_n527), .ZN(new_n775));
  INV_X1    g574(.A(new_n606), .ZN(new_n776));
  INV_X1    g575(.A(new_n666), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n776), .A2(new_n699), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n476), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g581(.A(new_n436), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT108), .Z(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1333gat));
  NAND3_X1  g586(.A1(new_n780), .A2(G71gat), .A3(new_n731), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT109), .B1(new_n779), .B2(new_n509), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n611), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n779), .A2(KEYINPUT109), .A3(new_n509), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g592(.A1(new_n779), .A2(new_n279), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(new_n612), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n776), .A2(new_n698), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n744), .A2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT51), .B1(new_n744), .B2(new_n796), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n801), .A2(new_n628), .A3(new_n476), .A4(new_n666), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n738), .A2(new_n666), .A3(new_n796), .ZN(new_n803));
  OAI21_X1  g602(.A(G85gat), .B1(new_n803), .B2(new_n346), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1336gat));
  OAI21_X1  g604(.A(G92gat), .B1(new_n803), .B2(new_n436), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(new_n801), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n777), .A2(new_n436), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n629), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT110), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n806), .B(new_n807), .C1(new_n808), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n806), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(new_n807), .ZN(G1337gat));
  NOR2_X1   g615(.A1(new_n509), .A2(G99gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n666), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G99gat), .B1(new_n803), .B2(new_n518), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1338gat));
  NOR2_X1   g619(.A1(new_n279), .A2(G106gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n666), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(G106gat), .B1(new_n803), .B2(new_n279), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n823), .B2(KEYINPUT112), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n822), .B(new_n823), .C1(KEYINPUT112), .C2(new_n825), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1339gat));
  AND2_X1   g628(.A1(new_n606), .A2(new_n700), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n609), .C1(new_n651), .C2(new_n654), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n832), .A2(new_n664), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n608), .B(new_n653), .C1(new_n656), .C2(KEYINPUT10), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n655), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n655), .A2(new_n657), .A3(new_n665), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n599), .A2(new_n603), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n595), .B2(new_n596), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n570), .B2(new_n589), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n595), .A2(new_n842), .A3(new_n596), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n584), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n698), .B1(new_n847), .B2(new_n721), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n587), .A2(new_n528), .A3(new_n598), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT97), .B1(new_n600), .B2(new_n602), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n666), .B(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n838), .A2(new_n839), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n851), .B(new_n682), .C1(new_n606), .C2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n830), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT114), .B(new_n830), .C1(new_n848), .C2(new_n853), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n464), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n509), .A2(new_n346), .A3(new_n454), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n606), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n346), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n520), .A2(new_n454), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n776), .A2(new_n286), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n862), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT115), .ZN(G1340gat));
  NOR3_X1   g667(.A1(new_n861), .A2(new_n287), .A3(new_n777), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n863), .A2(new_n666), .A3(new_n864), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n287), .B2(new_n870), .ZN(G1341gat));
  INV_X1    g670(.A(new_n861), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(G127gat), .A3(new_n698), .ZN(new_n873));
  INV_X1    g672(.A(new_n698), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(KEYINPUT116), .ZN(new_n876));
  AOI21_X1  g675(.A(G127gat), .B1(new_n875), .B2(KEYINPUT116), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(G1342gat));
  OR3_X1    g677(.A1(new_n865), .A2(G134gat), .A3(new_n682), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n872), .A2(new_n721), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n879), .A2(KEYINPUT56), .B1(new_n880), .B2(G134gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(KEYINPUT56), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n879), .A2(new_n884), .A3(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n881), .B1(new_n883), .B2(new_n885), .ZN(G1343gat));
  XNOR2_X1  g685(.A(new_n854), .B(new_n855), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n888), .A3(new_n464), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n731), .A2(new_n346), .A3(new_n454), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT118), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT57), .B1(new_n854), .B2(new_n279), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n606), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n731), .A2(new_n454), .A3(new_n279), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n863), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n606), .A2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(G148gat), .C1(new_n893), .C2(new_n777), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT119), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT57), .B(new_n464), .C1(new_n856), .C2(new_n857), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n888), .B1(new_n854), .B2(new_n279), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n906), .B(new_n888), .C1(new_n854), .C2(new_n279), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n903), .A2(KEYINPUT120), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n909), .A3(KEYINPUT57), .A4(new_n464), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n666), .A3(new_n891), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n900), .B1(new_n912), .B2(G148gat), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n777), .A2(G148gat), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n902), .A2(new_n913), .B1(new_n896), .B2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n893), .B2(new_n874), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n698), .A2(new_n210), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n896), .B2(new_n917), .ZN(G1346gat));
  NOR3_X1   g717(.A1(new_n893), .A2(new_n211), .A3(new_n682), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n863), .A2(new_n721), .A3(new_n895), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n211), .B2(new_n920), .ZN(G1347gat));
  NOR3_X1   g720(.A1(new_n509), .A2(new_n476), .A3(new_n436), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n887), .A2(new_n279), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(G169gat), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n924), .A3(new_n606), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n858), .A2(new_n476), .ZN(new_n926));
  INV_X1    g725(.A(new_n520), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n436), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n776), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n925), .B1(new_n930), .B2(new_n924), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n923), .B2(new_n777), .ZN(new_n932));
  INV_X1    g731(.A(G176gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n809), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n932), .B1(new_n928), .B2(new_n934), .ZN(G1349gat));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(new_n374), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n923), .B2(new_n874), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n874), .A2(new_n378), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n926), .A2(new_n454), .A3(new_n927), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n938), .A2(new_n940), .A3(KEYINPUT122), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n943), .A2(KEYINPUT123), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n946), .B1(new_n941), .B2(KEYINPUT60), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n945), .A2(new_n948), .ZN(G1350gat));
  OAI21_X1  g748(.A(G190gat), .B1(new_n923), .B2(new_n682), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n929), .A2(new_n375), .A3(new_n721), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1351gat));
  NAND3_X1  g752(.A1(new_n518), .A2(new_n346), .A3(new_n454), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n908), .B2(new_n910), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n230), .B1(new_n958), .B2(new_n776), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n731), .A2(new_n436), .A3(new_n279), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n887), .A2(new_n960), .A3(new_n346), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(G197gat), .A3(new_n606), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n959), .A2(KEYINPUT125), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n959), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n666), .A2(new_n231), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n956), .A2(new_n666), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n908), .B2(new_n910), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g770(.A(G204gat), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g771(.A(KEYINPUT126), .B(new_n969), .C1(new_n908), .C2(new_n910), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n968), .B(KEYINPUT127), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1353gat));
  INV_X1    g777(.A(new_n961), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n979), .A2(new_n224), .A3(new_n698), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n954), .A2(new_n874), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n911), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n982), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n983));
  AOI21_X1  g782(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n979), .B2(new_n721), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n682), .A2(new_n225), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n958), .B2(new_n987), .ZN(G1355gat));
endmodule


