//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G134gat), .ZN(new_n209));
  INV_X1    g008(.A(G134gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G127gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G113gat), .B2(G120gat), .ZN(new_n213));
  AND2_X1   g012(.A1(G113gat), .A2(G120gat), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n209), .A2(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(G113gat), .ZN(new_n217));
  INV_X1    g016(.A(G120gat), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT1), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(KEYINPUT68), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G113gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n218), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n215), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT69), .ZN(new_n226));
  XOR2_X1   g025(.A(G141gat), .B(G148gat), .Z(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(KEYINPUT2), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G141gat), .B(G148gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n231), .B(new_n230), .C1(new_n235), .C2(KEYINPUT2), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT68), .B(G113gat), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n219), .B(new_n216), .C1(new_n238), .C2(new_n218), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n215), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT77), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n245), .A3(KEYINPUT4), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n236), .A2(new_n234), .A3(new_n239), .A4(new_n215), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT4), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n244), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n236), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n254), .A3(new_n225), .ZN(new_n255));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n225), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n256), .B1(new_n259), .B2(new_n247), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT78), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n259), .A2(new_n247), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n263), .B(KEYINPUT5), .C1(new_n264), .C2(new_n256), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n250), .A2(new_n258), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n247), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(new_n242), .B2(new_n267), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n261), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n207), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n265), .A2(new_n262), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n248), .B1(new_n243), .B2(KEYINPUT77), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n257), .B1(new_n275), .B2(new_n246), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n206), .B(new_n270), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT6), .B(new_n207), .C1(new_n266), .C2(new_n271), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT85), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283));
  XNOR2_X1  g082(.A(G211gat), .B(G218gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G197gat), .B(G204gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT22), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n287), .A2(KEYINPUT73), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n291), .A2(KEYINPUT73), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(new_n284), .A3(new_n286), .A4(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G226gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n302), .B1(new_n303), .B2(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT23), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n305), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(KEYINPUT23), .B2(new_n303), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n307), .A2(KEYINPUT25), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT24), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT24), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(KEYINPUT65), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  OR3_X1    g115(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n313), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n314), .ZN(new_n320));
  NAND3_X1  g119(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G169gat), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT64), .B1(new_n328), .B2(new_n305), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n303), .A2(new_n302), .A3(KEYINPUT23), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n309), .B(new_n325), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n310), .A2(new_n318), .B1(new_n319), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n303), .A2(KEYINPUT26), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n326), .B2(new_n327), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n311), .B(new_n333), .C1(new_n335), .C2(new_n303), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT28), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT27), .B(G183gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G183gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n323), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n337), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n322), .A2(KEYINPUT27), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n347), .A2(new_n337), .A3(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n336), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n301), .B1(new_n332), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n319), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n318), .A2(KEYINPUT25), .A3(new_n307), .A4(new_n309), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(KEYINPUT67), .ZN(new_n356));
  AOI21_X1  g155(.A(G190gat), .B1(new_n342), .B2(new_n339), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT28), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n358), .B2(new_n348), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(KEYINPUT74), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n300), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n299), .A2(KEYINPUT29), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n332), .B2(new_n350), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n296), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n351), .A2(new_n360), .A3(new_n362), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n354), .A2(new_n299), .A3(new_n359), .ZN(new_n367));
  INV_X1    g166(.A(new_n296), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n283), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n360), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT74), .B1(new_n354), .B2(new_n359), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n299), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n368), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n374), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n374), .A2(KEYINPUT37), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n370), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT38), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n282), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n369), .A3(new_n373), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n369), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n374), .B1(new_n387), .B2(KEYINPUT37), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n366), .A2(new_n296), .A3(new_n367), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n390), .A2(KEYINPUT37), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n368), .B1(new_n361), .B2(new_n364), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT38), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n386), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n388), .C2(new_n370), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n281), .A2(new_n384), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n269), .A2(new_n255), .ZN(new_n397));
  INV_X1    g196(.A(new_n256), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT84), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n397), .A2(KEYINPUT84), .A3(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT39), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n264), .B2(new_n256), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n401), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT84), .B1(new_n397), .B2(new_n398), .ZN(new_n406));
  AOI211_X1 g205(.A(new_n400), .B(new_n256), .C1(new_n269), .C2(new_n255), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n403), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n408), .A3(new_n206), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT40), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n272), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n409), .B2(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n385), .A2(KEYINPUT76), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT76), .B1(new_n385), .B2(new_n414), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT75), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n419), .B1(new_n387), .B2(new_n374), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT75), .B(new_n373), .C1(new_n365), .C2(new_n369), .ZN(new_n421));
  OAI22_X1  g220(.A1(new_n420), .A2(new_n421), .B1(new_n414), .B2(new_n385), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n411), .B(new_n413), .C1(new_n418), .C2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(G228gat), .A2(G233gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n293), .A2(KEYINPUT80), .A3(new_n295), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT29), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n286), .A2(new_n289), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT80), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n284), .A4(new_n294), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n251), .ZN(new_n432));
  INV_X1    g231(.A(new_n295), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT29), .B1(new_n433), .B2(new_n429), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n426), .B1(new_n434), .B2(new_n425), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n253), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n427), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n368), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n424), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT3), .B1(new_n296), .B2(new_n427), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(KEYINPUT82), .A3(new_n253), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n438), .A2(new_n424), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n440), .B2(new_n237), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(G22gat), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n442), .A2(new_n443), .A3(new_n445), .ZN(new_n449));
  INV_X1    g248(.A(new_n438), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n293), .A2(KEYINPUT80), .A3(new_n295), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n430), .A2(new_n427), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT81), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n453), .A2(new_n251), .A3(new_n431), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n450), .B1(new_n454), .B2(new_n253), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n448), .B(new_n449), .C1(new_n455), .C2(new_n424), .ZN(new_n456));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(KEYINPUT31), .B(G50gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  NAND4_X1  g258(.A1(new_n447), .A2(KEYINPUT83), .A3(new_n456), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(new_n459), .B1(new_n456), .B2(new_n447), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n396), .A2(new_n423), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n226), .A2(new_n241), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n467), .B1(new_n332), .B2(new_n350), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n354), .A2(new_n359), .A3(new_n226), .A4(new_n241), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n473));
  NAND2_X1  g272(.A1(KEYINPUT70), .A2(KEYINPUT34), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI22_X1  g274(.A1(new_n470), .A2(new_n472), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n468), .A2(new_n469), .A3(new_n471), .A4(new_n474), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n470), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT32), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G15gat), .B(G43gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G71gat), .B(G99gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n471), .B1(new_n468), .B2(new_n469), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n487), .B2(KEYINPUT33), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT32), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n478), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n486), .A2(new_n491), .A3(new_n478), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n486), .A2(new_n478), .A3(KEYINPUT72), .A4(new_n491), .ZN(new_n496));
  AOI211_X1 g295(.A(KEYINPUT36), .B(new_n492), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n491), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n476), .A2(new_n477), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n488), .A2(new_n490), .ZN(new_n502));
  AOI221_X4 g301(.A(new_n489), .B1(KEYINPUT33), .B2(new_n485), .C1(new_n470), .C2(new_n472), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n498), .B(new_n500), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n495), .A2(new_n496), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n497), .B1(new_n508), .B2(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n380), .A2(KEYINPUT75), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n387), .A2(new_n419), .A3(new_n374), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n510), .A2(new_n511), .B1(new_n386), .B2(KEYINPUT30), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n279), .A2(new_n280), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n385), .A2(new_n414), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n415), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n464), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n460), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n466), .A2(new_n509), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n465), .A2(new_n506), .A3(new_n507), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT35), .B1(new_n523), .B2(new_n518), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n525));
  AOI211_X1 g324(.A(KEYINPUT35), .B(new_n492), .C1(new_n495), .C2(new_n496), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n465), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G50gat), .ZN(new_n532));
  INV_X1    g331(.A(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G43gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  INV_X1    g337(.A(G29gat), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n541), .A2(KEYINPUT89), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n541), .B2(KEYINPUT89), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n537), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT88), .B(G50gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(G43gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT87), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n533), .A3(G43gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n547), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n535), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n543), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g356(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n541), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n536), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n546), .A2(new_n554), .B1(new_n555), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n530), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n542), .ZN(new_n564));
  INV_X1    g363(.A(new_n537), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n554), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n560), .A2(new_n555), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(KEYINPUT90), .A3(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n573), .B(new_n574), .C1(G1gat), .C2(new_n571), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G8gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n568), .ZN(new_n579));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n577), .A2(new_n561), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n580), .B(KEYINPUT13), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n581), .A2(new_n582), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589));
  INV_X1    g388(.A(G197gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT11), .B(G169gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT12), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n576), .B1(new_n563), .B2(new_n569), .ZN(new_n595));
  INV_X1    g394(.A(new_n579), .ZN(new_n596));
  INV_X1    g395(.A(new_n580), .ZN(new_n597));
  NOR3_X1   g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n594), .B1(new_n598), .B2(KEYINPUT18), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n598), .A2(KEYINPUT18), .B1(new_n584), .B2(new_n586), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT92), .B1(new_n598), .B2(KEYINPUT18), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n604), .A3(new_n582), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n594), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n606), .A2(KEYINPUT93), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT93), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n601), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n529), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT94), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n529), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(G85gat), .A2(G92gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT7), .ZN(new_n618));
  NOR2_X1   g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n619), .B1(KEYINPUT8), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G99gat), .B(G106gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n624), .B1(new_n563), .B2(new_n569), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n628));
  INV_X1    g427(.A(new_n624), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n628), .B1(new_n629), .B2(new_n561), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n616), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(KEYINPUT99), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G134gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n229), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n625), .A2(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(new_n616), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n636), .A2(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G57gat), .B(G64gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(G71gat), .A2(G78gat), .ZN(new_n647));
  OAI22_X1  g446(.A1(new_n645), .A2(new_n646), .B1(KEYINPUT95), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(G71gat), .B(G78gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n576), .B1(KEYINPUT21), .B2(new_n650), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G127gat), .B(G155gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n658), .B(KEYINPUT96), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G183gat), .B(G211gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT98), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n655), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G230gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n298), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n622), .A2(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n629), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n624), .A2(new_n650), .A3(new_n668), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n624), .A2(KEYINPUT10), .A3(new_n650), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI211_X1 g474(.A(new_n666), .B(new_n298), .C1(new_n670), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g475(.A(G120gat), .B(G148gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT101), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n675), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(new_n675), .B2(new_n676), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n644), .A2(new_n665), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT102), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n281), .A2(KEYINPUT103), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n513), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n615), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g492(.A1(new_n418), .A2(new_n422), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n686), .B1(new_n612), .B2(new_n614), .ZN(new_n696));
  NAND2_X1  g495(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n697));
  INV_X1    g496(.A(G8gat), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n572), .A2(new_n698), .ZN(new_n699));
  AND4_X1   g498(.A1(new_n695), .A2(new_n696), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n696), .B2(new_n695), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT42), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(KEYINPUT42), .B2(new_n700), .ZN(G1325gat));
  INV_X1    g502(.A(new_n696), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n500), .B1(new_n502), .B2(new_n503), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n507), .A2(new_n705), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n704), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n704), .B2(new_n509), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1326gat));
  NAND3_X1  g508(.A1(new_n615), .A2(new_n520), .A3(new_n687), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT43), .B(G22gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  INV_X1    g511(.A(new_n644), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(new_n664), .A3(new_n684), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n612), .B2(new_n614), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n539), .A3(new_n691), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n529), .A2(new_n644), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n642), .B2(new_n643), .ZN(new_n725));
  INV_X1    g524(.A(new_n643), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(KEYINPUT105), .A3(new_n641), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n522), .B2(new_n528), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n723), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n664), .B(KEYINPUT104), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n606), .A2(new_n607), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n606), .A2(KEYINPUT93), .A3(new_n607), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n600), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n735), .A2(new_n740), .A3(new_n684), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n691), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n721), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G29gat), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n742), .A2(new_n721), .A3(new_n743), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n719), .B(new_n720), .C1(new_n745), .C2(new_n746), .ZN(G1328gat));
  NOR2_X1   g546(.A1(new_n694), .A2(G36gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n716), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n695), .A3(new_n741), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n750), .A2(new_n751), .B1(G36gat), .B2(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n750), .A2(KEYINPUT107), .A3(new_n751), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(G1329gat));
  INV_X1    g556(.A(new_n706), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n716), .A2(new_n531), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n509), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n730), .B1(new_n529), .B2(new_n644), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n760), .B(new_n741), .C1(new_n761), .C2(new_n732), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n764), .B2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n766), .B(new_n767), .C1(new_n759), .C2(new_n763), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n768), .ZN(G1330gat));
  INV_X1    g568(.A(new_n548), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n520), .A2(new_n734), .A3(new_n770), .A4(new_n741), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n716), .B2(new_n520), .ZN(new_n772));
  OR3_X1    g571(.A1(new_n771), .A2(new_n772), .A3(KEYINPUT48), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT48), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1331gat));
  INV_X1    g574(.A(new_n684), .ZN(new_n776));
  NOR4_X1   g575(.A1(new_n610), .A2(new_n644), .A3(new_n665), .A4(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT109), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(new_n529), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n691), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g580(.A(new_n694), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n783), .B(new_n784), .Z(G1333gat));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n760), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n706), .A2(G71gat), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n786), .A2(G71gat), .B1(new_n779), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n520), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n396), .A2(new_n423), .A3(new_n465), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n495), .A2(new_n496), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n705), .A2(KEYINPUT71), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n504), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT36), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT36), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n507), .A2(new_n799), .A3(new_n705), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n521), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n794), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n795), .A2(new_n797), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n803), .A2(new_n525), .A3(new_n465), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT35), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n507), .A2(new_n805), .A3(new_n705), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n520), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n804), .A2(KEYINPUT35), .B1(new_n525), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(KEYINPUT111), .B(new_n644), .C1(new_n802), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n610), .A2(new_n664), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT111), .B1(new_n529), .B2(new_n644), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n793), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n722), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n809), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(KEYINPUT112), .B(new_n793), .C1(new_n811), .C2(new_n812), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n743), .A2(G85gat), .A3(new_n776), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n610), .A2(new_n664), .A3(new_n776), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n723), .B2(new_n733), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825), .B2(new_n743), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n826), .ZN(G1336gat));
  NOR3_X1   g626(.A1(new_n694), .A2(G92gat), .A3(new_n776), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n818), .A2(new_n819), .A3(new_n828), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n695), .B(new_n822), .C1(new_n761), .C2(new_n732), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(new_n830), .B2(G92gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n828), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n813), .B2(new_n816), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n830), .A2(new_n835), .A3(G92gat), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n830), .B2(G92gat), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n834), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n832), .B1(new_n838), .B2(new_n839), .ZN(G1337gat));
  NOR3_X1   g639(.A1(new_n706), .A2(G99gat), .A3(new_n776), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n818), .A2(new_n819), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G99gat), .B1(new_n825), .B2(new_n509), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1338gat));
  NOR3_X1   g643(.A1(new_n465), .A2(G106gat), .A3(new_n776), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n818), .A2(new_n819), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(G106gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n824), .B2(new_n520), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n845), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n813), .B2(new_n816), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n853), .B2(new_n848), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(new_n854), .ZN(G1339gat));
  NAND2_X1  g654(.A1(new_n685), .A2(new_n740), .ZN(new_n856));
  INV_X1    g655(.A(new_n675), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n673), .A2(new_n667), .A3(new_n674), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n680), .B1(new_n675), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(KEYINPUT55), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n682), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n865), .B1(new_n584), .B2(new_n586), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n593), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n859), .A2(new_n861), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT55), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n864), .A2(new_n601), .A3(new_n867), .A4(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n728), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n601), .A2(new_n867), .A3(new_n684), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n864), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n740), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(new_n728), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n856), .B1(new_n876), .B2(new_n735), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n691), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n465), .A2(new_n878), .A3(new_n694), .A4(new_n803), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n238), .A3(new_n610), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n877), .A2(new_n465), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(new_n694), .A3(new_n758), .A4(new_n691), .ZN(new_n882));
  OAI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n740), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(G1340gat));
  NOR3_X1   g683(.A1(new_n882), .A2(new_n218), .A3(new_n776), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n879), .A2(new_n684), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n218), .B2(new_n886), .ZN(G1341gat));
  NAND3_X1  g686(.A1(new_n879), .A2(new_n208), .A3(new_n664), .ZN(new_n888));
  INV_X1    g687(.A(new_n735), .ZN(new_n889));
  OAI21_X1  g688(.A(G127gat), .B1(new_n882), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1342gat));
  NAND3_X1  g690(.A1(new_n879), .A2(new_n210), .A3(new_n644), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n894), .A3(new_n210), .A4(new_n644), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n882), .B2(new_n713), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  NAND3_X1  g696(.A1(new_n509), .A2(new_n694), .A3(new_n691), .ZN(new_n898));
  XNOR2_X1  g697(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n863), .B1(new_n868), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n873), .B1(new_n740), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n872), .B1(new_n902), .B2(new_n713), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n856), .B1(new_n903), .B2(new_n664), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n520), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n898), .B1(new_n905), .B2(KEYINPUT57), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n877), .A2(new_n907), .A3(new_n520), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n610), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n856), .ZN(new_n910));
  INV_X1    g709(.A(new_n873), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n911), .B1(new_n610), .B2(new_n900), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n912), .A2(new_n644), .B1(new_n728), .B2(new_n871), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n665), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT57), .B1(new_n914), .B2(new_n465), .ZN(new_n915));
  INV_X1    g714(.A(new_n898), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n915), .A2(new_n908), .A3(new_n610), .A4(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n909), .A2(new_n919), .A3(G141gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n740), .A2(G141gat), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT116), .Z(new_n922));
  NAND2_X1  g721(.A1(new_n509), .A2(new_n520), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n923), .A2(new_n695), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n877), .A2(new_n922), .A3(new_n691), .A4(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT58), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n917), .A2(G141gat), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT117), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n925), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT58), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n930), .A2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(G148gat), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n878), .A2(new_n936), .A3(new_n684), .A4(new_n924), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n915), .A2(new_n908), .A3(new_n916), .ZN(new_n938));
  AOI211_X1 g737(.A(KEYINPUT59), .B(new_n936), .C1(new_n938), .C2(new_n684), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n940));
  NAND2_X1  g739(.A1(new_n877), .A2(new_n520), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT57), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n686), .A2(new_n610), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n902), .A2(new_n713), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n871), .A2(new_n713), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n664), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n907), .B(new_n520), .C1(new_n943), .C2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n942), .A2(new_n947), .A3(new_n684), .A4(new_n916), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n940), .B1(new_n948), .B2(G148gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n937), .B1(new_n939), .B2(new_n949), .ZN(G1345gat));
  AND3_X1   g749(.A1(new_n878), .A2(new_n664), .A3(new_n924), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G155gat), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n889), .A2(new_n228), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n953), .A2(new_n954), .B1(new_n938), .B2(new_n955), .ZN(G1346gat));
  NAND4_X1  g755(.A1(new_n878), .A2(new_n229), .A3(new_n644), .A4(new_n924), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT122), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n938), .A2(new_n729), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n229), .B2(new_n959), .ZN(G1347gat));
  NAND2_X1  g759(.A1(new_n877), .A2(new_n743), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(new_n694), .A3(new_n523), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n326), .A3(new_n610), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n743), .A2(new_n695), .A3(new_n758), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n881), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n740), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(G1348gat));
  OAI21_X1  g769(.A(G176gat), .B1(new_n966), .B2(new_n776), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n962), .A2(new_n327), .A3(new_n684), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  OAI21_X1  g772(.A(G183gat), .B1(new_n966), .B2(new_n889), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n962), .A2(new_n338), .A3(new_n664), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT60), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT60), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1350gat));
  NAND3_X1  g779(.A1(new_n962), .A2(new_n323), .A3(new_n729), .ZN(new_n981));
  OAI21_X1  g780(.A(G190gat), .B1(new_n966), .B2(new_n713), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n982), .A2(KEYINPUT61), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(G1351gat));
  NOR2_X1   g784(.A1(new_n923), .A2(new_n694), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n877), .A2(new_n743), .A3(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(G197gat), .B1(new_n988), .B2(new_n610), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n942), .A2(new_n947), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n760), .A2(new_n691), .A3(new_n694), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n740), .A2(new_n590), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(G1352gat));
  XNOR2_X1  g794(.A(KEYINPUT125), .B(G204gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n992), .B2(new_n776), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n987), .A2(new_n776), .A3(new_n996), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n999), .ZN(G1353gat));
  OR3_X1    g799(.A1(new_n987), .A2(G211gat), .A3(new_n665), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n942), .A2(new_n947), .A3(new_n664), .A4(new_n991), .ZN(new_n1002));
  AND4_X1   g801(.A1(KEYINPUT126), .A2(new_n1002), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  AOI22_X1  g804(.A1(new_n1002), .A2(new_n1005), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1001), .B1(new_n1003), .B2(new_n1006), .ZN(G1354gat));
  INV_X1    g806(.A(G218gat), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n713), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n987), .B2(new_n728), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(KEYINPUT127), .ZN(new_n1011));
  OR2_X1    g810(.A1(new_n1010), .A2(KEYINPUT127), .ZN(new_n1012));
  AOI22_X1  g811(.A1(new_n993), .A2(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(G1355gat));
endmodule


