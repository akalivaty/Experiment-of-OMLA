

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765;

  XNOR2_X1 U371 ( .A(n573), .B(KEYINPUT35), .ZN(n758) );
  XNOR2_X1 U372 ( .A(n414), .B(n413), .ZN(n577) );
  AND2_X2 U373 ( .A1(n386), .A2(n399), .ZN(n378) );
  AND2_X2 U374 ( .A1(n434), .A2(KEYINPUT92), .ZN(n433) );
  XNOR2_X2 U375 ( .A(n748), .B(n441), .ZN(n726) );
  NOR2_X1 U376 ( .A1(G953), .A2(G237), .ZN(n562) );
  NOR2_X1 U377 ( .A1(n668), .A2(n667), .ZN(n665) );
  BUF_X1 U378 ( .A(G143), .Z(n711) );
  NAND2_X2 U379 ( .A1(n415), .A2(n424), .ZN(n619) );
  XNOR2_X2 U380 ( .A(n499), .B(n498), .ZN(n742) );
  XNOR2_X2 U381 ( .A(n464), .B(n484), .ZN(n499) );
  NAND2_X1 U382 ( .A1(n580), .A2(n583), .ZN(n617) );
  INV_X2 U383 ( .A(G953), .ZN(n394) );
  XNOR2_X1 U384 ( .A(G128), .B(G143), .ZN(n492) );
  XNOR2_X1 U385 ( .A(n591), .B(KEYINPUT110), .ZN(n762) );
  AND2_X1 U386 ( .A1(n621), .A2(n350), .ZN(n375) );
  AND2_X1 U387 ( .A1(n385), .A2(n423), .ZN(n372) );
  XNOR2_X1 U388 ( .A(n532), .B(n456), .ZN(n749) );
  XNOR2_X1 U389 ( .A(n379), .B(KEYINPUT99), .ZN(n464) );
  INV_X1 U390 ( .A(n492), .ZN(n494) );
  XNOR2_X1 U391 ( .A(n457), .B(G125), .ZN(n532) );
  XNOR2_X1 U392 ( .A(G119), .B(KEYINPUT3), .ZN(n379) );
  XNOR2_X1 U393 ( .A(KEYINPUT16), .B(G122), .ZN(n498) );
  XNOR2_X1 U394 ( .A(G137), .B(KEYINPUT70), .ZN(n544) );
  BUF_X1 U395 ( .A(n765), .Z(n348) );
  XNOR2_X2 U396 ( .A(n374), .B(KEYINPUT79), .ZN(n471) );
  AND2_X1 U397 ( .A1(n525), .A2(n401), .ZN(n427) );
  XNOR2_X1 U398 ( .A(n499), .B(n491), .ZN(n497) );
  XNOR2_X1 U399 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U400 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U401 ( .A1(n763), .A2(n706), .ZN(n380) );
  XNOR2_X1 U402 ( .A(n459), .B(KEYINPUT95), .ZN(n458) );
  NAND2_X1 U403 ( .A1(n593), .A2(n592), .ZN(n459) );
  NOR2_X1 U404 ( .A1(n483), .A2(n762), .ZN(n592) );
  INV_X1 U405 ( .A(G146), .ZN(n457) );
  INV_X1 U406 ( .A(n544), .ZN(n417) );
  XOR2_X1 U407 ( .A(n671), .B(KEYINPUT6), .Z(n587) );
  XNOR2_X1 U408 ( .A(n396), .B(KEYINPUT41), .ZN(n678) );
  AND2_X1 U409 ( .A1(n680), .A2(n395), .ZN(n396) );
  NAND2_X1 U410 ( .A1(n376), .A2(n375), .ZN(n374) );
  XNOR2_X1 U411 ( .A(n377), .B(n615), .ZN(n376) );
  NAND2_X1 U412 ( .A1(n402), .A2(n401), .ZN(n400) );
  NOR2_X1 U413 ( .A1(n640), .A2(n363), .ZN(n435) );
  NAND2_X1 U414 ( .A1(n640), .A2(n363), .ZN(n438) );
  NOR2_X1 U415 ( .A1(n390), .A2(n643), .ZN(n479) );
  NOR2_X1 U416 ( .A1(n481), .A2(KEYINPUT92), .ZN(n480) );
  NAND2_X1 U417 ( .A1(n432), .A2(G902), .ZN(n430) );
  NAND2_X1 U418 ( .A1(n401), .A2(G953), .ZN(n519) );
  INV_X1 U419 ( .A(KEYINPUT77), .ZN(n413) );
  NAND2_X1 U420 ( .A1(n619), .A2(n679), .ZN(n377) );
  INV_X1 U421 ( .A(KEYINPUT112), .ZN(n423) );
  XNOR2_X1 U422 ( .A(KEYINPUT90), .B(KEYINPUT45), .ZN(n605) );
  NAND2_X1 U423 ( .A1(n458), .A2(n604), .ZN(n606) );
  XNOR2_X1 U424 ( .A(n565), .B(n420), .ZN(n567) );
  XNOR2_X1 U425 ( .A(n566), .B(n421), .ZN(n420) );
  XNOR2_X1 U426 ( .A(n510), .B(n511), .ZN(n725) );
  XNOR2_X1 U427 ( .A(n546), .B(n742), .ZN(n511) );
  XNOR2_X1 U428 ( .A(n389), .B(n359), .ZN(n409) );
  NAND2_X1 U429 ( .A1(n471), .A2(n680), .ZN(n389) );
  XNOR2_X1 U430 ( .A(n383), .B(n517), .ZN(n412) );
  XNOR2_X1 U431 ( .A(n516), .B(KEYINPUT68), .ZN(n517) );
  NOR2_X1 U432 ( .A1(n634), .A2(n384), .ZN(n383) );
  NAND2_X1 U433 ( .A1(n398), .A2(n401), .ZN(n397) );
  NAND2_X1 U434 ( .A1(n587), .A2(KEYINPUT94), .ZN(n467) );
  XNOR2_X1 U435 ( .A(n586), .B(n470), .ZN(n597) );
  OR2_X1 U436 ( .A1(n587), .A2(KEYINPUT94), .ZN(n469) );
  XNOR2_X1 U437 ( .A(n453), .B(n362), .ZN(n452) );
  INV_X1 U438 ( .A(G898), .ZN(n393) );
  INV_X1 U439 ( .A(G952), .ZN(n392) );
  NOR2_X1 U440 ( .A1(n696), .A2(n405), .ZN(n404) );
  INV_X1 U441 ( .A(n525), .ZN(n432) );
  XNOR2_X1 U442 ( .A(G101), .B(G146), .ZN(n488) );
  INV_X1 U443 ( .A(KEYINPUT5), .ZN(n487) );
  XOR2_X1 U444 ( .A(G137), .B(KEYINPUT105), .Z(n486) );
  OR2_X1 U445 ( .A1(G237), .A2(G902), .ZN(n515) );
  XNOR2_X1 U446 ( .A(G113), .B(G131), .ZN(n566) );
  INV_X1 U447 ( .A(KEYINPUT108), .ZN(n421) );
  XOR2_X1 U448 ( .A(KEYINPUT12), .B(G104), .Z(n560) );
  INV_X1 U449 ( .A(G140), .ZN(n547) );
  XNOR2_X1 U450 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U451 ( .A(KEYINPUT80), .ZN(n501) );
  NAND2_X1 U452 ( .A1(n394), .A2(G224), .ZN(n502) );
  XNOR2_X1 U453 ( .A(KEYINPUT97), .B(KEYINPUT17), .ZN(n504) );
  XOR2_X1 U454 ( .A(KEYINPUT18), .B(KEYINPUT100), .Z(n505) );
  XNOR2_X1 U455 ( .A(n741), .B(n418), .ZN(n546) );
  XNOR2_X1 U456 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n418) );
  INV_X1 U457 ( .A(KEYINPUT4), .ZN(n495) );
  NOR2_X1 U458 ( .A1(n479), .A2(n724), .ZN(n478) );
  AND2_X1 U459 ( .A1(n668), .A2(n454), .ZN(n618) );
  NOR2_X1 U460 ( .A1(n667), .A2(n455), .ZN(n454) );
  INV_X1 U461 ( .A(n355), .ZN(n455) );
  INV_X1 U462 ( .A(G469), .ZN(n398) );
  XOR2_X1 U463 ( .A(n647), .B(KEYINPUT67), .Z(n648) );
  XNOR2_X1 U464 ( .A(G110), .B(KEYINPUT23), .ZN(n537) );
  XOR2_X1 U465 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n538) );
  XNOR2_X1 U466 ( .A(G119), .B(G128), .ZN(n533) );
  XNOR2_X1 U467 ( .A(G140), .B(KEYINPUT10), .ZN(n456) );
  XNOR2_X1 U468 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n536) );
  XNOR2_X1 U469 ( .A(G116), .B(G134), .ZN(n550) );
  XOR2_X1 U470 ( .A(G107), .B(G122), .Z(n551) );
  XNOR2_X1 U471 ( .A(n546), .B(n442), .ZN(n441) );
  XNOR2_X1 U472 ( .A(n545), .B(n443), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n547), .B(G146), .ZN(n443) );
  XNOR2_X1 U474 ( .A(n403), .B(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U475 ( .A1(n577), .A2(n610), .ZN(n403) );
  INV_X1 U476 ( .A(KEYINPUT106), .ZN(n448) );
  NOR2_X1 U477 ( .A1(n577), .A2(n576), .ZN(n449) );
  AND2_X1 U478 ( .A1(n425), .A2(n426), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n569), .B(n422), .ZN(n582) );
  XNOR2_X1 U480 ( .A(n570), .B(G475), .ZN(n422) );
  NAND2_X1 U481 ( .A1(n412), .A2(n411), .ZN(n523) );
  NOR2_X1 U482 ( .A1(n522), .A2(n361), .ZN(n411) );
  OR2_X2 U483 ( .A1(n678), .A2(n628), .ZN(n623) );
  XNOR2_X1 U484 ( .A(n388), .B(n387), .ZN(n765) );
  INV_X1 U485 ( .A(KEYINPUT40), .ZN(n387) );
  XNOR2_X1 U486 ( .A(n416), .B(n360), .ZN(n626) );
  NOR2_X1 U487 ( .A1(n625), .A2(n634), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n382), .B(n596), .ZN(n763) );
  NOR2_X1 U489 ( .A1(n468), .A2(n465), .ZN(n591) );
  NOR2_X1 U490 ( .A1(n597), .A2(n469), .ZN(n468) );
  XNOR2_X1 U491 ( .A(n451), .B(n368), .ZN(G57) );
  NAND2_X1 U492 ( .A1(n452), .A2(n369), .ZN(n451) );
  AND2_X1 U493 ( .A1(n393), .A2(G953), .ZN(n744) );
  INV_X1 U494 ( .A(KEYINPUT60), .ZN(n460) );
  INV_X1 U495 ( .A(KEYINPUT56), .ZN(n472) );
  NAND2_X1 U496 ( .A1(n406), .A2(n404), .ZN(n700) );
  XOR2_X1 U497 ( .A(G104), .B(G107), .Z(n349) );
  AND2_X1 U498 ( .A1(n665), .A2(n355), .ZN(n350) );
  AND2_X1 U499 ( .A1(n431), .A2(n430), .ZN(n351) );
  OR2_X1 U500 ( .A1(n726), .A2(n397), .ZN(n352) );
  XNOR2_X1 U501 ( .A(n513), .B(n512), .ZN(n353) );
  NOR2_X1 U502 ( .A1(n597), .A2(n587), .ZN(n354) );
  XOR2_X1 U503 ( .A(KEYINPUT84), .B(n609), .Z(n355) );
  XOR2_X1 U504 ( .A(G131), .B(G134), .Z(n356) );
  AND2_X1 U505 ( .A1(n590), .A2(n467), .ZN(n357) );
  AND2_X1 U506 ( .A1(n427), .A2(KEYINPUT112), .ZN(n358) );
  XNOR2_X1 U507 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n359) );
  XNOR2_X1 U508 ( .A(KEYINPUT36), .B(KEYINPUT115), .ZN(n360) );
  NAND2_X1 U509 ( .A1(G214), .A2(n515), .ZN(n679) );
  AND2_X1 U510 ( .A1(G898), .A2(G953), .ZN(n361) );
  INV_X1 U511 ( .A(G902), .ZN(n401) );
  XOR2_X1 U512 ( .A(n371), .B(KEYINPUT62), .Z(n362) );
  XNOR2_X1 U513 ( .A(n642), .B(KEYINPUT48), .ZN(n363) );
  XNOR2_X1 U514 ( .A(n496), .B(n417), .ZN(n748) );
  XNOR2_X1 U515 ( .A(n731), .B(KEYINPUT123), .ZN(n364) );
  XOR2_X1 U516 ( .A(n656), .B(n655), .Z(n365) );
  XOR2_X1 U517 ( .A(n725), .B(n482), .Z(n366) );
  XOR2_X1 U518 ( .A(n728), .B(n727), .Z(n367) );
  XOR2_X1 U519 ( .A(G902), .B(KEYINPUT15), .Z(n646) );
  XOR2_X1 U520 ( .A(n653), .B(KEYINPUT98), .Z(n368) );
  NAND2_X1 U521 ( .A1(n392), .A2(G953), .ZN(n369) );
  BUF_X1 U522 ( .A(n471), .Z(n370) );
  INV_X1 U523 ( .A(n428), .ZN(n371) );
  XNOR2_X1 U524 ( .A(n496), .B(n497), .ZN(n524) );
  NAND2_X1 U525 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U526 ( .A1(n428), .A2(n427), .ZN(n373) );
  NAND2_X1 U527 ( .A1(n428), .A2(n427), .ZN(n385) );
  NAND2_X1 U528 ( .A1(n621), .A2(n665), .ZN(n614) );
  NAND2_X2 U529 ( .A1(n378), .A2(n352), .ZN(n621) );
  XNOR2_X1 U530 ( .A(n380), .B(n600), .ZN(n603) );
  NAND2_X1 U531 ( .A1(n381), .A2(n668), .ZN(n706) );
  XNOR2_X1 U532 ( .A(n599), .B(KEYINPUT65), .ZN(n381) );
  NAND2_X1 U533 ( .A1(n354), .A2(n595), .ZN(n382) );
  INV_X1 U534 ( .A(n634), .ZN(n391) );
  INV_X1 U535 ( .A(n412), .ZN(n629) );
  INV_X1 U536 ( .A(n679), .ZN(n384) );
  NAND2_X1 U537 ( .A1(n351), .A2(n373), .ZN(n671) );
  NAND2_X1 U538 ( .A1(n726), .A2(G469), .ZN(n386) );
  NAND2_X1 U539 ( .A1(n409), .A2(n407), .ZN(n388) );
  NAND2_X1 U540 ( .A1(G902), .A2(G469), .ZN(n399) );
  OR2_X1 U541 ( .A1(n613), .A2(n391), .ZN(n390) );
  XNOR2_X2 U542 ( .A(n514), .B(n353), .ZN(n634) );
  NAND2_X1 U543 ( .A1(n394), .A2(G234), .ZN(n535) );
  AND2_X1 U544 ( .A1(n394), .A2(G227), .ZN(n545) );
  NAND2_X1 U545 ( .A1(n697), .A2(n394), .ZN(n405) );
  NAND2_X1 U546 ( .A1(n736), .A2(n394), .ZN(n740) );
  NAND2_X1 U547 ( .A1(n752), .A2(n394), .ZN(n757) );
  NAND2_X1 U548 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U549 ( .A1(n682), .A2(n384), .ZN(n395) );
  XNOR2_X2 U550 ( .A(n400), .B(n543), .ZN(n668) );
  INV_X1 U551 ( .A(n735), .ZN(n402) );
  NOR2_X1 U552 ( .A1(n688), .A2(n585), .ZN(n548) );
  NAND2_X1 U553 ( .A1(n663), .A2(n662), .ZN(n406) );
  INV_X1 U554 ( .A(n617), .ZN(n407) );
  AND2_X1 U555 ( .A1(n409), .A2(n408), .ZN(n724) );
  INV_X1 U556 ( .A(n718), .ZN(n408) );
  NOR2_X2 U557 ( .A1(n765), .A2(n760), .ZN(n410) );
  AND2_X2 U558 ( .A1(n657), .A2(n662), .ZN(n729) );
  NOR2_X2 U559 ( .A1(n477), .A2(n476), .ZN(n658) );
  NAND2_X1 U560 ( .A1(n649), .A2(n648), .ZN(n657) );
  NAND2_X1 U561 ( .A1(n440), .A2(n478), .ZN(n477) );
  NAND2_X1 U562 ( .A1(n733), .A2(G217), .ZN(n734) );
  BUF_X2 U563 ( .A(n729), .Z(n733) );
  NAND2_X1 U564 ( .A1(n436), .A2(n435), .ZN(n434) );
  XNOR2_X1 U565 ( .A(n410), .B(KEYINPUT46), .ZN(n632) );
  NAND2_X1 U566 ( .A1(n729), .A2(G475), .ZN(n463) );
  NOR2_X1 U567 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U568 ( .A1(n588), .A2(n665), .ZN(n414) );
  AND2_X2 U569 ( .A1(n450), .A2(n480), .ZN(n476) );
  NAND2_X1 U570 ( .A1(n372), .A2(n351), .ZN(n415) );
  XNOR2_X1 U571 ( .A(n621), .B(KEYINPUT1), .ZN(n588) );
  XNOR2_X2 U572 ( .A(n508), .B(n356), .ZN(n496) );
  NOR2_X1 U573 ( .A1(n645), .A2(n526), .ZN(n447) );
  NAND2_X1 U574 ( .A1(n729), .A2(G210), .ZN(n475) );
  NAND2_X1 U575 ( .A1(n447), .A2(n736), .ZN(n649) );
  NOR2_X1 U576 ( .A1(n419), .A2(n610), .ZN(n611) );
  NAND2_X1 U577 ( .A1(n712), .A2(n618), .ZN(n419) );
  NAND2_X1 U578 ( .A1(n437), .A2(n433), .ZN(n440) );
  XNOR2_X2 U579 ( .A(n553), .B(n495), .ZN(n508) );
  XNOR2_X2 U580 ( .A(n494), .B(n493), .ZN(n553) );
  NAND2_X1 U581 ( .A1(n428), .A2(n358), .ZN(n426) );
  NAND2_X1 U582 ( .A1(n429), .A2(KEYINPUT112), .ZN(n425) );
  INV_X1 U583 ( .A(n524), .ZN(n428) );
  NAND2_X1 U584 ( .A1(n524), .A2(n432), .ZN(n431) );
  NAND2_X1 U585 ( .A1(n437), .A2(n434), .ZN(n450) );
  INV_X1 U586 ( .A(n641), .ZN(n436) );
  AND2_X2 U587 ( .A1(n439), .A2(n438), .ZN(n437) );
  NAND2_X1 U588 ( .A1(n641), .A2(n363), .ZN(n439) );
  XNOR2_X1 U589 ( .A(n463), .B(n365), .ZN(n462) );
  XNOR2_X1 U590 ( .A(n475), .B(n366), .ZN(n474) );
  AND2_X1 U591 ( .A1(n444), .A2(n369), .ZN(G54) );
  XNOR2_X1 U592 ( .A(n730), .B(n367), .ZN(n444) );
  AND2_X1 U593 ( .A1(n445), .A2(n369), .ZN(G63) );
  XNOR2_X1 U594 ( .A(n732), .B(n364), .ZN(n445) );
  AND2_X1 U595 ( .A1(n446), .A2(n369), .ZN(G66) );
  XNOR2_X1 U596 ( .A(n734), .B(n402), .ZN(n446) );
  NAND2_X1 U597 ( .A1(n462), .A2(n369), .ZN(n461) );
  NAND2_X1 U598 ( .A1(n474), .A2(n369), .ZN(n473) );
  NAND2_X1 U599 ( .A1(n717), .A2(n702), .ZN(n581) );
  XNOR2_X1 U600 ( .A(n578), .B(KEYINPUT31), .ZN(n717) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(G51) );
  XNOR2_X1 U602 ( .A(n449), .B(n448), .ZN(n675) );
  NAND2_X1 U603 ( .A1(n652), .A2(n657), .ZN(n453) );
  XNOR2_X1 U604 ( .A(n461), .B(n460), .ZN(G60) );
  NAND2_X1 U605 ( .A1(n466), .A2(n357), .ZN(n465) );
  NAND2_X1 U606 ( .A1(n597), .A2(KEYINPUT94), .ZN(n466) );
  INV_X1 U607 ( .A(KEYINPUT22), .ZN(n470) );
  XNOR2_X2 U608 ( .A(KEYINPUT64), .B(KEYINPUT83), .ZN(n493) );
  NAND2_X1 U609 ( .A1(n370), .A2(n635), .ZN(n710) );
  INV_X1 U610 ( .A(n390), .ZN(n481) );
  XNOR2_X1 U611 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n482) );
  AND2_X1 U612 ( .A1(n581), .A2(n683), .ZN(n483) );
  INV_X1 U613 ( .A(KEYINPUT78), .ZN(n644) );
  XNOR2_X1 U614 ( .A(n503), .B(n532), .ZN(n507) );
  XNOR2_X1 U615 ( .A(KEYINPUT38), .B(KEYINPUT76), .ZN(n616) );
  INV_X1 U616 ( .A(KEYINPUT30), .ZN(n615) );
  BUF_X1 U617 ( .A(n658), .Z(n750) );
  XNOR2_X1 U618 ( .A(n540), .B(n539), .ZN(n541) );
  INV_X1 U619 ( .A(KEYINPUT63), .ZN(n653) );
  XNOR2_X1 U620 ( .A(n542), .B(n541), .ZN(n735) );
  XNOR2_X1 U621 ( .A(n700), .B(n699), .ZN(G75) );
  XNOR2_X1 U622 ( .A(G116), .B(G113), .ZN(n484) );
  NAND2_X1 U623 ( .A1(n562), .A2(G210), .ZN(n485) );
  XNOR2_X1 U624 ( .A(n486), .B(n485), .ZN(n490) );
  INV_X1 U625 ( .A(n646), .ZN(n526) );
  XNOR2_X1 U626 ( .A(G101), .B(G110), .ZN(n500) );
  XNOR2_X1 U627 ( .A(n349), .B(n500), .ZN(n741) );
  XNOR2_X1 U628 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U629 ( .A(n507), .B(n506), .Z(n509) );
  XNOR2_X1 U630 ( .A(n508), .B(n509), .ZN(n510) );
  NAND2_X1 U631 ( .A1(n526), .A2(n725), .ZN(n514) );
  XOR2_X1 U632 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n513) );
  NAND2_X1 U633 ( .A1(G210), .A2(n515), .ZN(n512) );
  INV_X1 U634 ( .A(KEYINPUT19), .ZN(n516) );
  NAND2_X1 U635 ( .A1(G234), .A2(G237), .ZN(n518) );
  XNOR2_X1 U636 ( .A(n518), .B(KEYINPUT14), .ZN(n693) );
  NAND2_X1 U637 ( .A1(n693), .A2(n519), .ZN(n521) );
  NOR2_X1 U638 ( .A1(G953), .A2(G952), .ZN(n520) );
  NOR2_X1 U639 ( .A1(n521), .A2(n520), .ZN(n608) );
  INV_X1 U640 ( .A(n608), .ZN(n522) );
  XNOR2_X2 U641 ( .A(n523), .B(KEYINPUT0), .ZN(n585) );
  XNOR2_X1 U642 ( .A(G472), .B(KEYINPUT75), .ZN(n525) );
  INV_X1 U643 ( .A(n587), .ZN(n610) );
  NAND2_X1 U644 ( .A1(n526), .A2(G234), .ZN(n527) );
  XNOR2_X1 U645 ( .A(n527), .B(KEYINPUT20), .ZN(n529) );
  NAND2_X1 U646 ( .A1(n529), .A2(G221), .ZN(n528) );
  XNOR2_X1 U647 ( .A(KEYINPUT21), .B(n528), .ZN(n667) );
  XOR2_X1 U648 ( .A(KEYINPUT103), .B(KEYINPUT25), .Z(n531) );
  NAND2_X1 U649 ( .A1(G217), .A2(n529), .ZN(n530) );
  XNOR2_X1 U650 ( .A(n531), .B(n530), .ZN(n543) );
  XOR2_X1 U651 ( .A(n533), .B(n544), .Z(n534) );
  XNOR2_X1 U652 ( .A(n749), .B(n534), .ZN(n542) );
  XNOR2_X1 U653 ( .A(n536), .B(n535), .ZN(n549) );
  NAND2_X1 U654 ( .A1(n549), .A2(G221), .ZN(n540) );
  XNOR2_X1 U655 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U656 ( .A(n548), .B(KEYINPUT34), .ZN(n572) );
  NAND2_X1 U657 ( .A1(n549), .A2(G217), .ZN(n557) );
  XNOR2_X1 U658 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U659 ( .A(n552), .B(KEYINPUT7), .Z(n555) );
  XNOR2_X1 U660 ( .A(n553), .B(KEYINPUT9), .ZN(n554) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U662 ( .A(n557), .B(n556), .ZN(n731) );
  NOR2_X1 U663 ( .A1(G902), .A2(n731), .ZN(n558) );
  XOR2_X1 U664 ( .A(G478), .B(n558), .Z(n579) );
  XNOR2_X1 U665 ( .A(KEYINPUT109), .B(KEYINPUT13), .ZN(n570) );
  XNOR2_X1 U666 ( .A(n711), .B(G122), .ZN(n559) );
  XNOR2_X1 U667 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U668 ( .A(n749), .B(n561), .ZN(n568) );
  XOR2_X1 U669 ( .A(KEYINPUT107), .B(KEYINPUT11), .Z(n564) );
  NAND2_X1 U670 ( .A1(G214), .A2(n562), .ZN(n563) );
  XNOR2_X1 U671 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U672 ( .A(n568), .B(n567), .ZN(n654) );
  NOR2_X1 U673 ( .A1(G902), .A2(n654), .ZN(n569) );
  INV_X1 U674 ( .A(n582), .ZN(n580) );
  NAND2_X1 U675 ( .A1(n579), .A2(n580), .ZN(n633) );
  XNOR2_X1 U676 ( .A(KEYINPUT81), .B(n633), .ZN(n571) );
  NAND2_X1 U677 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U678 ( .A1(n758), .A2(KEYINPUT44), .ZN(n593) );
  NOR2_X1 U679 ( .A1(n585), .A2(n614), .ZN(n574) );
  XNOR2_X1 U680 ( .A(n574), .B(KEYINPUT104), .ZN(n575) );
  INV_X1 U681 ( .A(n671), .ZN(n576) );
  NAND2_X1 U682 ( .A1(n575), .A2(n576), .ZN(n702) );
  NOR2_X1 U683 ( .A1(n675), .A2(n585), .ZN(n578) );
  NAND2_X1 U684 ( .A1(n579), .A2(n582), .ZN(n718) );
  INV_X1 U685 ( .A(n579), .ZN(n583) );
  NAND2_X1 U686 ( .A1(n718), .A2(n617), .ZN(n683) );
  NAND2_X1 U687 ( .A1(n583), .A2(n582), .ZN(n682) );
  OR2_X1 U688 ( .A1(n682), .A2(n667), .ZN(n584) );
  BUF_X1 U689 ( .A(n588), .Z(n664) );
  INV_X1 U690 ( .A(n664), .ZN(n627) );
  INV_X1 U691 ( .A(n668), .ZN(n589) );
  AND2_X1 U692 ( .A1(n627), .A2(n589), .ZN(n590) );
  INV_X1 U693 ( .A(KEYINPUT44), .ZN(n601) );
  NAND2_X1 U694 ( .A1(KEYINPUT96), .A2(n601), .ZN(n600) );
  XNOR2_X1 U695 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n596) );
  NAND2_X1 U696 ( .A1(n668), .A2(n664), .ZN(n594) );
  XNOR2_X1 U697 ( .A(KEYINPUT111), .B(n594), .ZN(n595) );
  NOR2_X1 U698 ( .A1(n597), .A2(n619), .ZN(n598) );
  NAND2_X1 U699 ( .A1(n627), .A2(n598), .ZN(n599) );
  NAND2_X1 U700 ( .A1(n758), .A2(n601), .ZN(n602) );
  NAND2_X1 U701 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X2 U702 ( .A(n606), .B(n605), .ZN(n736) );
  NAND2_X1 U703 ( .A1(G953), .A2(G900), .ZN(n607) );
  NAND2_X1 U704 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U705 ( .A(KEYINPUT113), .B(n617), .ZN(n712) );
  NAND2_X1 U706 ( .A1(n611), .A2(n679), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n664), .A2(n625), .ZN(n612) );
  XNOR2_X1 U708 ( .A(n612), .B(KEYINPUT43), .ZN(n613) );
  XNOR2_X2 U709 ( .A(n634), .B(n616), .ZN(n680) );
  XOR2_X1 U710 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n624) );
  AND2_X1 U711 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U712 ( .A(KEYINPUT28), .B(n620), .ZN(n622) );
  NAND2_X1 U713 ( .A1(n622), .A2(n621), .ZN(n628) );
  XNOR2_X1 U714 ( .A(n624), .B(n623), .ZN(n760) );
  NOR2_X1 U715 ( .A1(n627), .A2(n626), .ZN(n721) );
  NOR2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n713) );
  NAND2_X1 U717 ( .A1(n713), .A2(n683), .ZN(n636) );
  NOR2_X1 U718 ( .A1(KEYINPUT47), .A2(n636), .ZN(n630) );
  NOR2_X1 U719 ( .A1(n721), .A2(n630), .ZN(n631) );
  NAND2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n641) );
  NOR2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U722 ( .A(n710), .B(KEYINPUT88), .ZN(n638) );
  NAND2_X1 U723 ( .A1(KEYINPUT47), .A2(n636), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U725 ( .A(n639), .B(KEYINPUT87), .Z(n640) );
  XOR2_X1 U726 ( .A(KEYINPUT71), .B(KEYINPUT93), .Z(n642) );
  INV_X1 U727 ( .A(KEYINPUT92), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n658), .B(n644), .ZN(n645) );
  NAND2_X1 U729 ( .A1(KEYINPUT2), .A2(n646), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n658), .A2(KEYINPUT2), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n650), .B(KEYINPUT91), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n651), .A2(n736), .ZN(n662) );
  AND2_X1 U733 ( .A1(G472), .A2(n662), .ZN(n652) );
  XOR2_X1 U734 ( .A(KEYINPUT59), .B(KEYINPUT122), .Z(n656) );
  XNOR2_X1 U735 ( .A(n654), .B(KEYINPUT66), .ZN(n655) );
  OR2_X1 U736 ( .A1(n678), .A2(n688), .ZN(n697) );
  XNOR2_X1 U737 ( .A(KEYINPUT86), .B(KEYINPUT2), .ZN(n660) );
  AND2_X1 U738 ( .A1(n736), .A2(n750), .ZN(n659) );
  NOR2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n661), .B(KEYINPUT85), .ZN(n663) );
  NOR2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U742 ( .A(KEYINPUT50), .B(n666), .Z(n673) );
  NAND2_X1 U743 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(KEYINPUT49), .ZN(n670) );
  NOR2_X1 U745 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(KEYINPUT51), .B(n676), .ZN(n677) );
  NOR2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n691) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n687) );
  INV_X1 U752 ( .A(n683), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U757 ( .A(KEYINPUT52), .B(n692), .ZN(n695) );
  NAND2_X1 U758 ( .A1(n693), .A2(G952), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n695), .A2(n694), .ZN(n696) );
  INV_X1 U760 ( .A(KEYINPUT53), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT120), .ZN(n699) );
  INV_X1 U762 ( .A(n712), .ZN(n715) );
  NOR2_X1 U763 ( .A1(n702), .A2(n715), .ZN(n701) );
  XOR2_X1 U764 ( .A(G104), .B(n701), .Z(G6) );
  NOR2_X1 U765 ( .A1(n718), .A2(n702), .ZN(n704) );
  XNOR2_X1 U766 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n703) );
  XNOR2_X1 U767 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U768 ( .A(G107), .B(n705), .ZN(G9) );
  XNOR2_X1 U769 ( .A(G110), .B(n706), .ZN(G12) );
  XOR2_X1 U770 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n708) );
  NAND2_X1 U771 ( .A1(n713), .A2(n408), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n708), .B(n707), .ZN(n709) );
  XOR2_X1 U773 ( .A(G128), .B(n709), .Z(G30) );
  XNOR2_X1 U774 ( .A(n711), .B(n710), .ZN(G45) );
  NAND2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U776 ( .A(n714), .B(G146), .ZN(G48) );
  NOR2_X1 U777 ( .A1(n717), .A2(n715), .ZN(n716) );
  XOR2_X1 U778 ( .A(G113), .B(n716), .Z(G15) );
  NOR2_X1 U779 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U780 ( .A(KEYINPUT118), .B(n719), .Z(n720) );
  XNOR2_X1 U781 ( .A(G116), .B(n720), .ZN(G18) );
  XOR2_X1 U782 ( .A(KEYINPUT119), .B(KEYINPUT37), .Z(n723) );
  XNOR2_X1 U783 ( .A(G125), .B(n721), .ZN(n722) );
  XNOR2_X1 U784 ( .A(n723), .B(n722), .ZN(G27) );
  XOR2_X1 U785 ( .A(G134), .B(n724), .Z(G36) );
  XOR2_X1 U786 ( .A(G140), .B(n481), .Z(G42) );
  XNOR2_X1 U787 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n728) );
  XNOR2_X1 U788 ( .A(n726), .B(KEYINPUT57), .ZN(n727) );
  NAND2_X1 U789 ( .A1(n733), .A2(G469), .ZN(n730) );
  NAND2_X1 U790 ( .A1(n733), .A2(G478), .ZN(n732) );
  NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U792 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n738), .A2(G898), .ZN(n739) );
  NAND2_X1 U794 ( .A1(n740), .A2(n739), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n741), .B(n742), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n743), .B(KEYINPUT124), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(G69) );
  XOR2_X1 U799 ( .A(n749), .B(n748), .Z(n753) );
  INV_X1 U800 ( .A(n753), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U802 ( .A(G227), .B(n753), .ZN(n754) );
  NAND2_X1 U803 ( .A1(n754), .A2(G900), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(G953), .ZN(n756) );
  NAND2_X1 U805 ( .A1(n757), .A2(n756), .ZN(G72) );
  XNOR2_X1 U806 ( .A(n758), .B(G122), .ZN(n759) );
  XNOR2_X1 U807 ( .A(n759), .B(KEYINPUT125), .ZN(G24) );
  XOR2_X1 U808 ( .A(n760), .B(G137), .Z(G39) );
  XOR2_X1 U809 ( .A(G101), .B(KEYINPUT116), .Z(n761) );
  XNOR2_X1 U810 ( .A(n762), .B(n761), .ZN(G3) );
  XNOR2_X1 U811 ( .A(G119), .B(KEYINPUT126), .ZN(n764) );
  XNOR2_X1 U812 ( .A(n764), .B(n763), .ZN(G21) );
  XOR2_X1 U813 ( .A(n348), .B(G131), .Z(G33) );
endmodule

