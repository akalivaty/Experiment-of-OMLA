//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n188), .A2(new_n189), .A3(G143), .A4(G214), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n187), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n187), .A3(new_n193), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT17), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(KEYINPUT88), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G125), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n200), .A2(KEYINPUT16), .A3(G140), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(KEYINPUT16), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n194), .A2(KEYINPUT17), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT88), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n199), .A2(new_n207), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G113), .B(G122), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT87), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(G104), .ZN(new_n214));
  XOR2_X1   g028(.A(G125), .B(G140), .Z(new_n215));
  OAI21_X1  g029(.A(KEYINPUT72), .B1(new_n215), .B2(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT72), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n202), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(G146), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n220), .A2(new_n221), .B1(KEYINPUT18), .B2(new_n194), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n192), .B(new_n193), .C1(new_n223), .C2(new_n187), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT85), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT86), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT86), .B1(new_n222), .B2(new_n225), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n211), .B(new_n214), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n215), .B(KEYINPUT19), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n205), .B1(new_n229), .B2(G146), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(new_n197), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n225), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT86), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n236), .B2(new_n214), .ZN(new_n237));
  INV_X1    g051(.A(G475), .ZN(new_n238));
  INV_X1    g052(.A(G902), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n235), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n214), .B1(new_n243), .B2(new_n211), .ZN(new_n244));
  INV_X1    g058(.A(new_n228), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n239), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G475), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n237), .A2(KEYINPUT20), .A3(new_n238), .A4(new_n239), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G952), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(G234), .A2(G237), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT21), .B(G898), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n252), .A2(G902), .A3(G953), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT9), .B(G234), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(new_n261), .A3(G953), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G122), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G116), .ZN(new_n265));
  INV_X1    g079(.A(G116), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G122), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT14), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(KEYINPUT14), .A3(G122), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(G107), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G107), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT65), .B(G128), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n275), .B(new_n278), .C1(new_n279), .C2(new_n191), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(KEYINPUT65), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT65), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G128), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n191), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G134), .B1(new_n284), .B2(new_n277), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n274), .B1(new_n280), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT13), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n276), .B2(G143), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n191), .A2(KEYINPUT13), .A3(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G134), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n265), .A2(new_n267), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G107), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n273), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n291), .A2(new_n294), .A3(new_n280), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n263), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n285), .A2(new_n280), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(new_n273), .A3(new_n271), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n294), .A3(new_n280), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n262), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n296), .A2(KEYINPUT89), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n302), .A3(new_n299), .A4(new_n262), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n239), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT15), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n304), .B(new_n306), .Z(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n249), .A2(new_n259), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G221), .B1(new_n260), .B2(G902), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n310), .B(KEYINPUT74), .Z(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  INV_X1    g127(.A(G104), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(new_n314), .B2(G107), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n272), .A3(G104), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(G107), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(G101), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n319), .A2(new_n323), .A3(G101), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT0), .A2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT0), .A2(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n191), .A2(G146), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n218), .A2(G143), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n326), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n218), .A2(G143), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n191), .A2(G146), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT0), .A4(G128), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n319), .A2(G101), .ZN(new_n336));
  INV_X1    g150(.A(G101), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n315), .A2(new_n317), .A3(new_n337), .A4(new_n318), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(KEYINPUT4), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n325), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT10), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n272), .A2(G104), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n314), .A2(G107), .ZN(new_n343));
  OAI21_X1  g157(.A(G101), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n331), .A2(new_n332), .A3(new_n345), .A4(G128), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n348), .A2(G128), .B1(new_n331), .B2(new_n332), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n338), .B(new_n344), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n331), .A2(new_n332), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n281), .A2(new_n283), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n345), .B1(G143), .B2(new_n218), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n341), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n338), .A2(new_n344), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n341), .A2(new_n350), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT11), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n275), .B2(G137), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n275), .A2(G137), .ZN(new_n360));
  INV_X1    g174(.A(G137), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT11), .A3(G134), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G131), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n359), .A2(new_n362), .A3(new_n187), .A4(new_n360), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n340), .A2(new_n357), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n189), .A2(G227), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n368), .B2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n354), .A2(new_n346), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n350), .B1(new_n375), .B2(new_n356), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n366), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT12), .B1(new_n376), .B2(new_n366), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n373), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n367), .B1(new_n340), .B2(new_n357), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n372), .B1(new_n384), .B2(new_n368), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n313), .B(new_n239), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n372), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n368), .B1(new_n379), .B2(new_n380), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n368), .A2(new_n372), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n387), .A2(new_n388), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  OAI21_X1  g204(.A(G469), .B1(new_n390), .B2(G902), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n312), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n309), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n322), .A2(new_n324), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR3_X1   g211(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n399));
  INV_X1    g213(.A(G113), .ZN(new_n400));
  OAI22_X1  g214(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G116), .B(G119), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  OAI221_X1 g218(.A(new_n402), .B1(new_n399), .B2(new_n400), .C1(new_n397), .C2(new_n398), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n339), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n394), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  INV_X1    g223(.A(G119), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  OAI21_X1  g225(.A(G113), .B1(new_n411), .B2(KEYINPUT5), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(KEYINPUT5), .B2(new_n402), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n356), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n325), .A2(KEYINPUT78), .A3(new_n406), .A4(new_n339), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G122), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n408), .A2(new_n418), .A3(new_n415), .A4(new_n416), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT6), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n417), .A2(KEYINPUT79), .A3(KEYINPUT6), .A4(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n334), .A2(G125), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(G125), .B2(new_n375), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT80), .B(G224), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(G953), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n427), .B(new_n429), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n412), .B(KEYINPUT82), .Z(new_n433));
  NAND2_X1  g247(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n356), .B1(new_n437), .B2(new_n409), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n418), .B(KEYINPUT8), .ZN(new_n439));
  INV_X1    g253(.A(new_n356), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n414), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n438), .A2(KEYINPUT83), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n409), .B1(new_n433), .B2(new_n436), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n441), .B(new_n439), .C1(new_n443), .C2(new_n440), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT7), .B1(new_n428), .B2(G953), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n427), .B(new_n447), .Z(new_n448));
  NAND4_X1  g262(.A1(new_n442), .A2(new_n446), .A3(new_n421), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n239), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n432), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  INV_X1    g268(.A(new_n452), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n430), .B1(new_n423), .B2(new_n424), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(new_n450), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n456), .A2(new_n450), .A3(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT84), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n393), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n335), .A2(new_n366), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n361), .A2(G134), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n360), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G131), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n375), .A2(new_n365), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(new_n469), .A3(KEYINPUT30), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT64), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n334), .A2(new_n471), .B1(new_n364), .B2(new_n365), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n330), .A2(KEYINPUT64), .A3(new_n333), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n354), .A2(new_n346), .B1(G131), .B2(new_n467), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n472), .A2(new_n473), .B1(new_n365), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n406), .B(new_n470), .C1(new_n475), .C2(KEYINPUT30), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n474), .A2(new_n365), .B1(new_n335), .B2(new_n366), .ZN(new_n477));
  INV_X1    g291(.A(new_n406), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n476), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT31), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT28), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n477), .B2(new_n478), .ZN(new_n487));
  AND4_X1   g301(.A1(new_n486), .A2(new_n478), .A3(new_n465), .A4(new_n469), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n487), .A2(new_n488), .B1(new_n478), .B2(new_n475), .ZN(new_n489));
  INV_X1    g303(.A(new_n483), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT31), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n476), .A2(new_n492), .A3(new_n479), .A4(new_n483), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n485), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n494), .A2(KEYINPUT32), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT32), .B1(new_n494), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n464), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT67), .B1(new_n499), .B2(KEYINPUT32), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n476), .A2(new_n479), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n490), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n489), .A2(new_n483), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT29), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n477), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n406), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n506), .B1(new_n487), .B2(new_n488), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n483), .A2(KEYINPUT29), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n239), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G472), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n498), .A2(new_n500), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n279), .B2(new_n410), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n352), .A2(KEYINPUT68), .A3(G119), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT69), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n410), .B2(G128), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n276), .A2(KEYINPUT69), .A3(G119), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT24), .B(G110), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n279), .A2(new_n410), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT70), .B1(new_n410), .B2(G128), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n276), .A3(G119), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT23), .B1(new_n276), .B2(G119), .ZN(new_n528));
  AOI22_X1  g342(.A1(KEYINPUT23), .A2(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n519), .A2(new_n532), .A3(new_n520), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n205), .A3(new_n220), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n204), .A2(new_n205), .ZN(new_n536));
  OAI221_X1 g350(.A(new_n536), .B1(new_n530), .B2(new_n529), .C1(new_n520), .C2(new_n519), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(KEYINPUT73), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT22), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G137), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT73), .B1(new_n535), .B2(new_n537), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n537), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n239), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT25), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n261), .B1(G234), .B2(new_n239), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n546), .A2(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n538), .A3(new_n542), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n548), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT25), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n239), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n552), .A2(G902), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n511), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n463), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(G101), .ZN(G3));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n301), .A2(new_n565), .A3(new_n303), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT90), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n301), .A2(new_n568), .A3(new_n565), .A4(new_n303), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n300), .A2(KEYINPUT91), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n298), .A2(new_n572), .A3(new_n299), .A4(new_n262), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n571), .A2(KEYINPUT33), .A3(new_n296), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n305), .A2(G902), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT92), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n304), .A2(new_n305), .ZN(new_n578));
  INV_X1    g392(.A(new_n574), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n567), .B2(new_n569), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT92), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n575), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n249), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n459), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n586), .B(new_n259), .C1(new_n453), .C2(new_n457), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n386), .A2(new_n391), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n494), .A2(new_n239), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n494), .A2(new_n495), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n311), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n561), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  NOR2_X1   g412(.A1(new_n249), .A2(new_n307), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n587), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT35), .B(G107), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G9));
  NAND2_X1  g418(.A1(new_n592), .A2(new_n593), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n546), .B(KEYINPUT93), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n542), .A2(KEYINPUT36), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n606), .A2(KEYINPUT36), .A3(new_n542), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n559), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n605), .B1(new_n558), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n463), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT94), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT37), .B(G110), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G12));
  NAND3_X1  g430(.A1(new_n498), .A2(new_n500), .A3(new_n510), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n617), .A2(new_n392), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n452), .B1(new_n432), .B2(new_n451), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n459), .B1(new_n619), .B2(new_n460), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n558), .B2(new_n611), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT95), .B(G900), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n254), .B1(new_n258), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n249), .A2(new_n307), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n618), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  XNOR2_X1  g440(.A(new_n623), .B(KEYINPUT39), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n392), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n501), .A2(new_n490), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n506), .A2(new_n479), .A3(new_n490), .ZN(new_n633));
  OR3_X1    g447(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT96), .B1(new_n632), .B2(new_n633), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n634), .A2(new_n239), .A3(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n500), .B(new_n498), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n558), .A2(new_n611), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n586), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n631), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n458), .A2(new_n461), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT38), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n249), .A2(new_n308), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n458), .A2(new_n646), .A3(new_n461), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n643), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n641), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n191), .ZN(G45));
  INV_X1    g464(.A(new_n623), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n583), .A2(new_n249), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n621), .A2(new_n617), .A3(new_n392), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT97), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G146), .ZN(G48));
  INV_X1    g469(.A(new_n560), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n556), .B1(new_n555), .B2(new_n239), .ZN(new_n657));
  AOI211_X1 g471(.A(KEYINPUT25), .B(G902), .C1(new_n554), .C2(new_n548), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n656), .B1(new_n659), .B2(new_n552), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT98), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n313), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n368), .A2(new_n372), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT77), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n377), .B(new_n378), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n385), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n663), .B1(new_n670), .B2(new_n239), .ZN(new_n671));
  AOI211_X1 g485(.A(G902), .B(new_n662), .C1(new_n668), .C2(new_n669), .ZN(new_n672));
  INV_X1    g486(.A(new_n310), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n660), .A2(new_n617), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n588), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT41), .B(G113), .Z(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT99), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n676), .B(new_n678), .ZN(G15));
  NOR2_X1   g493(.A1(new_n675), .A2(new_n600), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n266), .ZN(G18));
  NAND3_X1  g495(.A1(new_n617), .A2(new_n309), .A3(new_n674), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n586), .B1(new_n453), .B2(new_n457), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n639), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n410), .ZN(G21));
  NAND2_X1  g500(.A1(new_n507), .A2(new_n490), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n485), .A2(new_n493), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n495), .B(KEYINPUT100), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT102), .B1(new_n591), .B2(G472), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n696));
  AOI211_X1 g510(.A(new_n696), .B(new_n637), .C1(new_n494), .C2(new_n239), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n660), .A2(new_n587), .A3(new_n674), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n644), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n264), .ZN(G24));
  NAND2_X1  g515(.A1(new_n683), .A2(new_n674), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n639), .A3(new_n652), .A4(new_n698), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  AOI211_X1 g519(.A(G469), .B(G902), .C1(new_n668), .C2(new_n669), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n388), .A2(new_n387), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n389), .A2(new_n384), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n313), .B1(new_n709), .B2(new_n239), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n310), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n586), .B(new_n711), .C1(new_n458), .C2(new_n461), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n713));
  OR3_X1    g527(.A1(new_n496), .A2(new_n497), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n713), .B1(new_n496), .B2(new_n497), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n510), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n660), .A3(new_n652), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n586), .B1(new_n458), .B2(new_n461), .ZN(new_n719));
  INV_X1    g533(.A(new_n711), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n718), .A2(new_n652), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n717), .A2(KEYINPUT42), .B1(new_n721), .B2(new_n562), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND3_X1  g537(.A1(new_n562), .A2(new_n624), .A3(new_n712), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT104), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G134), .ZN(G36));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n242), .A2(new_n247), .A3(new_n727), .A4(new_n248), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n242), .A2(new_n247), .A3(new_n248), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n583), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n583), .B(new_n731), .C1(new_n727), .C2(KEYINPUT43), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n605), .A3(new_n639), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT44), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n372), .B1(new_n666), .B2(new_n368), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n664), .A2(new_n383), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(G469), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(G469), .A2(G902), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n745), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n386), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n310), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n627), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n736), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n738), .A2(new_n719), .A3(new_n752), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT106), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n706), .B1(new_n746), .B2(new_n747), .ZN(new_n759));
  AOI211_X1 g573(.A(new_n758), .B(new_n673), .C1(new_n759), .C2(new_n749), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT47), .B1(new_n750), .B2(new_n310), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n652), .B(new_n719), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n660), .A2(new_n617), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n757), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n583), .A2(new_n249), .A3(new_n651), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n751), .A2(new_n758), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n310), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n719), .A4(new_n763), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n765), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G140), .ZN(G42));
  AND4_X1   g586(.A1(new_n660), .A2(new_n587), .A3(new_n674), .A4(new_n698), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n671), .A2(new_n672), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n310), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n511), .A2(new_n561), .A3(new_n775), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n773), .A2(new_n645), .B1(new_n776), .B2(new_n589), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n721), .A2(new_n562), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n617), .A2(new_n309), .A3(new_n674), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n776), .A2(new_n601), .B1(new_n780), .B2(new_n621), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(new_n778), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n652), .A2(new_n719), .A3(new_n698), .A4(new_n720), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n249), .A2(new_n308), .A3(new_n623), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n719), .A2(new_n617), .A3(new_n392), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n639), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n463), .B1(new_n562), .B2(new_n612), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n584), .A2(KEYINPUT109), .ZN(new_n789));
  INV_X1    g603(.A(new_n599), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n583), .A2(new_n791), .A3(new_n249), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n552), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n657), .A2(new_n658), .A3(new_n794), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n795), .A2(new_n594), .A3(new_n656), .A4(new_n259), .ZN(new_n796));
  INV_X1    g610(.A(new_n462), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n787), .A2(new_n724), .A3(new_n788), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n782), .A2(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n558), .A2(new_n611), .A3(new_n651), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n620), .A2(new_n644), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n638), .A3(new_n720), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n625), .A2(new_n653), .A3(new_n803), .A4(new_n704), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n639), .A2(new_n683), .A3(new_n624), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n592), .A2(new_n696), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n591), .A2(KEYINPUT102), .A3(G472), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n691), .A3(new_n693), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n558), .B2(new_n611), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n702), .A2(new_n766), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n806), .A2(new_n618), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n812), .A2(new_n813), .A3(new_n653), .A4(new_n803), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n805), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g629(.A(KEYINPUT110), .B(KEYINPUT53), .Z(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n800), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n788), .A2(new_n798), .A3(new_n724), .ZN(new_n819));
  OAI22_X1  g633(.A1(new_n699), .A2(new_n644), .B1(new_n675), .B2(new_n588), .ZN(new_n820));
  OAI22_X1  g634(.A1(new_n675), .A2(new_n600), .B1(new_n682), .B2(new_n684), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n822), .A3(new_n722), .A4(new_n787), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n805), .A2(new_n814), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT53), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT111), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n800), .A2(new_n815), .A3(KEYINPUT53), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n817), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT111), .A4(new_n829), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n253), .B1(new_n733), .B2(new_n734), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n642), .A2(new_n459), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n775), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT113), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n716), .A2(new_n660), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n834), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(KEYINPUT48), .B(new_n843), .C1(new_n840), .C2(new_n841), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n719), .A2(new_n674), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n558), .A2(new_n560), .A3(new_n254), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n848), .A2(new_n638), .A3(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n250), .B(G953), .C1(new_n850), .C2(new_n585), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n561), .A2(new_n809), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n835), .A2(new_n852), .A3(new_n703), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT114), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n835), .A2(new_n852), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT114), .A3(new_n703), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n857), .A4(new_n855), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n643), .A2(new_n647), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n674), .A2(new_n586), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT112), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n863), .A2(KEYINPUT112), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n856), .A2(new_n866), .A3(KEYINPUT50), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT50), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n835), .A2(new_n852), .A3(new_n867), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n865), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n760), .A2(new_n761), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n774), .A2(new_n312), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n836), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n583), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n848), .A2(new_n638), .A3(new_n849), .A4(new_n249), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n875), .A2(new_n856), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n842), .A2(new_n810), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n872), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT51), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n872), .A2(new_n878), .A3(new_n879), .A4(new_n882), .ZN(new_n883));
  AOI221_X4 g697(.A(new_n847), .B1(new_n860), .B2(new_n861), .C1(new_n881), .C2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n832), .A2(new_n833), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT116), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n250), .A2(new_n189), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n832), .A2(new_n884), .A3(new_n888), .A4(new_n833), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n561), .A2(new_n586), .A3(new_n312), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(KEYINPUT107), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT49), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n774), .A2(new_n894), .ZN(new_n895));
  OR4_X1    g709(.A1(new_n732), .A2(new_n892), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT108), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n638), .B1(new_n896), .B2(KEYINPUT108), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n774), .A2(new_n894), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n862), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n890), .A2(new_n900), .ZN(G75));
  AOI21_X1  g715(.A(new_n239), .B1(new_n828), .B2(new_n830), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(G210), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n425), .A2(new_n431), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n456), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n250), .A2(G953), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT117), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(G51));
  NAND2_X1  g727(.A1(new_n828), .A2(new_n830), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT118), .B1(new_n914), .B2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n831), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n828), .A2(new_n830), .A3(KEYINPUT118), .A4(new_n829), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n745), .B(KEYINPUT57), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n670), .ZN(new_n920));
  INV_X1    g734(.A(new_n744), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n902), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n912), .B1(new_n920), .B2(new_n922), .ZN(G54));
  INV_X1    g737(.A(new_n237), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n924), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT119), .B1(new_n925), .B2(new_n924), .ZN(new_n927));
  OAI221_X1 g741(.A(new_n911), .B1(new_n924), .B2(new_n925), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(G60));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n916), .A2(new_n580), .A3(new_n917), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n931), .B1(new_n832), .B2(new_n833), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n933), .B(new_n911), .C1(new_n934), .C2(new_n580), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n828), .B2(new_n830), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n609), .A2(new_n610), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n911), .B1(new_n939), .B2(new_n555), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n946));
  OAI221_X1 g760(.A(new_n911), .B1(KEYINPUT121), .B2(KEYINPUT61), .C1(new_n939), .C2(new_n555), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n942), .A2(new_n945), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n941), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT61), .B1(new_n949), .B2(new_n943), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(G66));
  NAND3_X1  g765(.A1(new_n822), .A2(new_n788), .A3(new_n798), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n189), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n256), .B2(new_n428), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n423), .B(new_n424), .C1(G898), .C2(new_n189), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  OAI21_X1  g771(.A(new_n470), .B1(new_n475), .B2(KEYINPUT30), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n229), .B(KEYINPUT122), .Z(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n625), .A2(new_n653), .A3(new_n704), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(KEYINPUT62), .C1(new_n648), .C2(new_n641), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n812), .A2(new_n653), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n649), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n836), .A2(new_n629), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(new_n562), .A3(new_n793), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT123), .Z(new_n969));
  NAND4_X1  g783(.A1(new_n966), .A2(new_n755), .A3(new_n771), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n960), .B1(new_n970), .B2(new_n189), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n752), .A2(new_n844), .A3(new_n802), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n722), .A2(new_n961), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n975), .A2(new_n771), .A3(new_n755), .A4(new_n724), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n189), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(G900), .B2(new_n189), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(KEYINPUT125), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n977), .B(new_n980), .C1(G900), .C2(new_n189), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n960), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n973), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n973), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n976), .B2(new_n952), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n502), .B(KEYINPUT127), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n912), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n970), .A2(new_n952), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n988), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT126), .B1(new_n993), .B2(new_n632), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  INV_X1    g809(.A(new_n632), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n995), .B(new_n996), .C1(new_n992), .C2(new_n988), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n991), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n818), .A2(new_n825), .ZN(new_n999));
  AND4_X1   g813(.A1(new_n502), .A2(new_n999), .A3(new_n996), .A4(new_n988), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n998), .A2(new_n1000), .ZN(G57));
endmodule


