//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(KEYINPUT0), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n187), .A2(new_n188), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n190), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT64), .B1(new_n193), .B2(G146), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n192), .B(new_n189), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(new_n191), .B2(G143), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n193), .A2(KEYINPUT64), .A3(G146), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n204), .A2(new_n205), .B1(G143), .B2(new_n191), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(new_n189), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n198), .B1(new_n202), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT80), .B(new_n211), .C1(new_n213), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G107), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G104), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n212), .A2(KEYINPUT3), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n216), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n217), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G101), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n223), .B(new_n222), .C1(new_n229), .C2(new_n218), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n230), .B2(new_n216), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n228), .B(KEYINPUT4), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n226), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n225), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT81), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT81), .ZN(new_n238));
  NOR4_X1   g052(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT4), .A4(new_n232), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n209), .B(new_n233), .C1(new_n237), .C2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n232), .B1(new_n234), .B2(new_n218), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n192), .B(new_n244), .C1(new_n199), .C2(new_n200), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n188), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n206), .B2(new_n246), .ZN(new_n247));
  AND4_X1   g061(.A1(KEYINPUT82), .A2(new_n228), .A3(new_n243), .A4(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n225), .B2(new_n227), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT82), .B1(new_n249), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n241), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT66), .B(new_n252), .C1(new_n253), .C2(G137), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G134), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT66), .B1(new_n257), .B2(new_n252), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n252), .A2(new_n253), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n256), .A2(G134), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n259), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(G137), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n269), .B2(new_n260), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT66), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n254), .ZN(new_n274));
  INV_X1    g088(.A(G131), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(G143), .B(G146), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n246), .A2(new_n279), .A3(KEYINPUT68), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G128), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n195), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n245), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n249), .A2(KEYINPUT10), .A3(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n240), .A2(new_n251), .A3(new_n278), .A4(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n249), .A2(new_n285), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n228), .A2(new_n243), .A3(new_n247), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n249), .A2(KEYINPUT82), .A3(new_n247), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT12), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n248), .A2(new_n250), .B1(new_n285), .B2(new_n249), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n277), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G140), .ZN(new_n299));
  INV_X1    g113(.A(G953), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n300), .A2(G227), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n299), .B(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n240), .A2(new_n251), .A3(new_n286), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n277), .A2(KEYINPUT85), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n240), .A2(new_n251), .A3(new_n306), .A4(new_n286), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n302), .ZN(new_n310));
  INV_X1    g124(.A(G469), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n304), .A2(new_n310), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n303), .B1(new_n298), .B2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n287), .A2(new_n294), .A3(new_n297), .A4(KEYINPUT84), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n308), .A2(new_n309), .A3(new_n303), .ZN(new_n320));
  AOI21_X1  g134(.A(G902), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI22_X1  g135(.A1(new_n314), .A2(new_n315), .B1(new_n321), .B2(new_n311), .ZN(new_n322));
  INV_X1    g136(.A(G221), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT9), .B(G234), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n323), .B1(new_n325), .B2(new_n312), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G113), .B(G122), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(new_n210), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT77), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n333), .A2(KEYINPUT77), .A3(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT16), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT16), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G146), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n191), .A3(new_n339), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(KEYINPUT78), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n347));
  INV_X1    g161(.A(G237), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n300), .A3(G214), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n193), .ZN(new_n350));
  NOR2_X1   g164(.A1(G237), .A2(G953), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(G143), .A3(G214), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n347), .B1(new_n353), .B2(G131), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(G131), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n275), .A3(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n357), .B2(new_n347), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n346), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT18), .A2(G131), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n353), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n335), .A2(new_n336), .A3(G146), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n332), .A2(new_n334), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n191), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n330), .B1(new_n360), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n343), .B2(new_n345), .ZN(new_n369));
  INV_X1    g183(.A(new_n330), .ZN(new_n370));
  INV_X1    g184(.A(new_n367), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n312), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT92), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT92), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(new_n312), .C1(new_n368), .C2(new_n372), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(G475), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n340), .A2(G146), .B1(new_n355), .B2(new_n356), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT19), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n335), .B2(new_n336), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n364), .A2(KEYINPUT19), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n191), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n379), .A2(new_n383), .B1(new_n362), .B2(new_n366), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT91), .B1(new_n384), .B2(new_n330), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n341), .A2(new_n383), .A3(new_n357), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n367), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n387), .A2(new_n388), .A3(new_n370), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n378), .B1(new_n390), .B2(new_n372), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT20), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n393), .B(new_n378), .C1(new_n390), .C2(new_n372), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n377), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT69), .ZN(new_n398));
  INV_X1    g212(.A(G116), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT69), .A2(G116), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(G122), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n399), .A2(G122), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n402), .B2(new_n404), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(G107), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT93), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n217), .B1(new_n410), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n397), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G107), .B1(new_n406), .B2(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n217), .A3(new_n405), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT94), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n193), .A2(G128), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n188), .A2(G143), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n418), .A2(new_n253), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(KEYINPUT95), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT95), .B1(new_n416), .B2(new_n420), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n417), .B1(new_n420), .B2(new_n416), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n419), .B1(new_n424), .B2(G134), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n415), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n400), .A2(KEYINPUT14), .A3(G122), .A4(new_n401), .ZN(new_n427));
  OAI211_X1 g241(.A(G107), .B(new_n427), .C1(new_n409), .C2(KEYINPUT14), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n418), .A2(new_n253), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n414), .B(new_n428), .C1(new_n419), .C2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G217), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n324), .A2(new_n431), .A3(G953), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n426), .B2(new_n430), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n312), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT15), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(G478), .ZN(new_n437));
  INV_X1    g251(.A(G478), .ZN(new_n438));
  OAI221_X1 g252(.A(new_n312), .B1(KEYINPUT15), .B2(new_n438), .C1(new_n433), .C2(new_n434), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n300), .A2(G952), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(G234), .B2(G237), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n312), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(G898), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n396), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT90), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n209), .A2(G125), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n285), .A2(new_n333), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n300), .A2(G224), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT88), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n452), .B(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n400), .A2(G119), .A3(new_n401), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n399), .A2(G119), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n458), .A2(KEYINPUT70), .A3(new_n460), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(KEYINPUT5), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G113), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT5), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT2), .B(G113), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n458), .A3(new_n460), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n472), .A3(new_n249), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n237), .A2(new_n239), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n471), .B1(new_n463), .B2(new_n464), .ZN(new_n476));
  INV_X1    g290(.A(new_n472), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT71), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n464), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT70), .B1(new_n458), .B2(new_n460), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n470), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n472), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n233), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT6), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n475), .B2(new_n484), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n474), .A2(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(KEYINPUT6), .A3(new_n488), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n457), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n455), .A2(KEYINPUT7), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n452), .B(new_n493), .Z(new_n494));
  XOR2_X1   g308(.A(new_n474), .B(KEYINPUT8), .Z(new_n495));
  OAI21_X1  g309(.A(new_n468), .B1(new_n461), .B2(new_n467), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n472), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n249), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n469), .A2(new_n472), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n249), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n500), .A2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n485), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n312), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n449), .B1(new_n492), .B2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n485), .A2(KEYINPUT6), .B1(new_n487), .B2(new_n488), .ZN(new_n509));
  INV_X1    g323(.A(new_n491), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n456), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n452), .B(new_n493), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n500), .A2(new_n501), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n502), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n514), .B2(new_n485), .ZN(new_n515));
  INV_X1    g329(.A(new_n449), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n446), .A2(new_n447), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n351), .A2(G210), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT27), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(G101), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n202), .A2(new_n208), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n270), .A2(new_n274), .A3(new_n275), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n275), .B1(new_n270), .B2(new_n274), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(new_n197), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n257), .B1(new_n269), .B2(G134), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G131), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n285), .A2(new_n276), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n532), .A2(KEYINPUT73), .B1(new_n478), .B2(new_n483), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n276), .A2(new_n530), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n285), .A2(new_n534), .B1(new_n277), .B2(new_n209), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT28), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n478), .A2(new_n483), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n532), .A2(new_n478), .A3(new_n483), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n524), .B1(new_n538), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g360(.A(new_n541), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n528), .A2(new_n548), .A3(new_n531), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n528), .B2(new_n531), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n523), .A3(new_n542), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT31), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n551), .A2(KEYINPUT31), .A3(new_n523), .A4(new_n542), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n557), .B(new_n524), .C1(new_n538), .C2(new_n544), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n546), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G472), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n312), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n559), .A2(KEYINPUT32), .A3(new_n560), .A4(new_n312), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT29), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n551), .A2(new_n542), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n524), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n538), .A2(new_n544), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n567), .C1(new_n568), .C2(new_n524), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n542), .A2(new_n543), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n538), .B1(KEYINPUT28), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n524), .A2(new_n565), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n563), .A2(new_n564), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n431), .B1(G234), .B2(new_n312), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G119), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G128), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(KEYINPUT75), .A3(G128), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n582), .B(new_n583), .C1(new_n579), .C2(G128), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT24), .B(G110), .ZN(new_n585));
  OR2_X1    g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n579), .A2(G128), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n580), .B(new_n587), .C1(new_n588), .C2(KEYINPUT23), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT76), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n343), .A2(new_n345), .A3(new_n586), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n589), .A2(G110), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n584), .A2(new_n585), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n341), .B(new_n365), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT22), .B(G137), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n300), .A2(G221), .A3(G234), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n597), .B(new_n598), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n596), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n312), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT25), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(KEYINPUT25), .A3(new_n312), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n578), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n577), .A2(G902), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n328), .A2(new_n519), .A3(new_n576), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  AND3_X1   g426(.A1(new_n559), .A2(new_n560), .A3(new_n312), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n560), .B1(new_n559), .B2(new_n312), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n448), .B1(new_n492), .B2(new_n507), .ZN(new_n616));
  INV_X1    g430(.A(new_n445), .ZN(new_n617));
  INV_X1    g431(.A(new_n448), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n511), .A2(new_n515), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n616), .A2(new_n447), .A3(new_n617), .A4(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n433), .B2(new_n434), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n426), .A2(new_n430), .ZN(new_n626));
  INV_X1    g440(.A(new_n432), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n622), .C1(new_n623), .C2(new_n621), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n438), .A2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(KEYINPUT97), .A3(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n438), .B(G902), .C1(new_n625), .C2(new_n629), .ZN(new_n633));
  AOI21_X1  g447(.A(KEYINPUT97), .B1(new_n435), .B2(new_n438), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n396), .B(new_n632), .C1(new_n633), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n620), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n615), .A2(new_n328), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND2_X1   g454(.A1(new_n440), .A2(new_n377), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n392), .A2(KEYINPUT98), .A3(new_n394), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n394), .A2(KEYINPUT98), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n620), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n328), .A2(new_n615), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(new_n599), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n596), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n607), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n605), .A2(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n613), .A2(new_n655), .A3(new_n614), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n328), .A2(new_n656), .A3(new_n519), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT99), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n657), .B(new_n659), .ZN(G12));
  INV_X1    g474(.A(new_n655), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n576), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n616), .A2(new_n447), .A3(new_n619), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n322), .A2(new_n327), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n442), .B(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n443), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n645), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G128), .ZN(G30));
  XOR2_X1   g487(.A(new_n670), .B(KEYINPUT39), .Z(new_n674));
  NAND2_X1  g488(.A1(new_n328), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  INV_X1    g490(.A(new_n518), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT38), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT38), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n518), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n447), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n396), .A2(new_n440), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n661), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT40), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n328), .A2(new_n686), .A3(new_n674), .ZN(new_n687));
  INV_X1    g501(.A(new_n566), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n524), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n312), .B1(new_n570), .B2(new_n523), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n563), .A2(new_n564), .A3(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n676), .A2(new_n685), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  NAND2_X1  g508(.A1(new_n630), .A2(new_n631), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n634), .ZN(new_n696));
  INV_X1    g510(.A(new_n670), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n396), .A3(new_n632), .A4(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n666), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  AND2_X1   g515(.A1(new_n576), .A2(new_n610), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n304), .A2(new_n312), .A3(new_n310), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n304), .A2(new_n310), .A3(KEYINPUT101), .A4(new_n312), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(G469), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n707), .B(new_n327), .C1(new_n315), .C2(new_n314), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n313), .A2(KEYINPUT86), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n706), .A2(G469), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n711), .A2(new_n712), .B1(new_n713), .B2(new_n705), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n327), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n702), .A2(new_n637), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n702), .A2(new_n646), .A3(new_n710), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  OAI21_X1  g534(.A(KEYINPUT103), .B1(new_n708), .B2(new_n663), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n714), .A2(new_n722), .A3(new_n327), .A4(new_n664), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n576), .A2(new_n446), .A3(new_n661), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  INV_X1    g541(.A(new_n570), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT28), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n524), .B1(new_n730), .B2(new_n538), .ZN(new_n731));
  AOI211_X1 g545(.A(G472), .B(G902), .C1(new_n731), .C2(new_n556), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n609), .A2(new_n614), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n620), .A2(new_n683), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n715), .A2(new_n710), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR4_X1   g550(.A1(new_n698), .A2(new_n655), .A3(new_n614), .A4(new_n732), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n724), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  NAND3_X1  g553(.A1(new_n613), .A2(KEYINPUT106), .A3(KEYINPUT32), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n561), .A2(new_n562), .B1(G472), .B2(new_n574), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n564), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n610), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n326), .A2(new_n682), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n508), .A2(new_n517), .A3(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n320), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n308), .A2(KEYINPUT105), .A3(new_n309), .A4(new_n303), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n319), .A2(G469), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(G469), .A2(G902), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT104), .Z(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n711), .A2(new_n712), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n747), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n699), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT42), .B1(new_n745), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n702), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  OAI21_X1  g577(.A(KEYINPUT107), .B1(new_n645), .B2(new_n670), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n641), .A2(new_n644), .A3(new_n765), .A4(new_n697), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n702), .A2(new_n767), .A3(new_n757), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n696), .A2(new_n632), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n377), .A2(new_n395), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n396), .B(KEYINPUT110), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n696), .A2(KEYINPUT43), .A3(new_n632), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT111), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n396), .B(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT111), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT43), .A4(new_n773), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n775), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n661), .B1(new_n613), .B2(new_n614), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n770), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n508), .A2(new_n447), .A3(new_n517), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n784), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n778), .A2(new_n782), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT44), .B(new_n789), .C1(new_n790), .C2(new_n775), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n319), .A2(KEYINPUT45), .A3(new_n749), .A4(new_n750), .ZN(new_n792));
  INV_X1    g606(.A(new_n320), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n318), .B2(new_n317), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n792), .B(G469), .C1(KEYINPUT45), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n754), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n796), .A2(new_n797), .B1(new_n711), .B2(new_n712), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n326), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(KEYINPUT108), .A3(new_n674), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT108), .B1(new_n800), .B2(new_n674), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n788), .B(new_n791), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XNOR2_X1  g619(.A(new_n800), .B(KEYINPUT47), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n699), .A2(new_n609), .A3(new_n787), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(new_n576), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  NAND4_X1  g625(.A1(new_n610), .A2(new_n780), .A3(new_n773), .A4(new_n746), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT112), .ZN(new_n813));
  INV_X1    g627(.A(new_n714), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n681), .B1(KEYINPUT49), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n563), .A2(new_n564), .A3(new_n691), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n814), .A2(KEYINPUT49), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n733), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n783), .A2(new_n667), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n724), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n708), .A2(new_n786), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n610), .A2(new_n822), .A3(new_n442), .A4(new_n816), .ZN(new_n823));
  INV_X1    g637(.A(new_n636), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n441), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n783), .A2(new_n667), .ZN(new_n826));
  INV_X1    g640(.A(new_n745), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n822), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT48), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n821), .B(new_n825), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n681), .A2(new_n447), .A3(new_n708), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n733), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n820), .A2(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n838), .A2(new_n839), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n655), .A2(new_n614), .A3(new_n732), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n826), .A2(new_n841), .A3(new_n822), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n820), .A2(new_n787), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n814), .A2(new_n327), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n806), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n773), .A2(new_n396), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n823), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n840), .A2(new_n844), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n832), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n842), .A2(new_n843), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n783), .A2(new_n667), .A3(new_n708), .A4(new_n786), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n854), .B2(new_n841), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n849), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n834), .A2(new_n837), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n820), .A2(new_n835), .A3(new_n836), .A4(new_n833), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(KEYINPUT117), .B2(KEYINPUT50), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT119), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n840), .A2(new_n844), .A3(new_n861), .A4(new_n849), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n847), .A2(KEYINPUT51), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n852), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n663), .A2(new_n683), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n751), .B(new_n754), .C1(new_n314), .C2(new_n315), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n605), .A2(new_n654), .A3(new_n326), .A4(new_n670), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT114), .B1(new_n870), .B2(new_n816), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n606), .A2(new_n327), .A3(new_n653), .A4(new_n697), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n872), .B1(new_n755), .B2(new_n756), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n692), .A4(new_n867), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n662), .B(new_n665), .C1(new_n671), .C2(new_n699), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(new_n738), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n877), .A3(new_n738), .A4(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n437), .A2(new_n439), .A3(new_n697), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(new_n377), .A3(new_n643), .A4(new_n642), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n786), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n885), .A2(new_n322), .A3(new_n327), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n662), .A2(new_n886), .B1(new_n737), .B2(new_n757), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n759), .A2(new_n887), .A3(new_n761), .A4(new_n768), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n726), .A2(new_n716), .A3(new_n719), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n636), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n774), .A2(new_n440), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n636), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(new_n890), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n677), .A2(new_n682), .A3(new_n445), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n894), .A2(new_n328), .A3(new_n615), .A4(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n611), .A3(new_n657), .A4(new_n735), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n888), .A2(new_n889), .A3(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n882), .A2(new_n898), .A3(KEYINPUT53), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n882), .B2(new_n898), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n882), .A2(new_n898), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n882), .A2(new_n898), .A3(KEYINPUT53), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT54), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n866), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n901), .B1(new_n899), .B2(new_n900), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(KEYINPUT54), .A3(new_n906), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT115), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n865), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n818), .B1(new_n912), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n300), .A2(G952), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n509), .A2(new_n510), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n456), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  OAI211_X1 g732(.A(G210), .B(G902), .C1(new_n899), .C2(new_n900), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT120), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n924), .A3(new_n920), .A4(new_n918), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n915), .B(new_n921), .C1(new_n923), .C2(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n753), .B(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n909), .A2(new_n910), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(new_n304), .A3(new_n310), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n905), .A2(new_n906), .ZN(new_n931));
  INV_X1    g745(.A(new_n795), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(G902), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n915), .B1(new_n930), .B2(new_n933), .ZN(G54));
  NAND4_X1  g748(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n390), .A2(new_n372), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n915), .ZN(G60));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT59), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n909), .A2(new_n910), .A3(new_n630), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n915), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n908), .A2(new_n911), .A3(new_n942), .ZN(new_n946));
  INV_X1    g760(.A(new_n630), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(G217), .A2(G902), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT60), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n652), .B(new_n951), .C1(new_n899), .C2(new_n900), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n905), .B2(new_n906), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n952), .B(new_n944), .C1(new_n953), .C2(new_n600), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(KEYINPUT61), .ZN(new_n956));
  AOI21_X1  g770(.A(KEYINPUT61), .B1(new_n954), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  INV_X1    g772(.A(G224), .ZN(new_n959));
  OAI21_X1  g773(.A(G953), .B1(new_n444), .B2(new_n959), .ZN(new_n960));
  OR3_X1    g774(.A1(new_n889), .A2(new_n897), .A3(KEYINPUT123), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT123), .B1(new_n889), .B2(new_n897), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n916), .B1(G898), .B2(new_n300), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  NAND2_X1  g780(.A1(G227), .A2(G900), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(G953), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n549), .A2(new_n550), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n381), .A2(new_n382), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n969), .B(new_n970), .Z(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  INV_X1    g786(.A(new_n693), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n877), .A2(new_n738), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n693), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n702), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n979), .A2(new_n675), .A3(new_n786), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n894), .B(KEYINPUT124), .ZN(new_n981));
  AOI22_X1  g795(.A1(new_n806), .A2(new_n809), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n982), .A3(new_n804), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n971), .B1(new_n984), .B2(G953), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n669), .A2(G953), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT125), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n791), .A2(new_n787), .A3(new_n785), .ZN(new_n990));
  INV_X1    g804(.A(new_n803), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n801), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n992), .B2(new_n974), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n804), .A2(KEYINPUT126), .A3(new_n976), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n827), .B(new_n867), .C1(new_n802), .C2(new_n803), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n762), .A2(new_n768), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(new_n810), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n988), .B1(new_n1000), .B2(new_n300), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n968), .B(new_n985), .C1(new_n1001), .C2(new_n971), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n998), .B1(new_n993), .B2(new_n994), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n987), .B1(new_n1003), .B2(G953), .ZN(new_n1004));
  OAI211_X1 g818(.A(G953), .B(new_n967), .C1(new_n1004), .C2(new_n971), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1002), .A2(new_n1005), .ZN(G72));
  INV_X1    g820(.A(new_n689), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n963), .A2(new_n978), .A3(new_n804), .A4(new_n982), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  AOI21_X1  g824(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1010), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n567), .B2(new_n552), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n915), .B1(new_n931), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1014), .B1(new_n1003), .B2(new_n963), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n688), .A2(new_n524), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1013), .A2(new_n1019), .ZN(G57));
endmodule


