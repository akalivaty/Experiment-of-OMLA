

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787;

  NOR2_X1 U375 ( .A1(n785), .A2(n787), .ZN(n463) );
  NOR2_X2 U376 ( .A1(n687), .A2(n689), .ZN(n731) );
  XNOR2_X1 U377 ( .A(n477), .B(n476), .ZN(n520) );
  XNOR2_X1 U378 ( .A(n465), .B(G107), .ZN(n500) );
  AND2_X1 U379 ( .A1(n772), .A2(n529), .ZN(n354) );
  OR2_X2 U380 ( .A1(n655), .A2(KEYINPUT44), .ZN(n656) );
  XNOR2_X2 U381 ( .A(n386), .B(n385), .ZN(n622) );
  NOR2_X2 U382 ( .A1(n626), .A2(n425), .ZN(n386) );
  XNOR2_X2 U383 ( .A(n381), .B(n494), .ZN(n501) );
  NOR2_X2 U384 ( .A1(n593), .A2(n592), .ZN(n595) );
  XNOR2_X2 U385 ( .A(n491), .B(n490), .ZN(n593) );
  XOR2_X2 U386 ( .A(KEYINPUT38), .B(n489), .Z(n726) );
  NAND2_X1 U387 ( .A1(n389), .A2(n388), .ZN(n772) );
  NAND2_X1 U388 ( .A1(n361), .A2(n355), .ZN(n417) );
  NOR2_X1 U389 ( .A1(n593), .A2(n488), .ZN(n439) );
  NOR2_X1 U390 ( .A1(n642), .A2(n570), .ZN(n571) );
  AND2_X1 U391 ( .A1(n406), .A2(n405), .ZN(n404) );
  XNOR2_X1 U392 ( .A(n545), .B(n544), .ZN(n624) );
  XNOR2_X1 U393 ( .A(KEYINPUT23), .B(KEYINPUT95), .ZN(n537) );
  XOR2_X1 U394 ( .A(G137), .B(G134), .Z(n495) );
  AND2_X2 U395 ( .A1(n469), .A2(n365), .ZN(n387) );
  XNOR2_X1 U396 ( .A(n575), .B(n574), .ZN(n612) );
  NOR2_X1 U397 ( .A1(n622), .A2(n710), .ZN(n617) );
  XNOR2_X2 U398 ( .A(G104), .B(G110), .ZN(n465) );
  NOR2_X1 U399 ( .A1(G237), .A2(G953), .ZN(n515) );
  XNOR2_X1 U400 ( .A(n467), .B(G140), .ZN(n548) );
  INV_X1 U401 ( .A(G131), .ZN(n467) );
  XNOR2_X1 U402 ( .A(n693), .B(KEYINPUT87), .ZN(n462) );
  XNOR2_X1 U403 ( .A(n463), .B(KEYINPUT46), .ZN(n443) );
  XNOR2_X1 U404 ( .A(n565), .B(n433), .ZN(n569) );
  XNOR2_X1 U405 ( .A(n566), .B(G478), .ZN(n433) );
  XNOR2_X1 U406 ( .A(n556), .B(n428), .ZN(n586) );
  XNOR2_X1 U407 ( .A(n429), .B(G475), .ZN(n428) );
  INV_X1 U408 ( .A(KEYINPUT13), .ZN(n429) );
  XNOR2_X1 U409 ( .A(n536), .B(KEYINPUT10), .ZN(n547) );
  NAND2_X1 U410 ( .A1(n399), .A2(n398), .ZN(n397) );
  OR2_X1 U411 ( .A1(n725), .A2(KEYINPUT30), .ZN(n398) );
  NAND2_X1 U412 ( .A1(n400), .A2(n391), .ZN(n390) );
  NAND2_X1 U413 ( .A1(G472), .A2(G902), .ZN(n405) );
  XOR2_X1 U414 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n516) );
  XNOR2_X1 U415 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n538) );
  XOR2_X1 U416 ( .A(G146), .B(G125), .Z(n536) );
  AND2_X1 U417 ( .A1(n462), .A2(n598), .ZN(n453) );
  AND2_X1 U418 ( .A1(n464), .A2(n462), .ZN(n444) );
  AND2_X1 U419 ( .A1(n443), .A2(n607), .ZN(n382) );
  OR2_X1 U420 ( .A1(G237), .A2(G902), .ZN(n513) );
  INV_X1 U421 ( .A(n623), .ZN(n642) );
  NAND2_X1 U422 ( .A1(n588), .A2(n725), .ZN(n575) );
  INV_X1 U423 ( .A(KEYINPUT22), .ZN(n385) );
  NAND2_X1 U424 ( .A1(n615), .A2(n426), .ZN(n425) );
  XNOR2_X1 U425 ( .A(n450), .B(n535), .ZN(n449) );
  XNOR2_X1 U426 ( .A(G119), .B(G137), .ZN(n535) );
  XNOR2_X1 U427 ( .A(n537), .B(n451), .ZN(n450) );
  INV_X1 U428 ( .A(KEYINPUT94), .ZN(n451) );
  XNOR2_X1 U429 ( .A(n427), .B(n770), .ZN(n668) );
  XNOR2_X1 U430 ( .A(n555), .B(n359), .ZN(n427) );
  XNOR2_X1 U431 ( .A(n357), .B(n554), .ZN(n555) );
  INV_X1 U432 ( .A(KEYINPUT73), .ZN(n490) );
  AND2_X1 U433 ( .A1(n581), .A2(n580), .ZN(n431) );
  NOR2_X1 U434 ( .A1(n356), .A2(n621), .ZN(n484) );
  NOR2_X1 U435 ( .A1(n356), .A2(n481), .ZN(n480) );
  NAND2_X1 U436 ( .A1(n379), .A2(KEYINPUT106), .ZN(n481) );
  INV_X2 U437 ( .A(G953), .ZN(n773) );
  XNOR2_X1 U438 ( .A(G116), .B(G122), .ZN(n563) );
  XNOR2_X1 U439 ( .A(n562), .B(n435), .ZN(n564) );
  NOR2_X1 U440 ( .A1(G952), .A2(n773), .ZN(n758) );
  NAND2_X1 U441 ( .A1(n708), .A2(n773), .ZN(n384) );
  AND2_X1 U442 ( .A1(n725), .A2(KEYINPUT30), .ZN(n400) );
  NAND2_X1 U443 ( .A1(n521), .A2(n403), .ZN(n402) );
  INV_X1 U444 ( .A(G902), .ZN(n403) );
  AND2_X1 U445 ( .A1(n636), .A2(n782), .ZN(n637) );
  AND2_X1 U446 ( .A1(n363), .A2(n408), .ZN(n407) );
  OR2_X1 U447 ( .A1(n582), .A2(n414), .ZN(n408) );
  XNOR2_X1 U448 ( .A(KEYINPUT3), .B(G116), .ZN(n499) );
  XNOR2_X1 U449 ( .A(G113), .B(G143), .ZN(n551) );
  XOR2_X1 U450 ( .A(G122), .B(G104), .Z(n552) );
  XOR2_X1 U451 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n550) );
  XNOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n549) );
  XNOR2_X1 U453 ( .A(n362), .B(n548), .ZN(n466) );
  NAND2_X1 U454 ( .A1(G234), .A2(G237), .ZN(n522) );
  XOR2_X1 U455 ( .A(KEYINPUT93), .B(KEYINPUT14), .Z(n523) );
  NAND2_X1 U456 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U457 ( .A1(n404), .A2(n401), .ZN(n623) );
  XOR2_X1 U458 ( .A(n642), .B(KEYINPUT6), .Z(n628) );
  XNOR2_X1 U459 ( .A(n514), .B(n460), .ZN(n666) );
  XNOR2_X1 U460 ( .A(n519), .B(n520), .ZN(n460) );
  XNOR2_X1 U461 ( .A(G119), .B(G113), .ZN(n476) );
  XNOR2_X1 U462 ( .A(n499), .B(n478), .ZN(n477) );
  INV_X1 U463 ( .A(G101), .ZN(n478) );
  XNOR2_X1 U464 ( .A(KEYINPUT68), .B(G122), .ZN(n475) );
  XNOR2_X1 U465 ( .A(n561), .B(n436), .ZN(n435) );
  INV_X1 U466 ( .A(KEYINPUT7), .ZN(n436) );
  XNOR2_X1 U467 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n502) );
  XOR2_X1 U468 ( .A(KEYINPUT92), .B(KEYINPUT76), .Z(n503) );
  NAND2_X1 U469 ( .A1(n441), .A2(n382), .ZN(n389) );
  NAND2_X1 U470 ( .A1(n442), .A2(n364), .ZN(n388) );
  NOR2_X1 U471 ( .A1(KEYINPUT2), .A2(n373), .ZN(n699) );
  AND2_X1 U472 ( .A1(n726), .A2(n376), .ZN(n589) );
  XNOR2_X1 U473 ( .A(n599), .B(n459), .ZN(n458) );
  INV_X1 U474 ( .A(KEYINPUT110), .ZN(n459) );
  INV_X1 U475 ( .A(n575), .ZN(n457) );
  XNOR2_X1 U476 ( .A(n635), .B(KEYINPUT35), .ZN(n640) );
  NAND2_X1 U477 ( .A1(n567), .A2(n587), .ZN(n596) );
  XNOR2_X1 U478 ( .A(n520), .B(n472), .ZN(n765) );
  XNOR2_X1 U479 ( .A(n500), .B(n473), .ZN(n472) );
  XNOR2_X1 U480 ( .A(n475), .B(n474), .ZN(n473) );
  INV_X1 U481 ( .A(KEYINPUT16), .ZN(n474) );
  XNOR2_X1 U482 ( .A(n452), .B(n448), .ZN(n468) );
  XNOR2_X1 U483 ( .A(n540), .B(n534), .ZN(n452) );
  XNOR2_X1 U484 ( .A(n547), .B(n449), .ZN(n448) );
  XOR2_X1 U485 ( .A(n668), .B(KEYINPUT59), .Z(n669) );
  AND2_X1 U486 ( .A1(n454), .A2(n621), .ZN(n693) );
  XNOR2_X1 U487 ( .A(n456), .B(n455), .ZN(n454) );
  INV_X1 U488 ( .A(KEYINPUT36), .ZN(n455) );
  NAND2_X1 U489 ( .A1(n458), .A2(n457), .ZN(n456) );
  XNOR2_X1 U490 ( .A(n643), .B(KEYINPUT31), .ZN(n690) );
  INV_X1 U491 ( .A(KEYINPUT108), .ZN(n438) );
  BUF_X1 U492 ( .A(n612), .Z(n383) );
  AND2_X1 U493 ( .A1(n485), .A2(n367), .ZN(n483) );
  NAND2_X1 U494 ( .A1(n482), .A2(n480), .ZN(n479) );
  XNOR2_X1 U495 ( .A(n753), .B(n432), .ZN(n755) );
  XNOR2_X1 U496 ( .A(n754), .B(KEYINPUT122), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n749), .B(n434), .ZN(n752) );
  OR2_X1 U498 ( .A1(n706), .A2(n384), .ZN(n742) );
  AND2_X1 U499 ( .A1(n424), .A2(n664), .ZN(n355) );
  INV_X1 U500 ( .A(n709), .ZN(n426) );
  OR2_X1 U501 ( .A1(n719), .A2(n625), .ZN(n356) );
  XOR2_X1 U502 ( .A(n552), .B(n551), .Z(n357) );
  AND2_X1 U503 ( .A1(n662), .A2(n639), .ZN(n358) );
  XOR2_X1 U504 ( .A(n550), .B(n549), .Z(n359) );
  AND2_X1 U505 ( .A1(n482), .A2(n379), .ZN(n360) );
  AND2_X1 U506 ( .A1(n423), .A2(n358), .ZN(n361) );
  AND2_X1 U507 ( .A1(G227), .A2(n773), .ZN(n362) );
  OR2_X1 U508 ( .A1(n585), .A2(n584), .ZN(n363) );
  AND2_X1 U509 ( .A1(n607), .A2(n461), .ZN(n364) );
  OR2_X1 U510 ( .A1(n700), .A2(n701), .ZN(n365) );
  NOR2_X1 U511 ( .A1(n734), .A2(n371), .ZN(n366) );
  OR2_X1 U512 ( .A1(n484), .A2(KEYINPUT106), .ZN(n367) );
  NAND2_X1 U513 ( .A1(n479), .A2(n483), .ZN(n784) );
  XNOR2_X1 U514 ( .A(n439), .B(n438), .ZN(n786) );
  XOR2_X1 U515 ( .A(n666), .B(KEYINPUT62), .Z(n368) );
  XNOR2_X1 U516 ( .A(KEYINPUT15), .B(G902), .ZN(n665) );
  INV_X1 U517 ( .A(n664), .ZN(n430) );
  INV_X1 U518 ( .A(KEYINPUT80), .ZN(n414) );
  INV_X1 U519 ( .A(n598), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT48), .B(KEYINPUT86), .ZN(n598) );
  OR2_X1 U521 ( .A1(n665), .A2(n701), .ZN(n369) );
  AND2_X2 U522 ( .A1(n469), .A2(n365), .ZN(n370) );
  INV_X1 U523 ( .A(n602), .ZN(n489) );
  INV_X1 U524 ( .A(n622), .ZN(n482) );
  BUF_X1 U525 ( .A(n487), .Z(n371) );
  NOR2_X1 U526 ( .A1(n404), .A2(n396), .ZN(n395) );
  NOR2_X1 U527 ( .A1(n397), .A2(n395), .ZN(n394) );
  INV_X1 U528 ( .A(n640), .ZN(n782) );
  XNOR2_X1 U529 ( .A(n447), .B(n368), .ZN(n446) );
  NAND2_X1 U530 ( .A1(n418), .A2(n417), .ZN(n372) );
  NAND2_X1 U531 ( .A1(n418), .A2(n417), .ZN(n373) );
  NAND2_X1 U532 ( .A1(n418), .A2(n417), .ZN(n698) );
  XNOR2_X1 U533 ( .A(n380), .B(n559), .ZN(n562) );
  NOR2_X1 U534 ( .A1(n783), .A2(n784), .ZN(n374) );
  XNOR2_X2 U535 ( .A(n620), .B(n619), .ZN(n783) );
  XNOR2_X2 U536 ( .A(n614), .B(n613), .ZN(n626) );
  INV_X1 U537 ( .A(n725), .ZN(n375) );
  NOR2_X1 U538 ( .A1(n729), .A2(n375), .ZN(n376) );
  BUF_X1 U539 ( .A(n751), .Z(n377) );
  XNOR2_X1 U540 ( .A(n514), .B(n498), .ZN(n751) );
  NAND2_X1 U541 ( .A1(n370), .A2(G472), .ZN(n447) );
  NAND2_X1 U542 ( .A1(n666), .A2(G472), .ZN(n406) );
  XNOR2_X1 U543 ( .A(n500), .B(n466), .ZN(n496) );
  XNOR2_X2 U544 ( .A(n378), .B(G469), .ZN(n416) );
  NOR2_X1 U545 ( .A1(n751), .A2(G902), .ZN(n378) );
  BUF_X1 U546 ( .A(n712), .Z(n379) );
  INV_X1 U547 ( .A(n381), .ZN(n380) );
  XNOR2_X2 U548 ( .A(n493), .B(G143), .ZN(n381) );
  NAND2_X1 U549 ( .A1(n470), .A2(n369), .ZN(n469) );
  OR2_X2 U550 ( .A1(n416), .A2(n713), .ZN(n578) );
  XNOR2_X1 U551 ( .A(n416), .B(KEYINPUT1), .ZN(n712) );
  NAND2_X1 U552 ( .A1(n657), .A2(n656), .ZN(n423) );
  NAND2_X1 U553 ( .A1(n387), .A2(G475), .ZN(n670) );
  NAND2_X1 U554 ( .A1(n387), .A2(G210), .ZN(n747) );
  AND2_X2 U555 ( .A1(n421), .A2(n419), .ZN(n418) );
  NAND2_X1 U556 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U557 ( .A1(n370), .A2(G469), .ZN(n749) );
  NAND2_X1 U558 ( .A1(n370), .A2(G478), .ZN(n753) );
  NAND2_X1 U559 ( .A1(n370), .A2(G217), .ZN(n756) );
  OR2_X1 U560 ( .A1(n666), .A2(n402), .ZN(n401) );
  OR2_X1 U561 ( .A1(n666), .A2(n390), .ZN(n399) );
  INV_X1 U562 ( .A(n402), .ZN(n391) );
  NAND2_X1 U563 ( .A1(n394), .A2(n392), .ZN(n581) );
  NAND2_X1 U564 ( .A1(n393), .A2(n404), .ZN(n392) );
  AND2_X1 U565 ( .A1(n401), .A2(n577), .ZN(n393) );
  INV_X1 U566 ( .A(n400), .ZN(n396) );
  NAND2_X1 U567 ( .A1(n409), .A2(n407), .ZN(n413) );
  NAND2_X1 U568 ( .A1(n410), .A2(KEYINPUT80), .ZN(n409) );
  INV_X1 U569 ( .A(n415), .ZN(n410) );
  NOR2_X2 U570 ( .A1(n413), .A2(n411), .ZN(n464) );
  AND2_X1 U571 ( .A1(n415), .A2(n412), .ZN(n411) );
  AND2_X1 U572 ( .A1(n582), .A2(n414), .ZN(n412) );
  XNOR2_X1 U573 ( .A(n786), .B(KEYINPUT82), .ZN(n415) );
  XNOR2_X1 U574 ( .A(n416), .B(KEYINPUT109), .ZN(n573) );
  NAND2_X1 U575 ( .A1(n420), .A2(n430), .ZN(n419) );
  NAND2_X1 U576 ( .A1(n358), .A2(n424), .ZN(n420) );
  NAND2_X1 U577 ( .A1(n422), .A2(n430), .ZN(n421) );
  INV_X1 U578 ( .A(n423), .ZN(n422) );
  NAND2_X1 U579 ( .A1(n637), .A2(n638), .ZN(n424) );
  NOR2_X2 U580 ( .A1(n612), .A2(n611), .ZN(n614) );
  NOR2_X1 U581 ( .A1(n712), .A2(n713), .ZN(n627) );
  NAND2_X1 U582 ( .A1(n372), .A2(n354), .ZN(n471) );
  NAND2_X1 U583 ( .A1(n645), .A2(n431), .ZN(n491) );
  NOR2_X1 U584 ( .A1(n487), .A2(n626), .ZN(n631) );
  NAND2_X1 U585 ( .A1(n640), .A2(n660), .ZN(n651) );
  NAND2_X1 U586 ( .A1(n782), .A2(KEYINPUT89), .ZN(n639) );
  XNOR2_X1 U587 ( .A(n471), .B(KEYINPUT84), .ZN(n470) );
  BUF_X1 U588 ( .A(n623), .Z(n719) );
  NOR2_X2 U589 ( .A1(n590), .A2(n383), .ZN(n685) );
  XNOR2_X1 U590 ( .A(n377), .B(n750), .ZN(n434) );
  NOR2_X1 U591 ( .A1(n605), .A2(n596), .ZN(n597) );
  XNOR2_X1 U592 ( .A(n437), .B(n673), .ZN(G60) );
  NOR2_X2 U593 ( .A1(n671), .A2(n758), .ZN(n437) );
  XNOR2_X1 U594 ( .A(n440), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U595 ( .A1(n748), .A2(n758), .ZN(n440) );
  AND2_X1 U596 ( .A1(n464), .A2(n453), .ZN(n441) );
  NAND2_X1 U597 ( .A1(n444), .A2(n443), .ZN(n442) );
  XNOR2_X1 U598 ( .A(n445), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U599 ( .A1(n446), .A2(n667), .ZN(n445) );
  NOR2_X1 U600 ( .A1(n468), .A2(G902), .ZN(n545) );
  XNOR2_X1 U601 ( .A(n756), .B(n468), .ZN(n757) );
  NAND2_X1 U602 ( .A1(n698), .A2(n772), .ZN(n700) );
  NAND2_X1 U603 ( .A1(n622), .A2(n486), .ZN(n485) );
  INV_X1 U604 ( .A(KEYINPUT106), .ZN(n486) );
  XNOR2_X2 U605 ( .A(n771), .B(G146), .ZN(n514) );
  XNOR2_X2 U606 ( .A(n501), .B(n495), .ZN(n771) );
  NOR2_X1 U607 ( .A1(n371), .A2(n724), .ZN(n707) );
  XNOR2_X1 U608 ( .A(n630), .B(n629), .ZN(n487) );
  NAND2_X1 U609 ( .A1(n632), .A2(n489), .ZN(n488) );
  INV_X1 U610 ( .A(n665), .ZN(n529) );
  XNOR2_X1 U611 ( .A(n492), .B(KEYINPUT20), .ZN(n530) );
  NAND2_X1 U612 ( .A1(n665), .A2(G234), .ZN(n492) );
  NOR2_X2 U613 ( .A1(n529), .A2(n745), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X2 U615 ( .A(n578), .B(KEYINPUT97), .ZN(n645) );
  OR2_X2 U616 ( .A1(n709), .A2(n624), .ZN(n713) );
  XNOR2_X1 U617 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U618 ( .A(n518), .B(G131), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n663), .B(KEYINPUT45), .ZN(n664) );
  INV_X1 U620 ( .A(KEYINPUT79), .ZN(n509) );
  INV_X1 U621 ( .A(n624), .ZN(n625) );
  XNOR2_X1 U622 ( .A(n510), .B(n509), .ZN(n511) );
  INV_X1 U623 ( .A(KEYINPUT19), .ZN(n574) );
  INV_X1 U624 ( .A(n758), .ZN(n667) );
  XNOR2_X1 U625 ( .A(n618), .B(KEYINPUT32), .ZN(n619) );
  XNOR2_X1 U626 ( .A(n672), .B(KEYINPUT60), .ZN(n673) );
  XNOR2_X2 U627 ( .A(G128), .B(KEYINPUT65), .ZN(n493) );
  XNOR2_X1 U628 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n494) );
  XNOR2_X1 U629 ( .A(G101), .B(KEYINPUT75), .ZN(n497) );
  XNOR2_X1 U630 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U631 ( .A(n501), .B(n765), .ZN(n508) );
  XNOR2_X1 U632 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U633 ( .A(n536), .B(n504), .Z(n506) );
  NAND2_X1 U634 ( .A1(G224), .A2(n773), .ZN(n505) );
  XNOR2_X1 U635 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U636 ( .A(n508), .B(n507), .ZN(n745) );
  NAND2_X1 U637 ( .A1(G210), .A2(n513), .ZN(n510) );
  XNOR2_X2 U638 ( .A(n512), .B(n511), .ZN(n588) );
  NAND2_X1 U639 ( .A1(G214), .A2(n513), .ZN(n725) );
  XNOR2_X1 U640 ( .A(n515), .B(KEYINPUT72), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n553), .A2(G210), .ZN(n517) );
  INV_X1 U642 ( .A(G472), .ZN(n521) );
  INV_X1 U643 ( .A(n628), .ZN(n659) );
  XNOR2_X1 U644 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U645 ( .A(KEYINPUT70), .B(n524), .ZN(n525) );
  NAND2_X1 U646 ( .A1(G952), .A2(n525), .ZN(n739) );
  NOR2_X1 U647 ( .A1(G953), .A2(n739), .ZN(n610) );
  NAND2_X1 U648 ( .A1(G902), .A2(n525), .ZN(n608) );
  NOR2_X1 U649 ( .A1(G900), .A2(n608), .ZN(n526) );
  NAND2_X1 U650 ( .A1(G953), .A2(n526), .ZN(n527) );
  XNOR2_X1 U651 ( .A(KEYINPUT107), .B(n527), .ZN(n528) );
  NOR2_X1 U652 ( .A1(n610), .A2(n528), .ZN(n579) );
  XNOR2_X1 U653 ( .A(KEYINPUT96), .B(n530), .ZN(n541) );
  NAND2_X1 U654 ( .A1(n541), .A2(G221), .ZN(n531) );
  XNOR2_X1 U655 ( .A(n531), .B(KEYINPUT21), .ZN(n709) );
  NOR2_X1 U656 ( .A1(n579), .A2(n709), .ZN(n546) );
  XOR2_X1 U657 ( .A(KEYINPUT24), .B(G140), .Z(n533) );
  XNOR2_X1 U658 ( .A(G110), .B(G128), .ZN(n532) );
  XNOR2_X1 U659 ( .A(n533), .B(n532), .ZN(n534) );
  NAND2_X1 U660 ( .A1(n773), .A2(G234), .ZN(n539) );
  XNOR2_X1 U661 ( .A(n539), .B(n538), .ZN(n560) );
  NAND2_X1 U662 ( .A1(n560), .A2(G221), .ZN(n540) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(KEYINPUT25), .Z(n543) );
  NAND2_X1 U664 ( .A1(G217), .A2(n541), .ZN(n542) );
  XNOR2_X1 U665 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U666 ( .A1(n546), .A2(n624), .ZN(n570) );
  XNOR2_X1 U667 ( .A(n548), .B(n547), .ZN(n770) );
  NAND2_X1 U668 ( .A1(G214), .A2(n553), .ZN(n554) );
  NOR2_X1 U669 ( .A1(G902), .A2(n668), .ZN(n556) );
  INV_X1 U670 ( .A(n586), .ZN(n567) );
  XNOR2_X1 U671 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n566) );
  XOR2_X1 U672 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n558) );
  XNOR2_X1 U673 ( .A(G134), .B(G107), .ZN(n557) );
  XNOR2_X1 U674 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U675 ( .A1(G217), .A2(n560), .ZN(n561) );
  XNOR2_X1 U676 ( .A(n564), .B(n563), .ZN(n754) );
  NOR2_X1 U677 ( .A1(G902), .A2(n754), .ZN(n565) );
  INV_X1 U678 ( .A(n569), .ZN(n587) );
  NOR2_X1 U679 ( .A1(n570), .A2(n596), .ZN(n568) );
  NAND2_X1 U680 ( .A1(n659), .A2(n568), .ZN(n599) );
  INV_X1 U681 ( .A(n596), .ZN(n687) );
  NAND2_X1 U682 ( .A1(n586), .A2(n569), .ZN(n604) );
  INV_X1 U683 ( .A(n604), .ZN(n689) );
  XNOR2_X1 U684 ( .A(KEYINPUT28), .B(n571), .ZN(n572) );
  NAND2_X1 U685 ( .A1(n573), .A2(n572), .ZN(n590) );
  INV_X1 U686 ( .A(n685), .ZN(n585) );
  OR2_X1 U687 ( .A1(n731), .A2(n585), .ZN(n576) );
  NAND2_X1 U688 ( .A1(n576), .A2(KEYINPUT47), .ZN(n582) );
  INV_X1 U689 ( .A(KEYINPUT30), .ZN(n577) );
  INV_X1 U690 ( .A(n579), .ZN(n580) );
  INV_X1 U691 ( .A(n588), .ZN(n602) );
  NOR2_X1 U692 ( .A1(n587), .A2(n586), .ZN(n632) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n731), .Z(n648) );
  NOR2_X1 U694 ( .A1(KEYINPUT47), .A2(n648), .ZN(n583) );
  XNOR2_X1 U695 ( .A(KEYINPUT69), .B(n583), .ZN(n584) );
  NAND2_X1 U696 ( .A1(n587), .A2(n586), .ZN(n729) );
  XNOR2_X1 U697 ( .A(n589), .B(KEYINPUT41), .ZN(n724) );
  NOR2_X1 U698 ( .A1(n590), .A2(n724), .ZN(n591) );
  XNOR2_X1 U699 ( .A(n591), .B(KEYINPUT42), .ZN(n787) );
  INV_X1 U700 ( .A(n726), .ZN(n592) );
  XNOR2_X1 U701 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n594) );
  XNOR2_X1 U702 ( .A(n595), .B(n594), .ZN(n605) );
  XNOR2_X1 U703 ( .A(n597), .B(KEYINPUT40), .ZN(n785) );
  INV_X1 U704 ( .A(n379), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n621), .A2(n599), .ZN(n600) );
  NAND2_X1 U706 ( .A1(n600), .A2(n725), .ZN(n601) );
  XNOR2_X1 U707 ( .A(n601), .B(KEYINPUT43), .ZN(n603) );
  NAND2_X1 U708 ( .A1(n603), .A2(n602), .ZN(n697) );
  NOR2_X1 U709 ( .A1(n605), .A2(n604), .ZN(n695) );
  INV_X1 U710 ( .A(n695), .ZN(n606) );
  AND2_X1 U711 ( .A1(n697), .A2(n606), .ZN(n607) );
  INV_X1 U712 ( .A(n729), .ZN(n615) );
  OR2_X1 U713 ( .A1(n773), .A2(G898), .ZN(n767) );
  NOR2_X1 U714 ( .A1(n608), .A2(n767), .ZN(n609) );
  NOR2_X1 U715 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U716 ( .A(KEYINPUT0), .ZN(n613) );
  XNOR2_X1 U717 ( .A(KEYINPUT105), .B(n624), .ZN(n710) );
  NOR2_X1 U718 ( .A1(n379), .A2(n659), .ZN(n616) );
  NAND2_X1 U719 ( .A1(n617), .A2(n616), .ZN(n620) );
  INV_X1 U720 ( .A(KEYINPUT78), .ZN(n618) );
  NOR2_X2 U721 ( .A1(n783), .A2(n784), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT90), .ZN(n638) );
  INV_X1 U723 ( .A(KEYINPUT44), .ZN(n636) );
  INV_X1 U724 ( .A(n626), .ZN(n644) );
  XNOR2_X1 U725 ( .A(n627), .B(KEYINPUT71), .ZN(n641) );
  NOR2_X1 U726 ( .A1(n641), .A2(n628), .ZN(n630) );
  XOR2_X1 U727 ( .A(KEYINPUT91), .B(KEYINPUT33), .Z(n629) );
  XNOR2_X1 U728 ( .A(n631), .B(KEYINPUT34), .ZN(n634) );
  XOR2_X1 U729 ( .A(n632), .B(KEYINPUT77), .Z(n633) );
  INV_X1 U730 ( .A(KEYINPUT89), .ZN(n660) );
  NOR2_X1 U731 ( .A1(n641), .A2(n642), .ZN(n721) );
  NAND2_X1 U732 ( .A1(n721), .A2(n644), .ZN(n643) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U734 ( .A1(n719), .A2(n646), .ZN(n677) );
  NOR2_X1 U735 ( .A1(n690), .A2(n677), .ZN(n647) );
  XNOR2_X1 U736 ( .A(n647), .B(KEYINPUT99), .ZN(n650) );
  INV_X1 U737 ( .A(n648), .ZN(n649) );
  NAND2_X1 U738 ( .A1(n650), .A2(n649), .ZN(n654) );
  AND2_X1 U739 ( .A1(n651), .A2(n654), .ZN(n652) );
  NAND2_X1 U740 ( .A1(n374), .A2(n652), .ZN(n657) );
  INV_X1 U741 ( .A(n654), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n360), .A2(n710), .ZN(n658) );
  NOR2_X1 U743 ( .A1(n659), .A2(n658), .ZN(n674) );
  NOR2_X1 U744 ( .A1(KEYINPUT44), .A2(n660), .ZN(n661) );
  NOR2_X1 U745 ( .A1(n674), .A2(n661), .ZN(n662) );
  XNOR2_X1 U746 ( .A(KEYINPUT64), .B(KEYINPUT85), .ZN(n663) );
  INV_X1 U747 ( .A(KEYINPUT2), .ZN(n701) );
  XNOR2_X1 U748 ( .A(n670), .B(n669), .ZN(n671) );
  INV_X1 U749 ( .A(KEYINPUT121), .ZN(n672) );
  XNOR2_X1 U750 ( .A(G101), .B(n674), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n675), .B(KEYINPUT111), .ZN(G3) );
  NAND2_X1 U752 ( .A1(n677), .A2(n687), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(G104), .ZN(G6) );
  XNOR2_X1 U754 ( .A(G107), .B(KEYINPUT112), .ZN(n681) );
  XOR2_X1 U755 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n679) );
  NAND2_X1 U756 ( .A1(n677), .A2(n689), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U758 ( .A(n681), .B(n680), .ZN(G9) );
  XOR2_X1 U759 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n683) );
  NAND2_X1 U760 ( .A1(n689), .A2(n685), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n683), .B(n682), .ZN(n684) );
  XOR2_X1 U762 ( .A(G128), .B(n684), .Z(G30) );
  NAND2_X1 U763 ( .A1(n685), .A2(n687), .ZN(n686) );
  XNOR2_X1 U764 ( .A(n686), .B(G146), .ZN(G48) );
  NAND2_X1 U765 ( .A1(n687), .A2(n690), .ZN(n688) );
  XNOR2_X1 U766 ( .A(G113), .B(n688), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U768 ( .A(n691), .B(KEYINPUT114), .ZN(n692) );
  XNOR2_X1 U769 ( .A(G116), .B(n692), .ZN(G18) );
  XNOR2_X1 U770 ( .A(G125), .B(n693), .ZN(n694) );
  XNOR2_X1 U771 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U772 ( .A(G134), .B(n695), .ZN(n696) );
  XNOR2_X1 U773 ( .A(n696), .B(KEYINPUT115), .ZN(G36) );
  XNOR2_X1 U774 ( .A(G140), .B(n697), .ZN(G42) );
  XNOR2_X1 U775 ( .A(n699), .B(KEYINPUT83), .ZN(n703) );
  OR2_X1 U776 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U777 ( .A1(n703), .A2(n702), .ZN(n705) );
  NOR2_X1 U778 ( .A1(KEYINPUT2), .A2(n772), .ZN(n704) );
  NOR2_X1 U779 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U780 ( .A(KEYINPUT120), .B(n707), .Z(n708) );
  NOR2_X1 U781 ( .A1(n710), .A2(n426), .ZN(n711) );
  XNOR2_X1 U782 ( .A(KEYINPUT49), .B(n711), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n713), .A2(n379), .ZN(n714) );
  XNOR2_X1 U784 ( .A(n714), .B(KEYINPUT50), .ZN(n715) );
  XNOR2_X1 U785 ( .A(KEYINPUT116), .B(n715), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U789 ( .A(KEYINPUT51), .B(n722), .Z(n723) );
  NOR2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n735) );
  NOR2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U792 ( .A(KEYINPUT117), .B(n727), .Z(n728) );
  NOR2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n733) );
  NOR2_X1 U794 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U795 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U796 ( .A1(n735), .A2(n366), .ZN(n736) );
  XNOR2_X1 U797 ( .A(n736), .B(KEYINPUT52), .ZN(n737) );
  XNOR2_X1 U798 ( .A(KEYINPUT118), .B(n737), .ZN(n738) );
  NOR2_X1 U799 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U800 ( .A(KEYINPUT119), .B(n740), .Z(n741) );
  NOR2_X1 U801 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U802 ( .A(KEYINPUT53), .B(n743), .ZN(G75) );
  XOR2_X1 U803 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n744) );
  XNOR2_X1 U804 ( .A(n745), .B(n744), .ZN(n746) );
  XOR2_X1 U805 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n750) );
  NOR2_X1 U806 ( .A1(n758), .A2(n752), .ZN(G54) );
  NOR2_X1 U807 ( .A1(n758), .A2(n755), .ZN(G63) );
  NOR2_X1 U808 ( .A1(n758), .A2(n757), .ZN(G66) );
  XOR2_X1 U809 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n760) );
  NAND2_X1 U810 ( .A1(G224), .A2(G953), .ZN(n759) );
  XNOR2_X1 U811 ( .A(n760), .B(n759), .ZN(n761) );
  NAND2_X1 U812 ( .A1(n761), .A2(G898), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n373), .A2(n773), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U815 ( .A(n764), .B(KEYINPUT125), .ZN(n769) );
  XOR2_X1 U816 ( .A(n765), .B(KEYINPUT124), .Z(n766) );
  NAND2_X1 U817 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U818 ( .A(n769), .B(n768), .ZN(G69) );
  XOR2_X1 U819 ( .A(n771), .B(n770), .Z(n775) );
  XOR2_X1 U820 ( .A(n772), .B(n775), .Z(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n781) );
  XNOR2_X1 U822 ( .A(G227), .B(KEYINPUT126), .ZN(n776) );
  XNOR2_X1 U823 ( .A(n776), .B(n775), .ZN(n777) );
  NAND2_X1 U824 ( .A1(G900), .A2(n777), .ZN(n778) );
  XOR2_X1 U825 ( .A(KEYINPUT127), .B(n778), .Z(n779) );
  NAND2_X1 U826 ( .A1(G953), .A2(n779), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n781), .A2(n780), .ZN(G72) );
  XNOR2_X1 U828 ( .A(n782), .B(G122), .ZN(G24) );
  XOR2_X1 U829 ( .A(n783), .B(G119), .Z(G21) );
  XOR2_X1 U830 ( .A(G110), .B(n784), .Z(G12) );
  XOR2_X1 U831 ( .A(n785), .B(G131), .Z(G33) );
  XNOR2_X1 U832 ( .A(G143), .B(n786), .ZN(G45) );
  XOR2_X1 U833 ( .A(n787), .B(G137), .Z(G39) );
endmodule

