//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT65), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n463), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G2105), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(KEYINPUT66), .A3(KEYINPUT3), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n465), .B2(G2104), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  AND3_X1   g054(.A1(new_n476), .A2(new_n472), .A3(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n483), .A3(new_n474), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n480), .A2(G124), .A3(G2105), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT68), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n474), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n500));
  OR3_X1    g075(.A1(new_n499), .A2(new_n467), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n476), .A2(new_n472), .A3(new_n496), .A4(new_n466), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT4), .B1(new_n502), .B2(KEYINPUT70), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n474), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n473), .A2(G2105), .A3(new_n476), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G126), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT72), .B(G88), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND2_X1  g104(.A1(new_n522), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(new_n531), .B1(new_n516), .B2(new_n517), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT73), .B(G51), .Z(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  INV_X1    g112(.A(new_n525), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n516), .B2(new_n517), .ZN(new_n541));
  AND2_X1   g116(.A1(G77), .A2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n518), .A2(new_n522), .A3(G90), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n520), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n523), .A2(new_n549), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n522), .A2(G53), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n561), .A2(new_n520), .B1(new_n562), .B2(new_n523), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(new_n523), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n538), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G73), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n515), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n518), .A2(G61), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n516), .B2(new_n517), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n520), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n523), .A2(new_n581), .B1(new_n525), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n520), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n523), .A2(new_n588), .B1(new_n525), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n520), .B1(new_n595), .B2(new_n525), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI221_X1 g173(.A(KEYINPUT76), .B1(new_n525), .B2(new_n595), .C1(new_n594), .C2(new_n520), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g175(.A1(new_n518), .A2(new_n522), .A3(G92), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n564), .ZN(G280));
  XOR2_X1   g184(.A(G280), .B(KEYINPUT77), .Z(G297));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n605), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND2_X1  g187(.A1(new_n605), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g191(.A1(new_n510), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n474), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(new_n617), .B1(new_n618), .B2(new_n619), .C1(new_n485), .C2(new_n620), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(G2096), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(G2096), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n622), .A2(new_n623), .A3(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT79), .Z(new_n642));
  NOR2_X1   g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n639), .A2(KEYINPUT78), .A3(new_n640), .ZN(new_n646));
  OAI21_X1  g221(.A(G14), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n642), .A2(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT80), .ZN(new_n651));
  NOR2_X1   g226(.A1(G2072), .A2(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n442), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n649), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(KEYINPUT17), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n649), .B(new_n650), .C1(new_n442), .C2(new_n652), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n651), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT81), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n669), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n676), .C1(new_n666), .C2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT84), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n681), .B2(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n664), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n663), .A3(new_n686), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NOR2_X1   g268(.A1(G162), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(G35), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT29), .ZN(new_n696));
  INV_X1    g271(.A(G2090), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n693), .A2(G32), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n510), .A2(G129), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n486), .A2(G141), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT26), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n707), .A2(new_n708), .B1(G105), .B2(new_n470), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n703), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT92), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n701), .B1(new_n711), .B2(new_n693), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT93), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n700), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n698), .A2(new_n699), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n717), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1971), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n584), .A2(G16), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G6), .B2(G16), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT32), .B(G1981), .Z(new_n723));
  AOI21_X1  g298(.A(new_n720), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(G16), .A2(G23), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT85), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G288), .B2(new_n717), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT33), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1976), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n724), .B(new_n729), .C1(new_n722), .C2(new_n723), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n732));
  NOR2_X1   g307(.A1(G25), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n486), .A2(G131), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  INV_X1    g310(.A(G107), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n510), .B2(G119), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(G29), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT35), .B(G1991), .Z(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n717), .A2(G24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n591), .B2(new_n717), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1986), .ZN(new_n747));
  INV_X1    g322(.A(new_n741), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n742), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n731), .A2(new_n732), .A3(new_n744), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT36), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(KEYINPUT86), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n717), .A2(G4), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n605), .B2(new_n717), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT87), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1348), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n717), .A2(G20), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT23), .Z(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G299), .B2(G16), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1956), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n717), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n717), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1961), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n717), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n717), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n717), .A2(G19), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n552), .B2(new_n717), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1341), .Z(new_n771));
  NAND3_X1  g346(.A1(new_n764), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT24), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(G34), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n478), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n761), .B(new_n772), .C1(G2084), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(G2084), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT97), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n757), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n693), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  INV_X1    g360(.A(G139), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n485), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT88), .ZN(new_n788));
  NAND2_X1  g363(.A1(G115), .A2(G2104), .ZN(new_n789));
  INV_X1    g364(.A(G127), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n467), .B2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(KEYINPUT89), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n474), .B1(new_n791), .B2(KEYINPUT89), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n788), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n783), .B1(new_n794), .B2(new_n693), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G2072), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n693), .A2(G26), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT28), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n486), .A2(G140), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n800));
  INV_X1    g375(.A(G116), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(G2105), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n510), .B2(G128), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(G29), .ZN(new_n805));
  INV_X1    g380(.A(G2067), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G164), .A2(new_n693), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G27), .B2(new_n693), .ZN(new_n809));
  INV_X1    g384(.A(G2078), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n796), .B(new_n812), .C1(new_n810), .C2(new_n809), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n795), .A2(G2072), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n621), .A2(KEYINPUT95), .A3(new_n693), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT95), .B1(new_n621), .B2(new_n693), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT30), .B(G28), .ZN(new_n817));
  OR2_X1    g392(.A1(KEYINPUT31), .A2(G11), .ZN(new_n818));
  NAND2_X1  g393(.A1(KEYINPUT31), .A2(G11), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n817), .A2(new_n693), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n815), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT96), .Z(new_n822));
  NOR4_X1   g397(.A1(new_n782), .A2(new_n813), .A3(new_n814), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n713), .A2(new_n700), .A3(new_n714), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT94), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n716), .A2(new_n753), .A3(new_n823), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NOR2_X1   g402(.A1(new_n604), .A2(new_n611), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT38), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(new_n520), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n518), .A2(new_n522), .A3(G93), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n522), .A2(G55), .A3(G543), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n834), .B1(new_n832), .B2(new_n833), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n548), .B2(new_n551), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n552), .B(new_n831), .C1(new_n835), .C2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n829), .B(new_n840), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n837), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  INV_X1    g422(.A(KEYINPUT40), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n794), .A2(new_n710), .ZN(new_n849));
  INV_X1    g424(.A(new_n711), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n794), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(G118), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(G2105), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n510), .B2(G130), .ZN(new_n855));
  INV_X1    g430(.A(G142), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n485), .B2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n625), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n739), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(new_n501), .C1(new_n504), .C2(new_n505), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT70), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n473), .A2(new_n863), .A3(new_n476), .A4(new_n496), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(KEYINPUT4), .A3(new_n503), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n865), .B2(new_n501), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n511), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n859), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n858), .B(new_n740), .ZN(new_n869));
  INV_X1    g444(.A(new_n511), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n506), .A2(KEYINPUT99), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n861), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n804), .B(KEYINPUT100), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n868), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n875), .B1(new_n873), .B2(new_n868), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n851), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n621), .B(new_n478), .ZN(new_n880));
  XOR2_X1   g455(.A(G162), .B(new_n880), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n868), .A2(new_n873), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n874), .ZN(new_n883));
  INV_X1    g458(.A(new_n851), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n883), .A2(new_n884), .A3(new_n876), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n881), .B1(new_n879), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n848), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n887), .A4(new_n886), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(G395));
  XNOR2_X1  g468(.A(G288), .B(KEYINPUT101), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n584), .ZN(new_n895));
  XNOR2_X1  g470(.A(G290), .B(G303), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n894), .B(G305), .ZN(new_n898));
  INV_X1    g473(.A(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT42), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n613), .B(new_n840), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT41), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n600), .A2(new_n564), .A3(new_n603), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n564), .B1(new_n600), .B2(new_n603), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n604), .A2(G299), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n600), .A2(new_n564), .A3(new_n603), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n905), .A2(new_n906), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n903), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n902), .B(new_n914), .ZN(new_n915));
  MUX2_X1   g490(.A(new_n837), .B(new_n915), .S(G868), .Z(G295));
  MUX2_X1   g491(.A(new_n837), .B(new_n915), .S(G868), .Z(G331));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n539), .A2(KEYINPUT102), .A3(new_n543), .A4(new_n544), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n919), .A2(G168), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n919), .B2(G168), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n840), .ZN(new_n924));
  NOR2_X1   g499(.A1(G171), .A2(KEYINPUT102), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n838), .B(new_n839), .C1(new_n921), .C2(new_n922), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n913), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n926), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n933), .A2(new_n907), .A3(new_n910), .A4(new_n927), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n928), .A2(new_n929), .A3(new_n911), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n901), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n901), .B1(new_n937), .B2(KEYINPUT105), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n930), .A2(new_n934), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n940), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  INV_X1    g524(.A(new_n901), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n936), .A2(new_n938), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n936), .B2(new_n938), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n951), .A2(new_n952), .A3(G37), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n918), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n947), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n946), .B1(new_n941), .B2(new_n943), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n954), .B1(new_n959), .B2(new_n940), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n936), .A2(new_n938), .A3(new_n950), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n940), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n918), .B1(new_n953), .B2(new_n954), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT107), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n956), .B1(new_n965), .B2(new_n968), .ZN(G397));
  NOR2_X1   g544(.A1(new_n872), .A2(G1384), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n469), .A2(G2105), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n470), .A2(G101), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(G40), .A3(new_n477), .A4(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT109), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n471), .A2(new_n978), .A3(G40), .A4(new_n477), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n711), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n804), .A2(G2067), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n799), .A2(new_n806), .A3(new_n803), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(G1996), .B2(new_n710), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n739), .A2(new_n743), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n740), .A2(new_n742), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n984), .A2(new_n988), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n591), .B(G1986), .Z(new_n992));
  OAI21_X1  g567(.A(new_n982), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT114), .B1(KEYINPUT115), .B2(KEYINPUT49), .ZN(new_n994));
  OAI21_X1  g569(.A(G1981), .B1(new_n580), .B2(new_n583), .ZN(new_n995));
  INV_X1    g570(.A(new_n579), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n578), .A2(KEYINPUT74), .B1(new_n572), .B2(new_n515), .ZN(new_n997));
  OAI21_X1  g572(.A(G651), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n583), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n994), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n995), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  AND2_X1   g580(.A1(new_n1005), .A2(KEYINPUT115), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1003), .B1(new_n1006), .B2(KEYINPUT49), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT112), .B(G8), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n970), .B2(new_n980), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n867), .A2(new_n980), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1008), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n568), .A2(new_n569), .A3(G1976), .A4(new_n570), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1007), .A2(new_n1009), .B1(new_n1014), .B2(KEYINPUT52), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  INV_X1    g591(.A(G1971), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n872), .A2(new_n1018), .A3(G1384), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n506), .B2(new_n511), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n980), .B1(new_n972), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1017), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n867), .A2(new_n1023), .A3(new_n1010), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n977), .A2(new_n979), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n512), .A2(new_n1010), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n1027), .A3(new_n697), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1016), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT55), .B(G8), .C1(new_n521), .C2(new_n527), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(KEYINPUT110), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(KEYINPUT111), .A3(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(G166), .B2(new_n1016), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT113), .B(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .A4(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1015), .A2(new_n1029), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT49), .B1(new_n1005), .B2(KEYINPUT115), .ZN(new_n1044));
  NOR4_X1   g619(.A1(new_n1044), .A2(G1976), .A3(G288), .A4(new_n1002), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1001), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1009), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT116), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1028), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n1010), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1025), .B1(new_n1026), .B2(new_n971), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1971), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(new_n1039), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1011), .B(new_n1012), .C1(new_n1044), .C2(new_n1002), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1042), .A3(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1047), .B(KEYINPUT116), .C1(new_n1053), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1048), .A2(new_n1058), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1060));
  AOI21_X1  g635(.A(new_n1025), .B1(new_n1023), .B2(new_n1020), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n697), .B(new_n1061), .C1(new_n970), .C2(new_n1023), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1008), .B1(new_n1022), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT117), .B1(new_n1063), .B2(new_n1039), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1023), .B1(new_n867), .B2(new_n1010), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n980), .B1(KEYINPUT50), .B2(new_n1026), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1065), .A2(new_n1066), .A3(G2090), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1012), .B1(new_n1067), .B2(new_n1052), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1039), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1056), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1064), .A2(new_n1071), .A3(new_n1053), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G2084), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1024), .A2(new_n1027), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1018), .B1(new_n872), .B2(G1384), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1025), .B1(new_n972), .B2(new_n1020), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1966), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(G168), .B(new_n1012), .C1(new_n1076), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT118), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT45), .B1(new_n867), .B2(new_n1010), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n980), .B1(new_n971), .B2(new_n1026), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n767), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1008), .B1(new_n1084), .B2(new_n1075), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(G168), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1060), .B1(new_n1073), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1053), .A2(KEYINPUT63), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1070), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1093), .A2(KEYINPUT120), .A3(new_n1072), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT120), .B1(new_n1093), .B2(new_n1072), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1091), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1059), .B1(new_n1089), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(G1956), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1050), .A2(new_n1051), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n564), .B(KEYINPUT57), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n872), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n980), .B1(new_n1023), .B2(new_n1020), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G1348), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1024), .A2(new_n1027), .A3(KEYINPUT122), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n970), .A2(new_n806), .A3(new_n980), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1099), .A2(new_n1103), .A3(new_n1101), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n605), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1105), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n605), .B2(KEYINPUT125), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1112), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n605), .A2(KEYINPUT125), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT60), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1115), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1103), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1105), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1112), .A2(new_n1113), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1050), .A2(new_n1051), .A3(new_n983), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1011), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1134), .A2(KEYINPUT123), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT123), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n552), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1117), .B1(new_n1133), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1012), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G168), .A2(new_n1008), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1149), .A2(KEYINPUT51), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1016), .B1(new_n1084), .B2(new_n1075), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT51), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1153));
  AOI211_X1 g728(.A(G168), .B(new_n1008), .C1(new_n1084), .C2(new_n1075), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1064), .A2(new_n1071), .A3(new_n1053), .A4(new_n1072), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT126), .B(G1961), .Z(new_n1158));
  NAND3_X1  g733(.A1(new_n1109), .A2(new_n1111), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1050), .A2(new_n1051), .A3(new_n810), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1159), .B(new_n1162), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(G301), .B(KEYINPUT54), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n973), .A2(new_n976), .A3(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1168), .B2(new_n1050), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1165), .A2(new_n1166), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1156), .A2(new_n1157), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1097), .B1(new_n1147), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT62), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1155), .A2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g749(.A(KEYINPUT62), .B(new_n1151), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1165), .A2(G171), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1174), .A2(new_n1157), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(KEYINPUT127), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1073), .A2(new_n1176), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1175), .A4(new_n1174), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n993), .B1(new_n1172), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n982), .A2(new_n983), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1185), .B(KEYINPUT46), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n982), .B1(new_n710), .B2(new_n987), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  OR3_X1    g764(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(KEYINPUT48), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n991), .A2(new_n982), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(KEYINPUT48), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n984), .A2(new_n988), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n986), .B1(new_n1196), .B2(new_n990), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1197), .A2(new_n982), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1189), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1184), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g775(.A1(G227), .A2(new_n460), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1202), .B1(new_n642), .B2(new_n647), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n689), .B2(new_n691), .ZN(new_n1204));
  OAI21_X1  g778(.A(new_n1204), .B1(new_n888), .B2(new_n889), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n949), .A2(new_n955), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n1206), .ZN(G308));
  OR2_X1    g781(.A1(new_n1205), .A2(new_n1206), .ZN(G225));
endmodule


