//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(KEYINPUT66), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT66), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G20), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G20), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(G250), .B1(G257), .B2(G264), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n222), .B1(new_n228), .B2(KEYINPUT0), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT67), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(KEYINPUT67), .B1(new_n230), .B2(new_n231), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n224), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT1), .ZN(new_n238));
  AOI211_X1 g0038(.A(new_n229), .B(new_n238), .C1(KEYINPUT0), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  INV_X1    g0040(.A(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G358));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G97), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n253), .B(new_n254), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(KEYINPUT9), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n215), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT74), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT72), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n217), .A3(KEYINPUT8), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT8), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT72), .B1(new_n264), .B2(G58), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n217), .A2(KEYINPUT8), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT73), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n269), .B(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n271), .B1(new_n211), .B2(new_n213), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n261), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n210), .B1(new_n201), .B2(new_n202), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n273), .A2(new_n261), .A3(new_n275), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n260), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n259), .B1(new_n281), .B2(G20), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G50), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n257), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n279), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n276), .A3(new_n277), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT9), .B(new_n285), .C1(new_n289), .C2(new_n260), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G222), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT70), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT3), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G33), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n296), .A2(new_n298), .A3(new_n292), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n300), .A3(G222), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n291), .A2(G223), .A3(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G77), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n295), .A2(new_n301), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n281), .B(G274), .C1(G41), .C2(G45), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  INV_X1    g0110(.A(G45), .ZN(new_n311));
  AOI21_X1  g0111(.A(G1), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G41), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n215), .B1(KEYINPUT69), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G33), .A3(G41), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n309), .B1(new_n317), .B2(G226), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n307), .A2(KEYINPUT71), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(G200), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n318), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n320), .B(new_n324), .C1(new_n305), .C2(new_n306), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT71), .B1(new_n307), .B2(new_n318), .ZN(new_n326));
  OAI21_X1  g0126(.A(G190), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n287), .A2(new_n290), .A3(new_n323), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT10), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n327), .A2(new_n323), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT10), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n290), .A4(new_n287), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n268), .A2(new_n270), .ZN(new_n334));
  INV_X1    g0134(.A(new_n284), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n282), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n336), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT82), .ZN(new_n339));
  AOI21_X1  g0139(.A(G20), .B1(new_n296), .B2(new_n298), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(KEYINPUT7), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT82), .B(new_n342), .C1(new_n291), .C2(G20), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n214), .A2(new_n303), .A3(KEYINPUT7), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT81), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G58), .A2(G68), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n210), .B1(new_n219), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n274), .A2(G159), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n347), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n348), .ZN(new_n353));
  OAI21_X1  g0153(.A(G20), .B1(new_n353), .B2(new_n201), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(KEYINPUT81), .A3(new_n350), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT16), .B1(new_n346), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT7), .B1(new_n291), .B2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n214), .A2(new_n303), .A3(new_n342), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(G68), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n352), .A4(new_n355), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n259), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n338), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n309), .B1(new_n317), .B2(G232), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n296), .A2(new_n298), .A3(G226), .A4(G1698), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n296), .A2(new_n298), .A3(G223), .A4(new_n292), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G33), .A2(G87), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n306), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n364), .A2(new_n369), .A3(G179), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n364), .B2(new_n369), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n352), .A2(new_n355), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n345), .B2(G68), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n259), .B(new_n361), .C1(new_n379), .C2(KEYINPUT16), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n373), .B1(new_n380), .B2(new_n338), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G200), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n364), .B2(new_n369), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n364), .A2(new_n369), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(G190), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(new_n387), .A3(new_n338), .ZN(new_n388));
  XNOR2_X1  g0188(.A(new_n388), .B(KEYINPUT17), .ZN(new_n389));
  XOR2_X1   g0189(.A(KEYINPUT15), .B(G87), .Z(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT66), .B(G20), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n272), .A2(new_n390), .B1(G77), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT8), .B(G58), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT77), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n210), .A2(new_n271), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n259), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT78), .B1(new_n337), .B2(new_n203), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n337), .A2(KEYINPUT78), .A3(new_n203), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(G77), .C2(new_n284), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n291), .A2(G238), .A3(G1698), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(new_n207), .B2(new_n291), .C1(new_n293), .C2(new_n241), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n306), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n309), .B1(new_n317), .B2(G244), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(G200), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n406), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT76), .B1(new_n408), .B2(G190), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT76), .ZN(new_n410));
  INV_X1    g0210(.A(G190), .ZN(new_n411));
  NOR3_X1   g0211(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n407), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G179), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n406), .A2(new_n371), .B1(new_n397), .B2(new_n400), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n383), .A2(new_n389), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n285), .B1(new_n289), .B2(new_n260), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n321), .A2(new_n322), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(G169), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT75), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n419), .B(new_n423), .C1(G169), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n414), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT12), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n337), .B2(new_n218), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n335), .A2(new_n218), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n272), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  OAI22_X1  g0232(.A1(new_n431), .A2(new_n432), .B1(new_n202), .B2(new_n395), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n260), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n430), .B1(new_n436), .B2(KEYINPUT11), .ZN(new_n437));
  INV_X1    g0237(.A(new_n435), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n259), .B1(new_n438), .B2(new_n433), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT11), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n308), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n312), .A2(KEYINPUT79), .A3(G274), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n317), .A2(G238), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n296), .A2(new_n298), .A3(G232), .A4(G1698), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n296), .A2(new_n298), .A3(G226), .A4(new_n292), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G97), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n306), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT13), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n446), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n371), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT14), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n453), .A2(new_n455), .ZN(new_n458));
  OAI22_X1  g0258(.A1(new_n456), .A2(new_n457), .B1(new_n458), .B2(new_n414), .ZN(new_n459));
  AOI211_X1 g0259(.A(KEYINPUT14), .B(new_n371), .C1(new_n453), .C2(new_n455), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n442), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(G190), .A3(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(G200), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n437), .A2(new_n441), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  AND4_X1   g0265(.A1(new_n333), .A2(new_n418), .A3(new_n426), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n337), .A2(new_n206), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n281), .A2(G33), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n260), .A2(new_n282), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(new_n206), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n345), .A2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n208), .A2(KEYINPUT83), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n475));
  AND2_X1   g0275(.A1(G97), .A2(G107), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G97), .A2(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n474), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n474), .A2(new_n478), .A3(KEYINPUT84), .A4(new_n479), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n391), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n274), .A2(G77), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n470), .B1(new_n486), .B2(new_n259), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n296), .A2(new_n298), .A3(G244), .A4(new_n292), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT85), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT86), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n299), .A2(new_n494), .A3(KEYINPUT4), .A4(G244), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n291), .A2(KEYINPUT4), .A3(G244), .A4(new_n292), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(G1698), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n306), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n281), .A2(G45), .ZN(new_n503));
  INV_X1    g0303(.A(G274), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g0305(.A(KEYINPUT5), .B(G41), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n503), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n316), .A2(new_n314), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G257), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n502), .A2(G190), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n487), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n500), .A2(new_n499), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(KEYINPUT86), .B2(new_n497), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n515), .A2(new_n493), .A3(new_n495), .A4(new_n491), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n513), .B1(new_n516), .B2(new_n306), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n384), .B1(new_n517), .B2(new_n507), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT87), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n502), .A2(new_n507), .A3(new_n510), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G200), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT87), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n487), .A4(new_n511), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n502), .A2(new_n414), .A3(new_n507), .A4(new_n510), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n484), .A2(new_n485), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n342), .B1(new_n291), .B2(G20), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n211), .A2(new_n213), .B1(new_n296), .B2(new_n298), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n526), .A2(new_n339), .B1(new_n527), .B2(KEYINPUT7), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n207), .B1(new_n528), .B2(new_n343), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n259), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n470), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n371), .A2(new_n520), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n519), .A2(new_n523), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n282), .A2(G116), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G116), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n469), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n271), .A2(G97), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n214), .A2(new_n499), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n536), .A2(G20), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n259), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n259), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(KEYINPUT20), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n505), .A2(new_n506), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n509), .B2(G270), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n296), .A2(new_n298), .A3(G257), .A4(new_n292), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n296), .A2(new_n298), .A3(G264), .A4(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(G303), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n291), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n306), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n371), .B1(new_n550), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n550), .A2(new_n555), .A3(G179), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n550), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n550), .A2(new_n555), .A3(G190), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n548), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n554), .A2(new_n306), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n566));
  INV_X1    g0366(.A(new_n215), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n316), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g0368(.A(KEYINPUT5), .B(G41), .Z(new_n569));
  OAI21_X1  g0369(.A(new_n568), .B1(new_n569), .B2(new_n503), .ZN(new_n570));
  INV_X1    g0370(.A(G270), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n507), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(G169), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT90), .B1(new_n548), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n537), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n259), .A2(new_n541), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT89), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n259), .A2(new_n540), .A3(new_n541), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT20), .B1(new_n579), .B2(new_n539), .ZN(new_n580));
  INV_X1    g0380(.A(new_n547), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT90), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n556), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT21), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n574), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT91), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n574), .A2(new_n584), .A3(KEYINPUT91), .A4(new_n585), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n559), .B(new_n564), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n296), .A2(new_n298), .A3(G250), .A4(new_n292), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n296), .A2(new_n298), .A3(G257), .A4(G1698), .ZN(new_n592));
  NAND2_X1  g0392(.A1(G33), .A2(G294), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n306), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n509), .A2(G264), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(G179), .A4(new_n507), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT92), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n596), .A3(new_n507), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n597), .A2(new_n598), .B1(new_n599), .B2(G169), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n597), .A2(new_n598), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n469), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT25), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n282), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n603), .A2(G107), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(KEYINPUT23), .B1(new_n210), .B2(G107), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G116), .ZN(new_n609));
  OR2_X1    g0409(.A1(KEYINPUT23), .A2(G107), .ZN(new_n610));
  OAI221_X1 g0410(.A(new_n608), .B1(G20), .B2(new_n609), .C1(new_n214), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n214), .A2(new_n291), .A3(G87), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT22), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT22), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n214), .A2(new_n291), .A3(new_n614), .A4(G87), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n259), .B1(new_n616), .B2(KEYINPUT24), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT24), .ZN(new_n618));
  AOI211_X1 g0418(.A(new_n618), .B(new_n611), .C1(new_n613), .C2(new_n615), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n607), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n602), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n599), .A2(G200), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n411), .B2(new_n599), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n391), .A2(new_n625), .B1(G87), .B2(new_n208), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n214), .A2(new_n291), .A3(G68), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT19), .B1(new_n272), .B2(G97), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n259), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n390), .A2(new_n282), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n603), .A2(G87), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n508), .B1(new_n314), .B2(new_n316), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n505), .B1(new_n635), .B2(G250), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n296), .A2(new_n298), .A3(G244), .A4(G1698), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n296), .A2(new_n298), .A3(G238), .A4(new_n292), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n609), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n306), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n636), .A2(new_n640), .A3(KEYINPUT88), .A4(G190), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n640), .A3(G190), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT88), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n636), .A2(new_n640), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n634), .A2(new_n641), .A3(new_n644), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n603), .A2(new_n390), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n630), .A2(new_n648), .A3(new_n632), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n645), .A2(new_n371), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n636), .A2(new_n640), .A3(new_n414), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n621), .A2(new_n624), .A3(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n466), .A2(new_n533), .A3(new_n590), .A4(new_n654), .ZN(G372));
  NAND2_X1  g0455(.A1(new_n520), .A2(new_n371), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n530), .A2(new_n531), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n524), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT26), .B1(new_n658), .B2(new_n653), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n391), .A2(new_n271), .A3(new_n206), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n627), .B(new_n626), .C1(new_n660), .C2(KEYINPUT19), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n631), .B1(new_n661), .B2(new_n259), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n646), .A2(new_n662), .A3(new_n642), .A4(new_n633), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n652), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n532), .A2(new_n665), .A3(new_n666), .A4(new_n524), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n659), .A2(new_n652), .A3(new_n667), .ZN(new_n668));
  AOI211_X1 g0468(.A(new_n559), .B(new_n621), .C1(new_n588), .C2(new_n589), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n519), .A2(new_n523), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n652), .B(new_n663), .C1(new_n620), .C2(new_n623), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n670), .A2(new_n658), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n668), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n466), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT93), .Z(new_n676));
  INV_X1    g0476(.A(new_n426), .ZN(new_n677));
  INV_X1    g0477(.A(new_n461), .ZN(new_n678));
  INV_X1    g0478(.A(new_n417), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n464), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n389), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  AOI211_X1 g0482(.A(new_n376), .B(new_n373), .C1(new_n380), .C2(new_n338), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT18), .B1(new_n363), .B2(new_n374), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n377), .A2(KEYINPUT94), .A3(new_n382), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n677), .B1(new_n688), .B2(new_n333), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n676), .A2(new_n689), .ZN(G369));
  INV_X1    g0490(.A(G13), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n391), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n281), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n214), .A2(new_n281), .A3(G13), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n694), .A2(new_n696), .A3(G213), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G343), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT95), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n548), .ZN(new_n701));
  INV_X1    g0501(.A(new_n559), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n582), .A2(new_n556), .ZN(new_n703));
  AOI21_X1  g0503(.A(KEYINPUT21), .B1(new_n703), .B2(KEYINPUT90), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT91), .B1(new_n704), .B2(new_n584), .ZN(new_n705));
  INV_X1    g0505(.A(new_n589), .ZN(new_n706));
  OAI211_X1 g0506(.A(new_n702), .B(new_n563), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n701), .B1(new_n707), .B2(KEYINPUT96), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n590), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n708), .A2(new_n710), .B1(new_n711), .B2(new_n701), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n699), .A2(new_n620), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n602), .A2(new_n620), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n715), .B(new_n716), .C1(new_n620), .C2(new_n623), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n621), .A2(new_n699), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n716), .A2(new_n699), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT97), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n711), .A2(new_n722), .A3(new_n700), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n559), .B1(new_n588), .B2(new_n589), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT97), .B1(new_n724), .B2(new_n699), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n720), .A2(new_n727), .ZN(G399));
  NOR2_X1   g0528(.A1(new_n226), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G1), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n732), .B1(new_n220), .B2(new_n730), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  XNOR2_X1  g0534(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n659), .A2(new_n652), .A3(new_n667), .ZN(new_n736));
  AOI221_X4 g0536(.A(new_n671), .B1(new_n532), .B2(new_n524), .C1(new_n519), .C2(new_n523), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n702), .B(new_n716), .C1(new_n705), .C2(new_n706), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n735), .B1(new_n739), .B2(new_n699), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(new_n533), .A3(new_n672), .ZN(new_n741));
  INV_X1    g0541(.A(new_n653), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n532), .A3(new_n666), .A4(new_n524), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT26), .B1(new_n658), .B2(new_n664), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n743), .A2(new_n744), .A3(new_n652), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT29), .A3(new_n700), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n740), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n599), .A2(new_n414), .A3(new_n645), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n520), .A2(new_n560), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT98), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n558), .A2(new_n599), .A3(new_n645), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n517), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n599), .A2(new_n645), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n550), .A2(G179), .A3(new_n555), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n502), .A3(new_n757), .A4(new_n510), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(KEYINPUT30), .ZN(new_n760));
  OAI211_X1 g0560(.A(KEYINPUT31), .B(new_n699), .C1(new_n755), .C2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n759), .A2(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(new_n754), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n750), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT31), .B1(new_n765), .B2(new_n699), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n590), .A2(new_n533), .A3(new_n654), .A4(new_n700), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n713), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n748), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n734), .B1(new_n770), .B2(G1), .ZN(G364));
  AOI21_X1  g0571(.A(new_n281), .B1(new_n692), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n729), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n714), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n708), .A2(new_n710), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n711), .A2(new_n701), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G330), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n712), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n411), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n214), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n303), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n391), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n789), .B1(G329), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n214), .A2(new_n414), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n795), .A2(new_n411), .A3(G200), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G322), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n414), .A2(G200), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT102), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(new_n411), .A3(new_n391), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n793), .B(new_n797), .C1(new_n798), .C2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n794), .A2(new_n411), .A3(new_n384), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n800), .A2(G20), .A3(G190), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT103), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n802), .B(new_n809), .C1(G303), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT101), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n795), .B2(new_n384), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n794), .A2(KEYINPUT101), .A3(G200), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n817), .A2(G190), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n817), .A2(new_n411), .A3(new_n818), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT33), .B(G317), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G326), .A2(new_n820), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n814), .A2(G87), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n792), .A2(G159), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT32), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G58), .B2(new_n796), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n801), .A2(new_n207), .ZN(new_n829));
  INV_X1    g0629(.A(new_n787), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n303), .B(new_n829), .C1(G97), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n806), .A2(G77), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n825), .A2(new_n828), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G50), .A2(new_n820), .B1(new_n822), .B2(G68), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n815), .A2(new_n824), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n215), .B1(G20), .B2(new_n371), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n783), .A2(new_n837), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n226), .A2(new_n303), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n841), .A2(G355), .B1(new_n536), .B2(new_n226), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n226), .A2(new_n291), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(G45), .B2(new_n220), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n252), .A2(new_n311), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n785), .B(new_n839), .C1(new_n840), .C2(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n775), .A2(new_n780), .B1(new_n784), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  NOR2_X1   g0649(.A1(new_n417), .A2(new_n699), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n699), .A2(new_n401), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n413), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n850), .B1(new_n852), .B2(new_n417), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n739), .B2(new_n699), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n674), .A2(new_n700), .A3(new_n853), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n769), .A3(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT106), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n769), .B1(new_n855), .B2(new_n856), .ZN(new_n860));
  NOR3_X1   g0660(.A1(new_n859), .A2(new_n774), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n858), .B2(new_n857), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n837), .A2(new_n781), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n774), .B1(G77), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT104), .Z(new_n866));
  AOI22_X1  g0666(.A1(new_n806), .A2(G159), .B1(G143), .B2(new_n796), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  INV_X1    g0668(.A(G150), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n819), .C1(new_n869), .C2(new_n821), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT34), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n801), .A2(new_n218), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n291), .B1(new_n791), .B2(new_n873), .C1(new_n787), .C2(new_n217), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n872), .B(new_n874), .C1(new_n814), .C2(G50), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n819), .A2(new_n553), .ZN(new_n876));
  INV_X1    g0676(.A(new_n801), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(G87), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n830), .A2(G97), .B1(new_n792), .B2(G311), .ZN(new_n879));
  INV_X1    g0679(.A(new_n796), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n878), .B(new_n879), .C1(new_n788), .C2(new_n880), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n876), .B(new_n881), .C1(G116), .C2(new_n806), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n822), .A2(G283), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n291), .B1(new_n814), .B2(G107), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT105), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n871), .A2(new_n875), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n866), .B1(new_n782), .B2(new_n853), .C1(new_n887), .C2(new_n838), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n862), .A2(new_n888), .ZN(G384));
  NAND2_X1  g0689(.A1(new_n482), .A2(new_n483), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT35), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n482), .A2(KEYINPUT35), .A3(new_n483), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n216), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  NAND3_X1  g0695(.A1(new_n221), .A2(G77), .A3(new_n348), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n202), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n281), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT108), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT37), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT16), .B1(new_n356), .B2(new_n360), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n338), .B1(new_n362), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n374), .B2(new_n697), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n901), .B1(new_n904), .B2(new_n388), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n363), .A2(new_n697), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n375), .A2(new_n907), .A3(new_n901), .A4(new_n388), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT107), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n903), .A2(new_n697), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n389), .B2(new_n383), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n380), .A2(new_n387), .A3(new_n338), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n381), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(KEYINPUT107), .A3(new_n901), .A4(new_n907), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n908), .A2(new_n909), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n905), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n921), .A2(new_n922), .A3(new_n914), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n900), .B1(new_n916), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n915), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n922), .B1(new_n921), .B2(new_n914), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT108), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n442), .A2(new_n699), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n461), .A2(new_n464), .A3(new_n928), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n442), .B(new_n699), .C1(new_n459), .C2(new_n460), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n853), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n767), .B2(new_n768), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n924), .A2(new_n927), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n907), .B1(new_n687), .B2(new_n389), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n901), .B1(new_n918), .B2(new_n907), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n920), .B2(new_n919), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n922), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n935), .B1(new_n940), .B2(new_n925), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n933), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n936), .A2(G330), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n466), .A2(new_n769), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n934), .A2(new_n935), .B1(new_n933), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n767), .A2(new_n768), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n466), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n740), .A2(new_n747), .A3(new_n466), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n689), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n949), .B(new_n951), .Z(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT39), .B1(new_n916), .B2(new_n923), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT39), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n940), .A2(new_n954), .A3(new_n925), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n678), .A2(new_n700), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT109), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n931), .ZN(new_n961));
  INV_X1    g0761(.A(new_n850), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(new_n856), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n963), .A2(new_n924), .A3(new_n927), .ZN(new_n964));
  INV_X1    g0764(.A(new_n697), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n685), .A2(new_n686), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n960), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n952), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n281), .B2(new_n692), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n952), .A2(new_n968), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n899), .B1(new_n970), .B2(new_n971), .ZN(G367));
  AOI21_X1  g0772(.A(new_n291), .B1(new_n792), .B2(G317), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n207), .B2(new_n787), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n880), .A2(new_n553), .B1(new_n206), .B2(new_n801), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(G283), .C2(new_n806), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n976), .B1(new_n788), .B2(new_n821), .C1(new_n808), .C2(new_n819), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n814), .A2(G116), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT46), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n806), .A2(G50), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n877), .A2(G77), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n291), .ZN(new_n982));
  INV_X1    g0782(.A(new_n814), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n980), .B1(KEYINPUT111), .B2(new_n982), .C1(new_n983), .C2(new_n217), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n787), .A2(new_n218), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G137), .B2(new_n792), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n880), .B2(new_n869), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(KEYINPUT111), .B2(new_n982), .ZN(new_n988));
  INV_X1    g0788(.A(G143), .ZN(new_n989));
  INV_X1    g0789(.A(G159), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n988), .B1(new_n989), .B2(new_n819), .C1(new_n990), .C2(new_n821), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n977), .A2(new_n979), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT47), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n838), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n993), .B2(new_n992), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n248), .A2(new_n843), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n783), .B(new_n837), .C1(new_n226), .C2(new_n390), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n785), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n783), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n700), .A2(new_n634), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n665), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n652), .B2(new_n1000), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n995), .B(new_n998), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n719), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n712), .B2(new_n713), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n720), .A2(new_n726), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n726), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n719), .B1(new_n778), .B2(G330), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n712), .A2(new_n713), .A3(new_n1004), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n726), .A2(new_n719), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n721), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n658), .A2(new_n700), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n699), .A2(new_n657), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n533), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1004), .B1(new_n723), .B2(new_n725), .ZN(new_n1019));
  OAI211_X1 g0819(.A(KEYINPUT44), .B(new_n1017), .C1(new_n1019), .C2(new_n721), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1017), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT45), .B1(new_n727), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT45), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1019), .A2(new_n1024), .A3(new_n721), .A4(new_n1017), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1018), .A2(new_n1021), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n1009), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n720), .B1(new_n1023), .B2(new_n1025), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1011), .A2(new_n1027), .A3(new_n770), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n770), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n729), .B(KEYINPUT41), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n773), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n533), .A2(new_n621), .A3(new_n1016), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n699), .B1(new_n1033), .B2(new_n658), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(new_n1035), .B2(KEYINPUT42), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(KEYINPUT42), .B2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OR3_X1    g0839(.A1(new_n720), .A2(KEYINPUT110), .A3(new_n1017), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1002), .A2(KEYINPUT43), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT110), .B1(new_n720), .B2(new_n1017), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1041), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1039), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n1043), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1003), .B1(new_n1032), .B2(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n244), .A2(G45), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n731), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1054), .A2(new_n843), .B1(new_n1055), .B2(new_n841), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n1055), .C1(G68), .C2(G77), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n394), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n202), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1057), .B1(new_n1059), .B2(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT50), .B2(new_n1059), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n1056), .A2(new_n1061), .B1(G107), .B2(new_n225), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n785), .B1(new_n1062), .B2(new_n840), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n719), .B2(new_n999), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n390), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n291), .B1(new_n791), .B2(new_n869), .C1(new_n787), .C2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n880), .A2(new_n202), .B1(new_n206), .B2(new_n801), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(G68), .C2(new_n806), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n814), .A2(G77), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n820), .A2(G159), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n822), .A2(new_n334), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n806), .A2(G303), .B1(G317), .B2(new_n796), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n820), .A2(G322), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(new_n808), .C2(new_n821), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT48), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n798), .B2(new_n787), .C1(new_n788), .C2(new_n983), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1078));
  XOR2_X1   g0878(.A(new_n1077), .B(new_n1078), .Z(new_n1079));
  AOI21_X1  g0879(.A(new_n291), .B1(new_n792), .B2(G326), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n536), .B2(new_n801), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1072), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1064), .B1(new_n1082), .B2(new_n837), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1011), .B2(new_n773), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1011), .A2(new_n770), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT113), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n770), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n729), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1087), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1084), .B1(new_n1090), .B2(new_n1091), .ZN(G393));
  INV_X1    g0892(.A(KEYINPUT114), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1027), .A2(new_n1093), .A3(new_n1028), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1026), .A2(KEYINPUT114), .A3(new_n1009), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n1085), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n729), .A3(new_n1029), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n787), .A2(new_n203), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n291), .B1(new_n791), .B2(new_n989), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n877), .C2(G87), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n394), .B2(new_n807), .C1(new_n983), .C2(new_n218), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n819), .A2(new_n869), .B1(new_n880), .B2(new_n990), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  AOI211_X1 g0903(.A(new_n1101), .B(new_n1103), .C1(G50), .C2(new_n822), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n303), .B1(new_n787), .B2(new_n536), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(G322), .B2(new_n792), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n207), .B2(new_n801), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n814), .B2(G283), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1108), .B1(new_n788), .B2(new_n807), .C1(new_n553), .C2(new_n821), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n820), .A2(G317), .B1(G311), .B2(new_n796), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n837), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n255), .A2(new_n226), .A3(new_n291), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n840), .B1(new_n225), .B2(new_n206), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1114), .B(new_n774), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n783), .B2(new_n1017), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n773), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1120), .ZN(G390));
  NOR2_X1   g0921(.A1(new_n956), .A2(new_n782), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n814), .A2(G150), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT53), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n291), .B1(new_n791), .B2(new_n1125), .C1(new_n787), .C2(new_n990), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n880), .A2(new_n873), .B1(new_n202), .B2(new_n801), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(KEYINPUT54), .B(G143), .Z(new_n1129));
  AOI22_X1  g0929(.A1(new_n822), .A2(G137), .B1(new_n806), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT116), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1130), .A2(KEYINPUT116), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1123), .A2(KEYINPUT53), .B1(G128), .B2(new_n820), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n822), .A2(G107), .B1(new_n806), .B2(G97), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT117), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n291), .B(new_n1098), .C1(G294), .C2(new_n792), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n872), .B1(G116), .B2(new_n796), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n825), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(new_n798), .C2(new_n819), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1134), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT118), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n838), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n774), .B1(new_n334), .B2(new_n864), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1122), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n940), .A2(new_n925), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n699), .B1(new_n741), .B2(new_n745), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n852), .A2(new_n417), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n850), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n958), .B(new_n1150), .C1(new_n1153), .C2(new_n961), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n947), .A2(G330), .A3(new_n853), .A4(new_n931), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n856), .A2(new_n962), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n959), .B1(new_n1156), .B2(new_n931), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1154), .B(new_n1155), .C1(new_n1157), .C2(new_n956), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n953), .B(new_n955), .C1(new_n963), .C2(new_n959), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1155), .B1(new_n1160), .B2(new_n1154), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1149), .B1(new_n1162), .B2(new_n773), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n931), .B1(new_n769), .B2(new_n853), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n713), .B(new_n932), .C1(new_n768), .C2(new_n767), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n713), .B(new_n854), .C1(new_n767), .C2(new_n768), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1155), .B(new_n1153), .C1(new_n1167), .C2(new_n931), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n950), .A2(new_n689), .A3(new_n944), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT115), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT115), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n950), .A2(new_n1172), .A3(new_n689), .A4(new_n944), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n729), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1154), .B1(new_n1157), .B2(new_n956), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1165), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1158), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(new_n1174), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1163), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT119), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT119), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1163), .B(new_n1183), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1182), .A2(new_n1184), .ZN(G378));
  AND2_X1   g0985(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1169), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1186), .B1(new_n1179), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n419), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(new_n965), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n333), .A2(new_n426), .A3(KEYINPUT55), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT55), .B1(new_n333), .B2(new_n426), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n333), .A2(new_n426), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT55), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1190), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n333), .A2(new_n426), .A3(KEYINPUT55), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1193), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n943), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n946), .A2(new_n1205), .A3(G330), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1204), .A2(new_n968), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n968), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1208));
  OAI211_X1 g1008(.A(KEYINPUT57), .B(new_n1188), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n943), .A2(new_n1203), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1205), .B1(new_n946), .B2(G330), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n967), .A2(KEYINPUT124), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1204), .A2(new_n1214), .A3(new_n1206), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1186), .A2(new_n1178), .A3(new_n1158), .A4(new_n1169), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1213), .A2(new_n1215), .B1(new_n1186), .B2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1209), .B(new_n729), .C1(new_n1217), .C2(KEYINPUT57), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1204), .A2(new_n1214), .A3(new_n1206), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1214), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n773), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1203), .A2(new_n781), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n291), .A2(G41), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G50), .B(new_n1223), .C1(new_n271), .C2(new_n310), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1223), .B1(new_n791), .B2(new_n798), .C1(new_n787), .C2(new_n218), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n880), .A2(new_n207), .B1(new_n217), .B2(new_n801), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n814), .C2(G77), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n807), .A2(new_n1065), .B1(new_n206), .B2(new_n821), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT120), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1227), .B1(new_n536), .B2(new_n819), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT58), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1224), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n796), .A2(G128), .B1(new_n830), .B2(G150), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n807), .B2(new_n868), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G125), .B2(new_n820), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n814), .A2(new_n1129), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1238), .A2(KEYINPUT121), .B1(G132), .B2(new_n822), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1237), .B(new_n1239), .C1(KEYINPUT121), .C2(new_n1238), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n990), .C2(new_n801), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1234), .B1(new_n1233), .B2(new_n1232), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n837), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT122), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n863), .A2(new_n202), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1222), .A2(new_n774), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1221), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1218), .A2(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n961), .A2(new_n781), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n864), .A2(G68), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n291), .B1(new_n787), .B2(new_n202), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n880), .A2(new_n868), .B1(new_n217), .B2(new_n801), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1255), .B(new_n1256), .C1(G128), .C2(new_n792), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n869), .B2(new_n807), .C1(new_n983), .C2(new_n990), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1129), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n873), .A2(new_n819), .B1(new_n821), .B2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n806), .A2(G107), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT125), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n981), .A2(new_n303), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .C1(new_n983), .C2(new_n206), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n787), .A2(new_n1065), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n791), .A2(new_n553), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n880), .B2(new_n798), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(new_n1263), .B2(new_n1262), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n1269), .B1(new_n536), .B2(new_n821), .C1(new_n788), .C2(new_n819), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1258), .A2(new_n1260), .B1(new_n1264), .B2(new_n1270), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n785), .B(new_n1254), .C1(new_n1271), .C2(new_n837), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1169), .A2(new_n773), .B1(new_n1253), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1174), .A2(new_n1031), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1169), .B1(new_n1173), .B2(new_n1171), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(G381));
  OAI21_X1  g1076(.A(new_n1188), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT57), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n967), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1204), .A2(new_n968), .A3(new_n1206), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1216), .B2(new_n1186), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n730), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1250), .B1(new_n1279), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n848), .B(new_n1084), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1286));
  NOR4_X1   g1086(.A1(G390), .A2(G384), .A3(new_n1286), .A4(G381), .ZN(new_n1287));
  INV_X1    g1087(.A(G387), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1181), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1285), .A2(new_n1287), .A3(new_n1288), .A4(new_n1289), .ZN(G407));
  NAND2_X1  g1090(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G343), .C2(new_n1291), .ZN(G409));
  AND2_X1   g1092(.A1(new_n1097), .A2(new_n1120), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT127), .B1(G387), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1286), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(G387), .A2(new_n1293), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1031), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(new_n1029), .B2(new_n770), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1051), .B(new_n1046), .C1(new_n1299), .C2(new_n773), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G390), .B1(new_n1003), .B2(new_n1300), .ZN(new_n1301));
  OAI22_X1  g1101(.A1(new_n1294), .A2(new_n1296), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1293), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1296), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1300), .A2(G390), .A3(new_n1003), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT127), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1302), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n1186), .B2(new_n1169), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1275), .A2(KEYINPUT60), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1309), .A2(new_n1310), .A3(new_n729), .A4(new_n1174), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1311), .A2(G384), .A3(new_n1273), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1311), .B2(new_n1273), .ZN(new_n1314));
  INV_X1    g1114(.A(G213), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1315), .A2(G343), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G2897), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1313), .A2(new_n1314), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1311), .A2(new_n1273), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1317), .B1(new_n1322), .B2(new_n1312), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1249), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1325), .B1(new_n1282), .B2(new_n773), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1031), .B(new_n1188), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1181), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1285), .B2(G378), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1324), .B1(new_n1329), .B2(new_n1316), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1312), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(G378), .A2(new_n1218), .A3(new_n1251), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1289), .ZN(new_n1335));
  AOI211_X1 g1135(.A(new_n1316), .B(new_n1332), .C1(new_n1333), .C2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  OAI211_X1 g1137(.A(new_n1330), .B(new_n1331), .C1(new_n1336), .C2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1316), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1322), .A4(new_n1312), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1341), .A2(KEYINPUT62), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1307), .B1(new_n1338), .B2(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1318), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1322), .A2(new_n1312), .A3(new_n1317), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1346), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1347), .A2(new_n1307), .A3(KEYINPUT61), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT126), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT63), .B1(new_n1336), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT63), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1341), .A2(KEYINPUT126), .A3(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1348), .A2(new_n1350), .A3(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1343), .A2(new_n1353), .ZN(G405));
  NAND2_X1  g1154(.A1(G375), .A2(new_n1289), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1355), .A2(new_n1333), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1332), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1356), .A2(new_n1332), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1307), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  OR2_X1    g1160(.A1(new_n1356), .A2(new_n1332), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1361), .A2(new_n1306), .A3(new_n1302), .A4(new_n1357), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1360), .A2(new_n1362), .ZN(G402));
endmodule


