//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1174, new_n1175, new_n1176,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1259, new_n1260;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT64), .B(G244), .Z(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT65), .Z(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n204), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n220), .B(new_n228), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n217), .A2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G274), .ZN(new_n247));
  AND2_X1   g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  AOI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n248), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n251), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n255), .B2(new_n234), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G223), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n258), .B1(new_n259), .B2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT74), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G33), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n260), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G87), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n257), .B(KEYINPUT77), .C1(new_n270), .C2(new_n254), .ZN(new_n271));
  INV_X1    g0071(.A(G200), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT77), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n254), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n271), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n257), .B1(new_n270), .B2(new_n254), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(G190), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n205), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n226), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT16), .ZN(new_n281));
  AOI21_X1  g0081(.A(G33), .B1(new_n263), .B2(new_n264), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n262), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(KEYINPUT7), .B(new_n204), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT7), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT3), .B(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G20), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n222), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G58), .A2(G68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT75), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(new_n223), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G20), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G159), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n281), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(G20), .B1(new_n265), .B2(new_n267), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n286), .ZN(new_n301));
  OAI21_X1  g0101(.A(G68), .B1(new_n300), .B2(new_n286), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT76), .ZN(new_n303));
  AND3_X1   g0103(.A1(new_n295), .A2(new_n303), .A3(new_n297), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n303), .B1(new_n295), .B2(new_n297), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n301), .A2(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n280), .B(new_n299), .C1(new_n306), .C2(new_n281), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n308), .A2(new_n204), .A3(G1), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n280), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n203), .A2(G20), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n310), .A2(new_n314), .B1(new_n311), .B2(new_n309), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n278), .A2(new_n307), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT17), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n316), .B(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n277), .A2(G179), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n271), .A2(new_n320), .A3(new_n275), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n307), .A2(new_n315), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n234), .A2(G1698), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n287), .B(new_n331), .C1(G226), .C2(G1698), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G238), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n253), .B1(new_n255), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n254), .B1(new_n332), .B2(new_n333), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT13), .B1(new_n342), .B2(new_n338), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n344), .A2(new_n345), .A3(G169), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n320), .B1(new_n341), .B2(new_n343), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n345), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n349), .A2(new_n345), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NOR4_X1   g0155(.A1(new_n280), .A2(new_n222), .A3(new_n309), .A4(new_n313), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT72), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n204), .A2(G33), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G77), .B1(G20), .B2(new_n222), .ZN(new_n360));
  INV_X1    g0160(.A(G50), .ZN(new_n361));
  INV_X1    g0161(.A(new_n296), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n363), .A2(new_n280), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n364), .A2(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(KEYINPUT11), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n309), .A2(new_n222), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT12), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n357), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n355), .A2(new_n369), .ZN(new_n370));
  AND4_X1   g0170(.A1(new_n357), .A2(new_n365), .A3(new_n366), .A4(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n344), .A2(G200), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n344), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n330), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n287), .A2(G222), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT66), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n267), .A2(new_n283), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n376), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G223), .B1(G77), .B2(new_n380), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT67), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n254), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n379), .A2(KEYINPUT67), .A3(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n253), .B1(new_n255), .B2(new_n259), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT69), .B1(new_n390), .B2(G179), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n248), .B1(new_n205), .B2(G33), .ZN(new_n392));
  INV_X1    g0192(.A(new_n311), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n359), .B1(G150), .B2(new_n296), .ZN(new_n394));
  NOR2_X1   g0194(.A1(G50), .A2(G58), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n204), .B1(new_n395), .B2(new_n222), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n392), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n309), .A2(new_n361), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n312), .A2(G50), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT68), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n310), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n400), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT69), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n352), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n390), .A2(new_n320), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n391), .A2(new_n404), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n310), .A2(G77), .A3(new_n312), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n410), .B(KEYINPUT70), .ZN(new_n411));
  XNOR2_X1  g0211(.A(KEYINPUT15), .B(G87), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n359), .B1(G20), .B2(G77), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n362), .B2(new_n311), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n280), .B1(new_n208), .B2(new_n309), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n253), .B1(new_n255), .B2(new_n207), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n381), .A2(G238), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n287), .A2(G232), .A3(new_n376), .ZN(new_n420));
  INV_X1    g0220(.A(G107), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(new_n287), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n422), .B2(new_n335), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n352), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n417), .B(new_n424), .C1(G169), .C2(new_n423), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n423), .A2(G190), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(new_n411), .A3(new_n416), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(new_n272), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT10), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n404), .A2(KEYINPUT9), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n403), .A2(new_n400), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n434), .A2(KEYINPUT9), .A3(new_n398), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n390), .A2(G200), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  AOI211_X1 g0236(.A(new_n373), .B(new_n388), .C1(new_n385), .C2(new_n386), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n432), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n435), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n405), .B2(new_n272), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n441), .A2(KEYINPUT10), .A3(new_n437), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n409), .B(new_n431), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(KEYINPUT71), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n375), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n309), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n203), .A2(G33), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n392), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(KEYINPUT25), .B1(new_n309), .B2(new_n421), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n309), .A2(KEYINPUT25), .A3(new_n421), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n449), .A2(G107), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT85), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n265), .A2(new_n204), .A3(G87), .A4(new_n267), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT84), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT22), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n456), .B2(KEYINPUT22), .ZN(new_n459));
  INV_X1    g0259(.A(G87), .ZN(new_n460));
  NOR4_X1   g0260(.A1(new_n380), .A2(KEYINPUT22), .A3(G20), .A4(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n204), .B2(G107), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n421), .A2(KEYINPUT23), .A3(G20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT81), .A2(G116), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT81), .A2(G116), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G33), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n471), .B2(G20), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n455), .B1(new_n462), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n456), .A2(KEYINPUT22), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT22), .ZN(new_n476));
  INV_X1    g0276(.A(new_n461), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n472), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(KEYINPUT85), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT85), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n392), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n454), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n265), .A2(new_n267), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n376), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G257), .B2(new_n376), .ZN(new_n489));
  INV_X1    g0289(.A(G294), .ZN(new_n490));
  OAI22_X1  g0290(.A1(new_n486), .A2(new_n489), .B1(new_n266), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n335), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT78), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(G41), .ZN(new_n495));
  INV_X1    g0295(.A(G41), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n203), .A2(G45), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n498), .A2(new_n501), .A3(new_n250), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT79), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n498), .A2(new_n501), .A3(new_n250), .A4(KEYINPUT79), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n498), .A2(new_n501), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n507), .A2(G264), .A3(new_n254), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n492), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n335), .B1(new_n498), .B2(new_n501), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT86), .A3(G264), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n492), .A2(new_n506), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(G169), .A2(new_n510), .B1(new_n516), .B2(G179), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n485), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n373), .A2(new_n509), .B1(new_n515), .B2(new_n272), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n454), .B(new_n519), .C1(new_n481), .C2(new_n484), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n470), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n449), .A2(G116), .B1(new_n309), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(G20), .B1(new_n266), .B2(G97), .ZN(new_n524));
  INV_X1    g0324(.A(G283), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n266), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n280), .B(new_n526), .C1(new_n204), .C2(new_n470), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(G257), .A2(G1698), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G264), .B2(new_n376), .ZN(new_n533));
  INV_X1    g0333(.A(G303), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n486), .A2(new_n533), .B1(new_n534), .B2(new_n287), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n335), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n513), .A2(G270), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n506), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(G200), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n373), .B2(new_n538), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT83), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT21), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n531), .A2(G169), .A3(new_n543), .A4(new_n538), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n531), .A2(G169), .A3(new_n538), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n541), .A3(new_n542), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n536), .A2(new_n506), .A3(G179), .A4(new_n537), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n531), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n540), .A2(new_n544), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n265), .A2(new_n204), .A3(G68), .A4(new_n267), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n333), .B2(new_n204), .ZN(new_n553));
  INV_X1    g0353(.A(G97), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n460), .A2(new_n554), .A3(new_n421), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n553), .A2(new_n555), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n551), .A2(new_n560), .A3(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n280), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n449), .A2(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n412), .A2(new_n309), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(G244), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n265), .A3(new_n267), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n254), .B1(new_n569), .B2(new_n471), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n500), .A2(new_n487), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n203), .A2(new_n247), .A3(G45), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n254), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G190), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n570), .B2(new_n574), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n449), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n562), .B(new_n564), .C1(new_n412), .C2(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n569), .A2(new_n471), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n352), .B(new_n573), .C1(new_n581), .C2(new_n254), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n320), .B1(new_n570), .B2(new_n574), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n565), .A2(new_n578), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n513), .A2(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT80), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n513), .A2(new_n588), .A3(G257), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n265), .A2(new_n267), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT4), .B1(new_n591), .B2(G244), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n567), .A3(G1698), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n287), .A2(new_n594), .B1(G33), .B2(G283), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n287), .B2(G250), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n376), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n335), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n590), .A2(new_n598), .A3(new_n506), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n320), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n285), .A2(new_n288), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G107), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n421), .A2(KEYINPUT6), .A3(G97), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n554), .A2(new_n421), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G97), .A2(G107), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(KEYINPUT6), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n280), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n447), .A2(G97), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n449), .B2(G97), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n590), .A2(new_n598), .A3(new_n352), .A4(new_n506), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n600), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n612), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n609), .B2(new_n280), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n590), .A2(new_n598), .A3(G190), .A4(new_n506), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n590), .A2(new_n598), .A3(new_n506), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n272), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n585), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n550), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n446), .A2(new_n521), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(G372));
  OAI21_X1  g0424(.A(KEYINPUT87), .B1(new_n520), .B2(new_n621), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n481), .A2(new_n484), .ZN(new_n626));
  INV_X1    g0426(.A(new_n519), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n453), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n615), .A2(new_n620), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT87), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .A4(new_n585), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n546), .A2(new_n544), .A3(new_n549), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n517), .B2(new_n485), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n625), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT88), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n625), .A2(new_n631), .A3(new_n633), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n578), .A2(new_n565), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n580), .A2(new_n584), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n640), .A2(new_n615), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n640), .B2(new_n615), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n639), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n635), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n446), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n409), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT89), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n650), .B1(new_n439), .B2(new_n442), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n436), .A2(new_n432), .A3(new_n438), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT10), .B1(new_n441), .B2(new_n437), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n369), .A2(new_n355), .B1(new_n426), .B2(new_n374), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n326), .B(new_n328), .C1(new_n656), .C2(new_n318), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n648), .A2(new_n658), .ZN(G369));
  NAND3_X1  g0459(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT27), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(new_n662), .A3(G213), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT90), .Z(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n521), .B1(new_n485), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n518), .A2(new_n667), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n531), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n632), .A2(new_n540), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n632), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n632), .A2(new_n667), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n521), .A2(new_n679), .B1(new_n518), .B2(new_n668), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(G399));
  NAND3_X1  g0481(.A1(new_n218), .A2(KEYINPUT91), .A3(new_n496), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT91), .B1(new_n218), .B2(new_n496), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n555), .A2(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n224), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n633), .A2(new_n628), .A3(new_n638), .A4(new_n629), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n667), .B1(new_n646), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n645), .B1(new_n634), .B2(KEYINPUT88), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n667), .B1(new_n694), .B2(new_n637), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n695), .B2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g0496(.A(new_n575), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n492), .A2(new_n512), .A3(new_n514), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n619), .A2(new_n548), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n619), .A2(KEYINPUT30), .A3(new_n548), .A4(new_n699), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n575), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n599), .A2(new_n515), .A3(new_n538), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT31), .B1(new_n706), .B2(new_n667), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n521), .A2(new_n622), .A3(new_n668), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n696), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n690), .B1(new_n716), .B2(G1), .ZN(new_n717));
  XOR2_X1   g0517(.A(new_n717), .B(KEYINPUT92), .Z(G364));
  AOI21_X1  g0518(.A(new_n226), .B1(G20), .B2(new_n320), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n204), .A2(G190), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G179), .A2(G200), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G159), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT32), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n204), .A2(new_n352), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(G190), .A3(G200), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n725), .A2(new_n726), .B1(new_n361), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n726), .B2(new_n725), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n204), .A2(new_n373), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n272), .A2(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n287), .B1(new_n733), .B2(new_n460), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n727), .A2(new_n373), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n734), .B1(G68), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n204), .B1(new_n722), .B2(G190), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT93), .Z(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G97), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n352), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n731), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n721), .A2(new_n732), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n221), .B1(new_n743), .B2(new_n421), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n741), .A2(new_n721), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n744), .B1(G77), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n730), .A2(new_n737), .A3(new_n740), .A4(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G322), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n380), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n728), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n750), .B1(G326), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n743), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G283), .A2(new_n753), .B1(new_n746), .B2(G311), .ZN(new_n754));
  INV_X1    g0554(.A(new_n733), .ZN(new_n755));
  INV_X1    g0555(.A(new_n723), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G303), .A2(new_n755), .B1(new_n756), .B2(G329), .ZN(new_n757));
  XNOR2_X1  g0557(.A(KEYINPUT33), .B(G317), .ZN(new_n758));
  INV_X1    g0558(.A(new_n738), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n736), .A2(new_n758), .B1(new_n759), .B2(G294), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n752), .A2(new_n754), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n720), .B1(new_n748), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n218), .A2(new_n287), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n218), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n242), .A2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n218), .A2(new_n486), .ZN(new_n767));
  INV_X1    g0567(.A(G45), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n225), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n719), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n308), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n203), .B1(new_n777), .B2(G45), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n686), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n762), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n773), .B(KEYINPUT94), .Z(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n675), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n676), .A2(new_n779), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n675), .A2(G330), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT95), .Z(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT96), .Z(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  INV_X1    g0588(.A(new_n779), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n720), .A2(new_n772), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(G77), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n425), .A2(new_n667), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n667), .A2(new_n417), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n428), .B2(new_n429), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(new_n425), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n772), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n380), .B1(new_n723), .B2(new_n797), .C1(new_n728), .C2(new_n534), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G283), .B2(new_n736), .ZN(new_n799));
  INV_X1    g0599(.A(new_n742), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G294), .A2(new_n800), .B1(new_n746), .B2(new_n470), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n743), .A2(new_n460), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(G107), .B2(new_n755), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n799), .A2(new_n740), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n800), .B1(new_n746), .B2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  INV_X1    g0606(.A(G150), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n806), .B2(new_n728), .C1(new_n807), .C2(new_n735), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n743), .A2(new_n222), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G50), .B2(new_n755), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  INV_X1    g0612(.A(G132), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n591), .B1(new_n813), .B2(new_n723), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G58), .B2(new_n759), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n812), .A2(KEYINPUT98), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT98), .B1(new_n812), .B2(new_n815), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n804), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n791), .B(new_n796), .C1(new_n719), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n431), .A2(new_n668), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n647), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n695), .B2(new_n795), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(new_n714), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT99), .Z(new_n826));
  AOI21_X1  g0626(.A(new_n789), .B1(new_n824), .B2(new_n714), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n820), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  NOR2_X1   g0629(.A1(new_n777), .A2(new_n203), .ZN(new_n830));
  INV_X1    g0630(.A(new_n315), .ZN(new_n831));
  INV_X1    g0631(.A(new_n306), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n392), .B1(new_n832), .B2(KEYINPUT16), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n306), .A2(new_n281), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n665), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n318), .B2(new_n329), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n316), .B1(new_n835), .B2(new_n665), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n322), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n324), .A2(new_n664), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n325), .A2(new_n841), .A3(new_n316), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n837), .A2(new_n844), .A3(KEYINPUT38), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT38), .B1(new_n837), .B2(new_n844), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n369), .A2(new_n667), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n353), .B1(new_n348), .B2(new_n350), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n374), .B(new_n848), .C1(new_n849), .C2(new_n371), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n355), .A2(new_n369), .A3(new_n667), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n792), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT100), .B1(new_n823), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT100), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n855), .B(new_n792), .C1(new_n647), .C2(new_n822), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n847), .B(new_n852), .C1(new_n854), .C2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT39), .B1(new_n845), .B2(new_n846), .ZN(new_n858));
  XNOR2_X1  g0658(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n324), .B(new_n664), .C1(new_n318), .C2(new_n329), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n325), .A2(new_n841), .A3(new_n316), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n843), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n859), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n845), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n858), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n370), .A2(new_n667), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n868), .A2(new_n869), .B1(new_n329), .B2(new_n665), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n446), .B(new_n693), .C1(new_n695), .C2(KEYINPUT29), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n658), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n871), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n852), .A2(new_n795), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n710), .B2(new_n711), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n845), .B2(new_n846), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n876), .B(KEYINPUT40), .C1(new_n845), .C2(new_n864), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n446), .A2(new_n712), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n881), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(G330), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n830), .B1(new_n874), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n874), .B2(new_n885), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n607), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n227), .A4(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT36), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n225), .A2(G77), .A3(new_n292), .A4(new_n293), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(G50), .B2(new_n222), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G1), .A3(new_n308), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n887), .A2(new_n891), .A3(new_n894), .ZN(G367));
  OAI21_X1  g0695(.A(new_n629), .B1(new_n617), .B2(new_n668), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n615), .A2(new_n668), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(new_n521), .A3(new_n679), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT103), .Z(new_n901));
  INV_X1    g0701(.A(new_n518), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n615), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n899), .A2(KEYINPUT42), .B1(new_n903), .B2(new_n668), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n585), .B1(new_n565), .B2(new_n668), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n668), .A2(new_n565), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n639), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n901), .A2(new_n904), .B1(KEYINPUT43), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n908), .B(new_n909), .Z(new_n910));
  INV_X1    g0710(.A(new_n898), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n678), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT108), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n778), .B(KEYINPUT107), .Z(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n680), .A2(new_n898), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(KEYINPUT105), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n680), .A2(new_n898), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n926), .B(KEYINPUT45), .Z(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n677), .A2(KEYINPUT106), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n521), .A2(new_n679), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n671), .B2(new_n679), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(new_n676), .Z(new_n933));
  NAND2_X1  g0733(.A1(new_n716), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n930), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n716), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n685), .B(KEYINPUT41), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n917), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n914), .A2(new_n915), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n915), .B1(new_n914), .B2(new_n940), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n774), .B1(new_n218), .B2(new_n412), .C1(new_n238), .C2(new_n767), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n789), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n745), .A2(new_n525), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n755), .A2(KEYINPUT46), .A3(G116), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(G303), .C2(new_n800), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n743), .A2(new_n554), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n949), .B(new_n591), .C1(G317), .C2(new_n756), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n736), .A2(G294), .B1(new_n759), .B2(G107), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n755), .A2(new_n470), .ZN(new_n952));
  XNOR2_X1  g0752(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(G311), .B2(new_n751), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n948), .A2(new_n950), .A3(new_n951), .A4(new_n954), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n733), .A2(new_n221), .B1(new_n723), .B2(new_n806), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT110), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n739), .A2(G68), .ZN(new_n958));
  INV_X1    g0758(.A(G143), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n735), .A2(new_n724), .B1(new_n728), .B2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n742), .A2(new_n807), .B1(new_n745), .B2(new_n361), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n287), .B1(new_n743), .B2(new_n208), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n945), .B1(new_n907), .B2(new_n781), .C1(new_n967), .C2(new_n720), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT112), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n943), .A2(new_n970), .ZN(G387));
  OAI22_X1  g0771(.A1(new_n733), .A2(new_n490), .B1(new_n738), .B2(new_n525), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G317), .A2(new_n800), .B1(new_n746), .B2(G303), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n973), .B1(new_n797), .B2(new_n735), .C1(new_n749), .C2(new_n728), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT48), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n975), .B2(new_n974), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT49), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n470), .A2(new_n753), .B1(new_n756), .B2(G326), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n979), .A2(new_n486), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n486), .B(new_n949), .C1(G77), .C2(new_n755), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n739), .A2(new_n413), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n742), .A2(new_n361), .B1(new_n745), .B2(new_n222), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G150), .B2(new_n756), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G159), .A2(new_n751), .B1(new_n736), .B2(new_n393), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n983), .A2(new_n984), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n720), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n763), .A2(new_n687), .B1(G107), .B2(new_n218), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n235), .A2(G45), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n311), .A2(KEYINPUT50), .A3(G50), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT50), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n393), .B2(new_n361), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT113), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n687), .B(new_n768), .C1(new_n222), .C2(new_n208), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n992), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n995), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n767), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n990), .B1(new_n991), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n789), .B1(new_n1000), .B2(new_n775), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n781), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n989), .B(new_n1001), .C1(new_n672), .C2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n933), .B2(new_n917), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n934), .A2(new_n685), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n716), .A2(new_n933), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(G393));
  AOI21_X1  g0807(.A(new_n686), .B1(new_n930), .B2(new_n935), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n935), .B2(new_n930), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n930), .A2(new_n917), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n911), .A2(new_n773), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n751), .A2(G317), .B1(new_n800), .B2(G311), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n745), .A2(new_n490), .B1(new_n723), .B2(new_n749), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G283), .B2(new_n755), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n380), .B1(new_n743), .B2(new_n421), .C1(new_n735), .C2(new_n534), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n470), .B2(new_n759), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n728), .A2(new_n807), .B1(new_n742), .B2(new_n724), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT51), .Z(new_n1020));
  OAI22_X1  g0820(.A1(new_n745), .A2(new_n311), .B1(new_n723), .B2(new_n959), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n802), .B(new_n1021), .C1(G68), .C2(new_n755), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n739), .A2(G77), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n486), .B1(G50), .B2(new_n736), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1018), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n719), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n774), .B1(new_n554), .B2(new_n218), .C1(new_n245), .C2(new_n767), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1011), .A2(new_n789), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1009), .A2(new_n1010), .A3(new_n1029), .ZN(G390));
  NAND2_X1  g0830(.A1(new_n446), .A2(new_n713), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n872), .A2(new_n658), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n712), .A2(G330), .A3(new_n795), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1034), .A2(new_n852), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n852), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n854), .A2(new_n856), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1037), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n794), .A2(new_n425), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n792), .B1(new_n692), .B2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n852), .B(KEYINPUT114), .Z(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1041), .C1(new_n1034), .C2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1032), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n868), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n821), .B1(new_n694), .B2(new_n637), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n855), .B1(new_n1047), .B2(new_n792), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n823), .A2(KEYINPUT100), .A3(new_n853), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1036), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1050), .B2(new_n869), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n869), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1042), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1052), .B(new_n865), .C1(new_n1041), .C2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1051), .A2(new_n1039), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1039), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1045), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n852), .B1(new_n854), .B2(new_n856), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n868), .B1(new_n1059), .B2(new_n1052), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1054), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1037), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1062), .A2(new_n1055), .A3(new_n1044), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(new_n685), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n789), .B1(new_n393), .B2(new_n790), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n868), .A2(new_n772), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n745), .A2(new_n554), .B1(new_n723), .B2(new_n490), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n810), .B(new_n1067), .C1(G116), .C2(new_n800), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n380), .B1(new_n733), .B2(new_n460), .C1(new_n525), .C2(new_n728), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G107), .B2(new_n736), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(new_n1070), .A3(new_n1023), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n742), .A2(new_n813), .B1(new_n743), .B2(new_n361), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n380), .B(new_n1072), .C1(G125), .C2(new_n756), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n736), .A2(G137), .B1(new_n751), .B2(G128), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n733), .A2(new_n807), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT53), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT54), .B(G143), .Z(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n746), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .A4(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n739), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1081), .A2(new_n724), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1071), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1065), .B(new_n1066), .C1(new_n719), .C2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1084), .B1(new_n1085), .B2(new_n917), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1064), .A2(new_n1086), .ZN(G378));
  NOR2_X1   g0887(.A1(new_n434), .A2(new_n398), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n665), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n655), .B2(new_n409), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1091), .B(new_n649), .C1(new_n651), .C2(new_n654), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR3_X1   g0895(.A1(new_n439), .A2(new_n442), .A3(new_n650), .ZN(new_n1096));
  AOI21_X1  g0896(.A(KEYINPUT89), .B1(new_n652), .B2(new_n653), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n409), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n1091), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n655), .A2(new_n409), .A3(new_n1092), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(new_n1100), .A3(new_n1089), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1095), .A2(new_n1101), .A3(new_n771), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n789), .B1(G50), .B2(new_n790), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n591), .A2(G41), .ZN(new_n1104));
  AOI211_X1 g0904(.A(G50), .B(new_n1104), .C1(new_n266), .C2(new_n496), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n742), .A2(new_n421), .B1(new_n745), .B2(new_n412), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1104), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G283), .C2(new_n756), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G77), .A2(new_n755), .B1(new_n753), .B2(G58), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n554), .B2(new_n735), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n751), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n958), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT58), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1105), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G128), .A2(new_n800), .B1(new_n746), .B2(G137), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n751), .A2(G125), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n813), .C2(new_n735), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1078), .A2(new_n755), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1118), .A2(KEYINPUT116), .B1(new_n1081), .B2(new_n807), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1117), .B(new_n1119), .C1(KEYINPUT116), .C2(new_n1118), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT59), .Z(new_n1121));
  AOI211_X1 g0921(.A(G33), .B(G41), .C1(new_n756), .C2(G124), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n724), .B2(new_n743), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1114), .B1(new_n1113), .B2(new_n1112), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1103), .B1(new_n1124), .B2(new_n719), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1102), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n879), .A2(G330), .A3(new_n880), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1095), .A2(new_n1101), .A3(KEYINPUT118), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1095), .A2(new_n1101), .A3(KEYINPUT118), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1132), .A2(G330), .A3(new_n879), .A4(new_n880), .ZN(new_n1133));
  AND4_X1   g0933(.A1(new_n857), .A2(new_n1131), .A3(new_n870), .A4(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n857), .A2(new_n870), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1136), .B2(new_n916), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT57), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1032), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1139), .C1(new_n1063), .C2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1063), .A2(new_n1140), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1139), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1136), .B1(new_n1063), .B2(new_n1140), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n685), .B1(new_n1146), .B2(KEYINPUT57), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1137), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(G375));
  AOI22_X1  g0950(.A1(G159), .A2(new_n755), .B1(new_n756), .B2(G128), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT121), .Z(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n361), .B2(new_n1081), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1078), .A2(new_n736), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n742), .A2(new_n806), .B1(new_n743), .B2(new_n221), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G150), .B2(new_n746), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n486), .B1(G132), .B2(new_n751), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n733), .A2(new_n554), .B1(new_n723), .B2(new_n534), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT120), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n287), .B1(new_n753), .B2(G77), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G283), .A2(new_n800), .B1(new_n746), .B2(G107), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n470), .A2(new_n736), .B1(new_n751), .B2(G294), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n984), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1153), .A2(new_n1158), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n719), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n789), .C1(G68), .C2(new_n790), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1053), .B2(new_n771), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n917), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1045), .A2(new_n939), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1169), .A2(new_n1140), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(G381));
  AOI211_X1 g0973(.A(new_n969), .B(G390), .C1(new_n941), .C2(new_n942), .ZN(new_n1174));
  OR2_X1    g0974(.A1(G396), .A2(G393), .ZN(new_n1175));
  NOR4_X1   g0975(.A1(G378), .A2(G384), .A3(G381), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1149), .A3(new_n1176), .ZN(G407));
  INV_X1    g0977(.A(G378), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n666), .A2(G213), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1149), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(G407), .A2(G213), .A3(new_n1181), .ZN(G409));
  AOI21_X1  g0982(.A(new_n938), .B1(new_n1063), .B2(new_n1140), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1183), .A2(new_n917), .B1(new_n1135), .B2(new_n1134), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G378), .B1(new_n1184), .B2(new_n1126), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1149), .B2(G378), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT62), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1172), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1044), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n686), .B1(new_n1172), .B2(KEYINPUT60), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT123), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(KEYINPUT123), .A3(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(G384), .A3(new_n1170), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G384), .B1(new_n1198), .B2(new_n1170), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1137), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1138), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1142), .A2(KEYINPUT119), .A3(new_n1143), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(G378), .B(new_n1203), .C1(new_n1207), .C2(new_n1147), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1185), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(KEYINPUT122), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1188), .A2(new_n1189), .A3(new_n1202), .A4(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(KEYINPUT125), .B1(new_n1186), .B2(new_n1180), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT125), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1210), .A2(new_n1214), .A3(new_n1179), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1180), .A2(G2897), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT124), .Z(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1201), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1199), .A3(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1213), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT61), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1212), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1189), .B1(new_n1226), .B2(new_n1202), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT126), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1214), .B1(new_n1210), .B2(new_n1179), .ZN(new_n1229));
  AOI211_X1 g1029(.A(KEYINPUT125), .B(new_n1180), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1222), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1202), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1234), .A3(new_n1235), .A4(new_n1212), .ZN(new_n1236));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n943), .B2(new_n970), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1174), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(G393), .B(new_n787), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1238), .B2(new_n1174), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1243), .A2(new_n1244), .A3(KEYINPUT127), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT127), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1228), .A2(new_n1236), .A3(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(KEYINPUT61), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1188), .A2(new_n1202), .A3(new_n1211), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1202), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1188), .A2(new_n1211), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1222), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1250), .A2(new_n1253), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1248), .A2(new_n1257), .ZN(G405));
  XNOR2_X1  g1058(.A(new_n1149), .B(G378), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(new_n1202), .Z(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(new_n1249), .Z(G402));
endmodule


