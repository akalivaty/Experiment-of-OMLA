//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT74), .Z(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(KEYINPUT28), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT68), .B1(new_n208), .B2(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n205), .ZN(new_n210));
  AOI211_X1 g009(.A(G190gat), .B(new_n209), .C1(KEYINPUT68), .C2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n211), .B2(KEYINPUT28), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n213), .A2(new_n206), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n215), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(KEYINPUT26), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n214), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n216), .A2(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n219), .B1(new_n215), .B2(KEYINPUT23), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(new_n214), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT67), .Z(new_n232));
  NOR2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(KEYINPUT24), .B2(new_n214), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT64), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n235), .B(new_n239), .C1(KEYINPUT24), .C2(new_n214), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n226), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n242), .A2(new_n227), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n224), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n204), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247));
  INV_X1    g046(.A(new_n203), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n246), .A2(new_n247), .B1(new_n244), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n245), .ZN(new_n250));
  INV_X1    g049(.A(new_n204), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT75), .ZN(new_n253));
  XNOR2_X1  g052(.A(G197gat), .B(G204gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255));
  INV_X1    g054(.A(G211gat), .ZN(new_n256));
  INV_X1    g055(.A(G218gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G211gat), .B(G218gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n260), .A2(new_n254), .A3(new_n258), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT73), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n253), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n263), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n250), .A2(new_n203), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n244), .A2(new_n204), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(new_n266), .B2(new_n267), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n202), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT38), .ZN(new_n275));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n265), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n250), .A2(new_n247), .A3(new_n251), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n244), .A2(new_n248), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n246), .A2(new_n247), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n269), .A3(new_n271), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n275), .B(new_n279), .C1(new_n287), .C2(KEYINPUT37), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n274), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G141gat), .B(G148gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT76), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  OR2_X1    g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(KEYINPUT2), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n291), .C2(KEYINPUT2), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  OR2_X1    g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(G134gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n300), .B(new_n301), .C1(KEYINPUT69), .C2(KEYINPUT1), .ZN(new_n302));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT1), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n302), .B(new_n304), .Z(new_n305));
  NOR2_X1   g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n302), .B(new_n304), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT77), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n308), .B2(new_n298), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n309), .A2(KEYINPUT5), .A3(G225gat), .A4(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT5), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n313), .B1(KEYINPUT4), .B2(new_n306), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n298), .A2(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(KEYINPUT77), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n317), .A3(new_n297), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n315), .A2(new_n316), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT78), .A3(new_n315), .A4(new_n318), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n296), .A2(new_n297), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n330), .A2(KEYINPUT80), .A3(new_n312), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n332), .B1(new_n306), .B2(new_n311), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(KEYINPUT4), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT5), .B1(new_n335), .B2(new_n325), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n310), .B1(new_n328), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT0), .ZN(new_n339));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n310), .C1(new_n328), .C2(new_n336), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n279), .B1(new_n287), .B2(KEYINPUT37), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n265), .B1(new_n249), .B2(new_n253), .ZN(new_n351));
  INV_X1    g150(.A(new_n286), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n202), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT38), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n285), .A2(new_n286), .A3(new_n278), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n290), .A2(new_n349), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G78gat), .ZN(new_n358));
  INV_X1    g157(.A(G228gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n269), .A2(new_n245), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(KEYINPUT81), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT3), .B1(new_n362), .B2(KEYINPUT81), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n298), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n318), .A2(new_n245), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n264), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n318), .A2(new_n245), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n265), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n315), .B(new_n361), .C1(new_n329), .C2(new_n362), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(G22gat), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n371), .A2(new_n372), .ZN(new_n375));
  INV_X1    g174(.A(new_n368), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n329), .B1(new_n363), .B2(new_n364), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n376), .A2(new_n377), .B1(new_n359), .B2(new_n360), .ZN(new_n378));
  INV_X1    g177(.A(G22gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n375), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n358), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n374), .A2(new_n380), .A3(new_n358), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  INV_X1    g183(.A(G106gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  INV_X1    g187(.A(new_n383), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n381), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT40), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n327), .B1(new_n335), .B2(new_n325), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT39), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n341), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n309), .A2(new_n327), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT39), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n342), .B1(new_n394), .B2(new_n395), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n402), .B(KEYINPUT40), .C1(new_n394), .C2(new_n399), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n343), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n279), .B1(new_n351), .B2(new_n352), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n356), .A3(KEYINPUT30), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n353), .A2(new_n407), .A3(new_n278), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n392), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n357), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G227gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n244), .A2(new_n307), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n224), .B(new_n305), .C1(new_n236), .C2(new_n243), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(new_n417), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n414), .A3(new_n416), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n424), .B(KEYINPUT32), .C1(new_n425), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(KEYINPUT32), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n425), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n428), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT71), .B1(new_n417), .B2(new_n419), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n423), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n430), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n415), .A2(new_n416), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n421), .B(new_n418), .C1(new_n437), .C2(new_n414), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n422), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n435), .B1(new_n441), .B2(KEYINPUT72), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT72), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n436), .B2(new_n440), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT36), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n435), .A2(new_n441), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n446), .A2(KEYINPUT36), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n346), .A2(new_n347), .B1(new_n406), .B2(new_n408), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n447), .C1(new_n448), .C2(new_n392), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n442), .A2(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n392), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n348), .A2(new_n409), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT35), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n391), .A2(new_n446), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT35), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n448), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n412), .A2(new_n450), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G229gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT13), .ZN(new_n460));
  INV_X1    g259(.A(G43gat), .ZN(new_n461));
  INV_X1    g260(.A(G50gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G43gat), .A2(G50gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT83), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(KEYINPUT83), .A3(new_n464), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(KEYINPUT15), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G29gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n470), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n471));
  INV_X1    g270(.A(G36gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT14), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(G29gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(KEYINPUT15), .B2(new_n465), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n467), .A2(new_n476), .A3(KEYINPUT15), .A4(new_n468), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G8gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  OR2_X1    g281(.A1(new_n482), .A2(G1gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT16), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n484), .B2(G1gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n483), .A2(new_n481), .A3(new_n485), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n486), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n478), .A2(new_n479), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n460), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(KEYINPUT17), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n494), .A3(new_n479), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n459), .A3(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT18), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n496), .A2(KEYINPUT18), .A3(new_n488), .A4(new_n459), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(new_n501), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(G197gat), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT11), .B(G169gat), .Z(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT12), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n509), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(KEYINPUT85), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n504), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n458), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G71gat), .B(G78gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G57gat), .B(G64gat), .Z(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  INV_X1    g322(.A(G71gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n358), .A3(KEYINPUT9), .ZN(new_n525));
  NAND2_X1  g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G64gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(KEYINPUT86), .A3(G57gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT88), .ZN(new_n536));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT20), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n536), .A2(new_n538), .ZN(new_n540));
  XOR2_X1   g339(.A(G183gat), .B(G211gat), .Z(new_n541));
  OR3_X1    g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  AOI211_X1 g344(.A(new_n486), .B(new_n487), .C1(new_n545), .C2(KEYINPUT21), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n546), .B(new_n549), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n542), .A2(new_n550), .A3(new_n543), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G232gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT90), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT41), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G85gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT91), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G85gat), .ZN(new_n565));
  INV_X1    g364(.A(G92gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT7), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G99gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT8), .B1(new_n573), .B2(new_n385), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT92), .ZN(new_n576));
  XOR2_X1   g375(.A(G99gat), .B(G106gat), .Z(new_n577));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n567), .A2(new_n572), .A3(new_n578), .A4(new_n574), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n577), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n585), .B1(G99gat), .B2(G106gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT91), .B(G85gat), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n566), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n578), .B1(new_n588), .B2(new_n572), .ZN(new_n589));
  INV_X1    g388(.A(new_n579), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n584), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT93), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT94), .B1(new_n583), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n493), .A2(new_n495), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT94), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n591), .A2(KEYINPUT93), .A3(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n480), .A3(new_n598), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n556), .A2(new_n557), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n605), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n561), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n600), .B2(new_n603), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n608), .B(new_n561), .C1(new_n611), .C2(KEYINPUT95), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(KEYINPUT95), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n608), .A2(new_n561), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n611), .A2(KEYINPUT95), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT96), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n609), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n554), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G230gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(new_n360), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n545), .A2(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n596), .A2(new_n598), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT97), .B(KEYINPUT10), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n531), .B1(new_n580), .B2(new_n581), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n591), .A2(new_n592), .A3(new_n545), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n624), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n580), .A2(new_n581), .A3(new_n531), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n545), .B1(new_n591), .B2(new_n592), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n634), .A2(new_n635), .A3(new_n624), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  NAND3_X1  g439(.A1(new_n633), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n633), .B2(new_n637), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n621), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n517), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n348), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n346), .A2(KEYINPUT98), .A3(new_n347), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT99), .B(G1gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  INV_X1    g453(.A(new_n409), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n517), .A2(new_n655), .A3(new_n646), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT16), .B(G8gat), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n656), .A2(KEYINPUT100), .A3(G8gat), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n656), .B2(G8gat), .ZN(new_n662));
  OAI22_X1  g461(.A1(new_n659), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(G1325gat));
  NAND2_X1  g462(.A1(new_n445), .A2(new_n447), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G15gat), .B1(new_n647), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n446), .A2(G15gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n647), .B2(new_n667), .ZN(G1326gat));
  OR3_X1    g467(.A1(new_n647), .A2(KEYINPUT101), .A3(new_n392), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT101), .B1(new_n647), .B2(new_n392), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(new_n554), .ZN(new_n675));
  INV_X1    g474(.A(new_n620), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n644), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n517), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n651), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n470), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n458), .B2(new_n620), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n346), .A2(new_n356), .A3(new_n347), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n289), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n410), .B1(new_n687), .B2(new_n355), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n442), .A2(new_n391), .A3(new_n444), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n456), .B1(new_n689), .B2(new_n448), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n448), .A2(new_n456), .A3(new_n455), .ZN(new_n691));
  OAI22_X1  g490(.A1(new_n688), .A2(new_n449), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(KEYINPUT44), .A3(new_n676), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n554), .A2(new_n516), .A3(new_n645), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(G29gat), .B1(new_n696), .B2(new_n651), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n683), .A2(new_n697), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n679), .A2(G36gat), .A3(new_n409), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT46), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G36gat), .B1(new_n696), .B2(new_n409), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1329gat));
  NAND4_X1  g502(.A1(new_n685), .A2(new_n664), .A3(new_n693), .A4(new_n695), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(new_n461), .ZN(new_n708));
  INV_X1    g507(.A(new_n446), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n680), .A2(new_n461), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n704), .A2(G43gat), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n708), .A2(new_n711), .B1(new_n713), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g513(.A1(new_n679), .A2(KEYINPUT105), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n517), .A2(new_n716), .A3(new_n678), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n715), .A2(new_n462), .A3(new_n391), .A4(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n685), .A2(new_n391), .A3(new_n693), .A4(new_n695), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n719), .B1(new_n718), .B2(new_n721), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n722), .A2(new_n723), .ZN(G1331gat));
  INV_X1    g523(.A(new_n516), .ZN(new_n725));
  NOR4_X1   g524(.A1(new_n458), .A2(new_n725), .A3(new_n621), .A4(new_n644), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n681), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g527(.A(new_n409), .B(KEYINPUT106), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n726), .B(new_n730), .C1(new_n731), .C2(new_n528), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n528), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1333gat));
  AOI21_X1  g533(.A(new_n524), .B1(new_n726), .B2(new_n664), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n446), .A2(G71gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n726), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1334gat));
  NAND2_X1  g538(.A1(new_n726), .A2(new_n391), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g540(.A1(new_n554), .A2(new_n725), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n692), .A2(new_n676), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n692), .A2(new_n745), .A3(new_n676), .A4(new_n742), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n744), .A2(new_n645), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n587), .A3(new_n681), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n554), .A2(new_n725), .A3(new_n644), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n694), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n651), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n751), .B2(new_n587), .ZN(G1336gat));
  NAND4_X1  g551(.A1(new_n685), .A2(new_n655), .A3(new_n693), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n729), .A2(G92gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n744), .A2(new_n645), .A3(new_n746), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT52), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n685), .A2(new_n693), .A3(new_n730), .A4(new_n749), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G92gat), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT108), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AND4_X1   g562(.A1(KEYINPUT108), .A2(new_n762), .A3(new_n759), .A4(new_n756), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n758), .B1(new_n763), .B2(new_n764), .ZN(G1337gat));
  XOR2_X1   g564(.A(KEYINPUT109), .B(G99gat), .Z(new_n766));
  NAND3_X1  g565(.A1(new_n747), .A2(new_n709), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n665), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n766), .ZN(G1338gat));
  NOR2_X1   g568(.A1(new_n392), .A2(new_n385), .ZN(new_n770));
  AND4_X1   g569(.A1(new_n685), .A2(new_n693), .A3(new_n749), .A4(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n744), .A2(new_n391), .A3(new_n645), .A4(new_n746), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n385), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT53), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n772), .A2(new_n385), .ZN(new_n777));
  OAI211_X1 g576(.A(KEYINPUT110), .B(new_n776), .C1(new_n777), .C2(new_n771), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1339gat));
  AOI21_X1  g578(.A(new_n459), .B1(new_n496), .B2(new_n488), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n488), .A2(new_n491), .A3(new_n460), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n508), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n512), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n645), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(new_n623), .A3(new_n626), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n785), .A2(new_n788), .A3(new_n623), .A4(new_n626), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n787), .A2(KEYINPUT54), .A3(new_n633), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n623), .B1(new_n785), .B2(new_n626), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n640), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(KEYINPUT55), .A3(new_n793), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(new_n641), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n784), .B1(new_n798), .B2(new_n516), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n620), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n796), .A2(new_n641), .A3(new_n797), .A4(new_n783), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n620), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n554), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n554), .A2(new_n516), .A3(new_n644), .A4(new_n620), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT112), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n620), .A2(new_n801), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n620), .B2(new_n799), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n807), .B(new_n804), .C1(new_n809), .C2(new_n554), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n651), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n729), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n516), .A2(G113gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n689), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n811), .A2(new_n455), .A3(new_n725), .A4(new_n729), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n815), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n815), .B2(G113gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT114), .ZN(G1340gat));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n455), .A3(new_n645), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G120gat), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n644), .A2(G120gat), .ZN(new_n822));
  XOR2_X1   g621(.A(new_n822), .B(KEYINPUT115), .Z(new_n823));
  NAND3_X1  g622(.A1(new_n812), .A2(new_n689), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n825), .B(new_n826), .ZN(G1341gat));
  NOR2_X1   g626(.A1(new_n675), .A2(new_n299), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n812), .A2(new_n455), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n689), .A3(new_n554), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n299), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n812), .A2(new_n833), .A3(new_n455), .A4(new_n828), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT118), .A4(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n812), .A2(new_n455), .A3(new_n676), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G134gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n676), .A2(new_n409), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n452), .A2(new_n842), .A3(G134gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n811), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT119), .B1(new_n844), .B2(KEYINPUT56), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n844), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n846));
  OAI221_X1 g645(.A(new_n841), .B1(KEYINPUT56), .B2(new_n844), .C1(new_n845), .C2(new_n846), .ZN(G1343gat));
  NAND3_X1  g646(.A1(new_n681), .A2(new_n665), .A3(new_n729), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n392), .B(new_n848), .C1(new_n806), .C2(new_n810), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n725), .ZN(new_n850));
  INV_X1    g649(.A(G141gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n681), .A2(new_n665), .A3(KEYINPUT120), .A4(new_n729), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n804), .B1(new_n809), .B2(new_n554), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n391), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n392), .B1(new_n806), .B2(new_n810), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n857), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n725), .A2(G141gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n852), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(G1344gat));
  INV_X1    g666(.A(G148gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(KEYINPUT59), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n869), .B1(new_n863), .B2(new_n644), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n858), .A2(new_n857), .A3(new_n391), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n645), .B(new_n871), .C1(new_n861), .C2(new_n857), .ZN(new_n872));
  OAI21_X1  g671(.A(G148gat), .B1(new_n872), .B2(new_n856), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(KEYINPUT121), .A3(KEYINPUT59), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT121), .B1(new_n873), .B2(KEYINPUT59), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n868), .A3(new_n645), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1345gat));
  INV_X1    g677(.A(G155gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n849), .A2(new_n879), .A3(new_n554), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n863), .A2(new_n675), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n879), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n880), .C1(new_n881), .C2(new_n879), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n863), .B2(new_n620), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n651), .A2(new_n664), .A3(G162gat), .A4(new_n842), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n861), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(G1347gat));
  INV_X1    g689(.A(G169gat), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n806), .A2(new_n810), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n651), .ZN(new_n894));
  AOI211_X1 g693(.A(KEYINPUT123), .B(new_n681), .C1(new_n806), .C2(new_n810), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n689), .B(new_n730), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n891), .B1(new_n896), .B2(new_n516), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n651), .A2(new_n655), .A3(new_n455), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n806), .B2(new_n810), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(G169gat), .A3(new_n725), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT124), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n899), .A2(G176gat), .A3(new_n645), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT125), .Z(new_n907));
  OR2_X1    g706(.A1(new_n896), .A2(new_n644), .ZN(new_n908));
  INV_X1    g707(.A(G176gat), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n554), .A2(new_n205), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n899), .A2(new_n554), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n896), .A2(new_n911), .B1(new_n912), .B2(new_n213), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g713(.A1(new_n676), .A2(new_n206), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n676), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(G190gat), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT61), .B(new_n206), .C1(new_n899), .C2(new_n676), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n896), .A2(new_n915), .B1(new_n918), .B2(new_n919), .ZN(G1351gat));
  INV_X1    g719(.A(G197gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n729), .A2(new_n664), .A3(new_n392), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n894), .B2(new_n895), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n516), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n651), .A2(new_n655), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(new_n664), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n871), .B(new_n926), .C1(new_n861), .C2(new_n857), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n725), .A2(G197gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n924), .B(new_n931), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1352gat));
  NOR2_X1   g732(.A1(new_n644), .A2(G204gat), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n922), .B(new_n934), .C1(new_n894), .C2(new_n895), .ZN(new_n935));
  OR3_X1    g734(.A1(new_n935), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n935), .B2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(KEYINPUT62), .ZN(new_n938));
  INV_X1    g737(.A(new_n926), .ZN(new_n939));
  OAI21_X1  g738(.A(G204gat), .B1(new_n872), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(G1353gat));
  OR2_X1    g740(.A1(new_n927), .A2(new_n675), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n554), .A2(new_n256), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n944), .A2(new_n945), .B1(new_n923), .B2(new_n946), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n927), .B2(new_n620), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n676), .A2(new_n257), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n923), .B2(new_n949), .ZN(G1355gat));
endmodule


