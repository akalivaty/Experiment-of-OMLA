

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X2 U322 ( .A(n389), .B(n388), .ZN(n513) );
  XNOR2_X1 U323 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n376) );
  OR2_X1 U324 ( .A1(n465), .A2(n464), .ZN(n479) );
  XOR2_X1 U325 ( .A(n335), .B(n334), .Z(n290) );
  XNOR2_X1 U326 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n361) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n363) );
  NOR2_X1 U328 ( .A1(n520), .A2(n525), .ZN(n454) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U330 ( .A(n336), .B(n290), .ZN(n337) );
  XNOR2_X1 U331 ( .A(n375), .B(n374), .ZN(n521) );
  NOR2_X1 U332 ( .A1(n578), .A2(n481), .ZN(n482) );
  XNOR2_X1 U333 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U334 ( .A(n447), .B(n446), .ZN(n522) );
  XNOR2_X1 U335 ( .A(n484), .B(KEYINPUT38), .ZN(n492) );
  XNOR2_X1 U336 ( .A(n449), .B(KEYINPUT58), .ZN(n450) );
  XNOR2_X1 U337 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U338 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n292) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G29GAT), .ZN(n291) );
  XNOR2_X1 U341 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U342 ( .A(KEYINPUT71), .B(n293), .Z(n360) );
  INV_X1 U343 ( .A(n360), .ZN(n309) );
  XOR2_X1 U344 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n295) );
  XNOR2_X1 U345 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n307) );
  XOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .Z(n380) );
  XOR2_X1 U348 ( .A(KEYINPUT11), .B(n380), .Z(n297) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G85GAT), .Z(n328) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(n328), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n303) );
  XNOR2_X1 U352 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n298), .B(G162GAT), .ZN(n424) );
  INV_X1 U354 ( .A(KEYINPUT66), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n424), .B(n299), .ZN(n301) );
  NAND2_X1 U356 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U358 ( .A(n303), .B(n302), .Z(n305) );
  XNOR2_X1 U359 ( .A(G134GAT), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n535) );
  INV_X1 U363 ( .A(n535), .ZN(n550) );
  XNOR2_X1 U364 ( .A(G71GAT), .B(G57GAT), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n310), .B(KEYINPUT13), .ZN(n333) );
  XOR2_X1 U366 ( .A(G8GAT), .B(G183GAT), .Z(n311) );
  XOR2_X1 U367 ( .A(G211GAT), .B(n311), .Z(n383) );
  XOR2_X1 U368 ( .A(n333), .B(n383), .Z(n324) );
  XOR2_X1 U369 ( .A(G22GAT), .B(G155GAT), .Z(n415) );
  XOR2_X1 U370 ( .A(G15GAT), .B(G127GAT), .Z(n433) );
  XOR2_X1 U371 ( .A(n415), .B(n433), .Z(n313) );
  NAND2_X1 U372 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U374 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U377 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT72), .B(G1GAT), .Z(n352) );
  XOR2_X1 U379 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n319) );
  XNOR2_X1 U380 ( .A(G78GAT), .B(G64GAT), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U382 ( .A(n352), .B(n320), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U384 ( .A(n324), .B(n323), .Z(n573) );
  XOR2_X1 U385 ( .A(KEYINPUT112), .B(n573), .Z(n560) );
  XOR2_X1 U386 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n326) );
  XNOR2_X1 U387 ( .A(G120GAT), .B(G204GAT), .ZN(n325) );
  XOR2_X1 U388 ( .A(n326), .B(n325), .Z(n340) );
  XNOR2_X1 U389 ( .A(G176GAT), .B(G92GAT), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n327), .B(G64GAT), .ZN(n387) );
  XOR2_X1 U391 ( .A(n387), .B(n328), .Z(n330) );
  NAND2_X1 U392 ( .A1(G230GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n338) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n423) );
  XNOR2_X1 U397 ( .A(n423), .B(n333), .ZN(n336) );
  XOR2_X1 U398 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n335) );
  XNOR2_X1 U399 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n570) );
  XOR2_X1 U401 ( .A(n570), .B(KEYINPUT41), .Z(n556) );
  XOR2_X1 U402 ( .A(G22GAT), .B(G141GAT), .Z(n342) );
  XNOR2_X1 U403 ( .A(G15GAT), .B(G197GAT), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(G8GAT), .Z(n344) );
  XNOR2_X1 U406 ( .A(KEYINPUT68), .B(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U408 ( .A(n346), .B(n345), .Z(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT74), .B(KEYINPUT69), .Z(n348) );
  XNOR2_X1 U410 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n356) );
  XOR2_X1 U412 ( .A(G113GAT), .B(G50GAT), .Z(n350) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U415 ( .A(n352), .B(n351), .Z(n354) );
  NAND2_X1 U416 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U420 ( .A(n360), .B(n359), .Z(n526) );
  INV_X1 U421 ( .A(n526), .ZN(n565) );
  OR2_X1 U422 ( .A1(n556), .A2(n565), .ZN(n362) );
  NOR2_X1 U423 ( .A1(n560), .A2(n363), .ZN(n364) );
  NAND2_X1 U424 ( .A1(n364), .A2(n550), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n365), .B(KEYINPUT47), .ZN(n373) );
  INV_X1 U426 ( .A(n570), .ZN(n371) );
  XOR2_X1 U427 ( .A(KEYINPUT36), .B(KEYINPUT100), .Z(n366) );
  XNOR2_X1 U428 ( .A(n535), .B(n366), .ZN(n578) );
  NOR2_X1 U429 ( .A1(n573), .A2(n578), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n367), .B(KEYINPUT114), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n368), .B(KEYINPUT45), .ZN(n369) );
  NAND2_X1 U432 ( .A1(n369), .A2(n565), .ZN(n370) );
  NOR2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n372) );
  NOR2_X1 U434 ( .A1(n373), .A2(n372), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n376), .B(KEYINPUT21), .ZN(n377) );
  XOR2_X1 U436 ( .A(n377), .B(KEYINPUT88), .Z(n379) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(G218GAT), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n379), .B(n378), .ZN(n428) );
  XOR2_X1 U439 ( .A(n380), .B(n428), .Z(n382) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U442 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U443 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n386) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n442) );
  XNOR2_X1 U446 ( .A(n442), .B(n387), .ZN(n388) );
  XOR2_X1 U447 ( .A(KEYINPUT122), .B(n513), .Z(n390) );
  NOR2_X1 U448 ( .A1(n521), .A2(n390), .ZN(n392) );
  INV_X1 U449 ( .A(KEYINPUT54), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n414) );
  XOR2_X1 U451 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n394) );
  XNOR2_X1 U452 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n413) );
  XOR2_X1 U454 ( .A(G155GAT), .B(G148GAT), .Z(n396) );
  XNOR2_X1 U455 ( .A(G127GAT), .B(G162GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U457 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n398) );
  XNOR2_X1 U458 ( .A(G1GAT), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U460 ( .A(n400), .B(n399), .Z(n406) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n401), .B(KEYINPUT2), .ZN(n416) );
  XOR2_X1 U463 ( .A(G85GAT), .B(n416), .Z(n403) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U468 ( .A(n407), .B(KEYINPUT6), .Z(n411) );
  XOR2_X1 U469 ( .A(G120GAT), .B(KEYINPUT0), .Z(n409) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(G134GAT), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n443) );
  XNOR2_X1 U472 ( .A(n443), .B(KEYINPUT92), .ZN(n410) );
  XNOR2_X1 U473 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X2 U474 ( .A(n413), .B(n412), .Z(n510) );
  NOR2_X1 U475 ( .A1(n414), .A2(n510), .ZN(n564) );
  XOR2_X1 U476 ( .A(n416), .B(n415), .Z(n418) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U479 ( .A(G211GAT), .B(KEYINPUT24), .Z(n420) );
  XNOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U482 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U485 ( .A(n428), .B(n427), .ZN(n458) );
  NAND2_X1 U486 ( .A1(n564), .A2(n458), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n429), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U488 ( .A(G183GAT), .B(G190GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(G43GAT), .B(G99GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U491 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT83), .B(G71GAT), .Z(n437) );
  XNOR2_X1 U495 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U497 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n439) );
  XNOR2_X1 U498 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n448), .A2(n522), .ZN(n559) );
  NOR2_X1 U504 ( .A1(n550), .A2(n559), .ZN(n451) );
  INV_X1 U505 ( .A(G190GAT), .ZN(n449) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n471) );
  XOR2_X1 U507 ( .A(KEYINPUT98), .B(KEYINPUT34), .Z(n469) );
  NAND2_X1 U508 ( .A1(n526), .A2(n570), .ZN(n483) );
  NOR2_X1 U509 ( .A1(n573), .A2(n535), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n452), .B(KEYINPUT16), .ZN(n466) );
  XNOR2_X1 U511 ( .A(n513), .B(KEYINPUT27), .ZN(n460) );
  NAND2_X1 U512 ( .A1(n510), .A2(n460), .ZN(n520) );
  XNOR2_X1 U513 ( .A(KEYINPUT67), .B(KEYINPUT28), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(n458), .ZN(n525) );
  XOR2_X1 U515 ( .A(KEYINPUT94), .B(n454), .Z(n455) );
  NOR2_X1 U516 ( .A1(n522), .A2(n455), .ZN(n465) );
  NAND2_X1 U517 ( .A1(n513), .A2(n522), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n458), .A2(n456), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n457), .B(KEYINPUT25), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n522), .A2(n458), .ZN(n459) );
  XNOR2_X1 U521 ( .A(KEYINPUT26), .B(n459), .ZN(n563) );
  AND2_X1 U522 ( .A1(n460), .A2(n563), .ZN(n461) );
  NOR2_X1 U523 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n510), .A2(n463), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n466), .A2(n479), .ZN(n497) );
  NOR2_X1 U526 ( .A1(n483), .A2(n497), .ZN(n467) );
  XOR2_X1 U527 ( .A(KEYINPUT95), .B(n467), .Z(n477) );
  NAND2_X1 U528 ( .A1(n477), .A2(n510), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT96), .B(n472), .ZN(G1324GAT) );
  NAND2_X1 U532 ( .A1(n477), .A2(n513), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n475) );
  NAND2_X1 U535 ( .A1(n477), .A2(n522), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U537 ( .A(G15GAT), .B(n476), .Z(G1326GAT) );
  NAND2_X1 U538 ( .A1(n525), .A2(n477), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G22GAT), .ZN(G1327GAT) );
  AND2_X1 U540 ( .A1(n479), .A2(n573), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT101), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n482), .ZN(n508) );
  NOR2_X1 U543 ( .A1(n483), .A2(n508), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n510), .A2(n492), .ZN(n486) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n485) );
  XNOR2_X1 U546 ( .A(G29GAT), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U547 ( .A1(n492), .A2(n513), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n490) );
  NAND2_X1 U550 ( .A1(n492), .A2(n522), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n494) );
  NAND2_X1 U554 ( .A1(n492), .A2(n525), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(n495), .ZN(G1331GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n499) );
  INV_X1 U558 ( .A(n556), .ZN(n528) );
  NAND2_X1 U559 ( .A1(n528), .A2(n565), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT106), .ZN(n509) );
  NOR2_X1 U561 ( .A1(n509), .A2(n497), .ZN(n503) );
  NAND2_X1 U562 ( .A1(n510), .A2(n503), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n513), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U567 ( .A1(n503), .A2(n522), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U570 ( .A1(n503), .A2(n525), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n507) );
  XOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT108), .Z(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n508), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n510), .A2(n517), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT110), .B(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  XOR2_X1 U578 ( .A(G92GAT), .B(KEYINPUT111), .Z(n515) );
  NAND2_X1 U579 ( .A1(n517), .A2(n513), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NAND2_X1 U581 ( .A1(n522), .A2(n517), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U583 ( .A1(n525), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n540) );
  NAND2_X1 U587 ( .A1(n540), .A2(n522), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT115), .B(n523), .Z(n524) );
  NOR2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n526), .A2(n536), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U593 ( .A1(n536), .A2(n528), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(KEYINPUT117), .ZN(n534) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n532) );
  NAND2_X1 U597 ( .A1(n536), .A2(n560), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n538) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n540), .A2(n563), .ZN(n549) );
  NOR2_X1 U605 ( .A1(n565), .A2(n549), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  NOR2_X1 U608 ( .A1(n556), .A2(n549), .ZN(n547) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n544) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(KEYINPUT120), .B(n545), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n573), .A2(n549), .ZN(n548) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n565), .A2(n559), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G169GAT), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT123), .ZN(G1348GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n555) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n556), .A2(n559), .ZN(n557) );
  XOR2_X1 U625 ( .A(n558), .B(n557), .Z(G1349GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n577) );
  NOR2_X1 U630 ( .A1(n565), .A2(n577), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n577), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n577), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n576) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

