//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT66), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT68), .Z(G261));
  AOI22_X1  g032(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G137), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n459), .B2(new_n460), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n473), .B2(G2105), .ZN(G160));
  NOR2_X1   g049(.A1(new_n459), .A2(new_n460), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(new_n476), .B2(G112), .ZN(new_n480));
  INV_X1    g055(.A(G100), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(new_n476), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n475), .A2(G2105), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n479), .B(new_n483), .C1(G136), .C2(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n464), .A2(new_n470), .A3(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n467), .B2(new_n469), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n476), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n467), .B2(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n466), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n488), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n501), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n512), .A2(new_n514), .A3(G543), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n512), .A2(new_n514), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n511), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(new_n515), .B(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n508), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n525), .B(new_n530), .C1(new_n531), .C2(new_n519), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  INV_X1    g108(.A(new_n519), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(G90), .B1(G52), .B2(new_n524), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n506), .A2(new_n507), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  INV_X1    g112(.A(G77), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n538), .B2(new_n504), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT73), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  OAI221_X1 g116(.A(new_n541), .B1(new_n538), .B2(new_n504), .C1(new_n536), .C2(new_n537), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(G651), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n535), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n524), .A2(G43), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT75), .B(G81), .Z(new_n547));
  NAND3_X1  g122(.A1(new_n508), .A2(new_n518), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n506), .A2(G56), .A3(new_n507), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n510), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n546), .B(new_n548), .C1(KEYINPUT74), .C2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(G860), .A3(new_n554), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n506), .A2(new_n560), .A3(new_n507), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n560), .B1(new_n506), .B2(new_n507), .ZN(new_n562));
  OAI21_X1  g137(.A(G65), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n510), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n566));
  AND2_X1   g141(.A1(G53), .A2(G543), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n518), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n566), .B1(new_n518), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n508), .A2(G91), .A3(new_n518), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n565), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  OAI21_X1  g148(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n508), .A2(G87), .A3(new_n518), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n516), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND4_X1  g152(.A1(new_n518), .A2(new_n506), .A3(G86), .A4(new_n507), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n515), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n506), .A2(G61), .A3(new_n507), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n510), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n510), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n518), .A2(KEYINPUT72), .A3(G543), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n515), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n519), .A2(new_n588), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G290));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(G301), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n508), .A2(G92), .A3(new_n518), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n508), .A2(KEYINPUT10), .A3(G92), .A4(new_n518), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n524), .A2(G54), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n506), .A2(new_n560), .A3(new_n507), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n603), .B(new_n604), .C1(new_n608), .C2(new_n510), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT78), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(new_n597), .ZN(G284));
  AOI21_X1  g186(.A(new_n598), .B1(new_n610), .B2(new_n597), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n572), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n572), .B2(G868), .ZN(G280));
  XOR2_X1   g190(.A(KEYINPUT79), .B(G559), .Z(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(G860), .B2(new_n616), .ZN(G148));
  NAND2_X1  g192(.A1(new_n553), .A2(new_n554), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n616), .ZN(new_n619));
  MUX2_X1   g194(.A(new_n618), .B(new_n619), .S(G868), .Z(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g196(.A1(new_n464), .A2(new_n470), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n622), .A2(new_n466), .A3(G2105), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n623), .B(new_n624), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n484), .A2(G135), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT81), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n477), .A2(G123), .ZN(new_n631));
  NOR2_X1   g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(new_n476), .B2(G111), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G2096), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n627), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT82), .Z(G156));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT14), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n644), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n644), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n653), .A3(G14), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT85), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT84), .Z(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  INV_X1    g242(.A(new_n657), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n662), .B1(new_n668), .B2(new_n661), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n635), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(G2096), .ZN(new_n674));
  INV_X1    g249(.A(G2100), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n688), .B(new_n691), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT87), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  NAND2_X1  g274(.A1(G303), .A2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(new_n701), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n701), .B2(G23), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n704), .A2(new_n705), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n703), .A2(G1971), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(G305), .A2(G16), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT32), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n701), .A2(G6), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n715), .B1(new_n714), .B2(new_n716), .ZN(new_n718));
  OAI21_X1  g293(.A(G1981), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT34), .ZN(new_n720));
  OR3_X1    g295(.A1(new_n717), .A2(new_n718), .A3(G1981), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n719), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n708), .A2(new_n709), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n703), .B2(G1971), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n724), .A2(new_n721), .A3(new_n710), .A4(new_n719), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n701), .B1(G290), .B2(KEYINPUT90), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(KEYINPUT90), .B2(G290), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n701), .A2(G24), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n728), .A2(new_n690), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n690), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n484), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n477), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT89), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT89), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  MUX2_X1   g316(.A(G25), .B(new_n736), .S(new_n741), .Z(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT35), .B(G1991), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n730), .A2(new_n731), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n722), .A2(new_n726), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n722), .A2(new_n726), .A3(new_n748), .A4(new_n745), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n737), .A2(G33), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT93), .B(KEYINPUT25), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n484), .A2(G139), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT95), .ZN(new_n758));
  INV_X1    g333(.A(new_n622), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n759), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(new_n476), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n751), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n701), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n572), .B2(new_n701), .ZN(new_n767));
  INV_X1    g342(.A(G1956), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n741), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n741), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT29), .B(G2090), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n466), .A2(G2105), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n477), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT26), .Z(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n737), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n737), .B2(G32), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n771), .A2(new_n772), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n771), .B2(new_n772), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n741), .A2(G27), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n741), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G2078), .Z(new_n787));
  INV_X1    g362(.A(G160), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n740), .B1(new_n789), .B2(G34), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT96), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(G34), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n788), .A2(new_n737), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n787), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n701), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n701), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1966), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT31), .B(G11), .Z(new_n803));
  INV_X1    g378(.A(KEYINPUT30), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n737), .B1(new_n804), .B2(G28), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT97), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(KEYINPUT97), .B1(new_n804), .B2(G28), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n808), .B1(new_n634), .B2(new_n740), .C1(new_n781), .C2(new_n782), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n784), .A2(new_n799), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n701), .A2(G5), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G171), .B2(new_n701), .ZN(new_n812));
  INV_X1    g387(.A(G1961), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n764), .A2(new_n769), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n740), .A2(G26), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT91), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n484), .A2(G140), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n477), .A2(G128), .ZN(new_n821));
  NOR2_X1   g396(.A1(G104), .A2(G2105), .ZN(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(new_n476), .B2(G116), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n820), .B(new_n821), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(new_n818), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n819), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G2067), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n701), .A2(G19), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n618), .B2(G16), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(G1341), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(G1341), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n610), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G4), .B2(G16), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G1348), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(G1348), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT92), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(new_n833), .C1(new_n836), .C2(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n815), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n750), .A2(new_n842), .ZN(G311));
  AND3_X1   g418(.A1(new_n750), .A2(new_n842), .A3(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT98), .B1(new_n750), .B2(new_n842), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(G150));
  NAND3_X1  g421(.A1(new_n508), .A2(G93), .A3(new_n518), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n589), .A2(G55), .A3(new_n591), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n506), .A2(G67), .A3(new_n507), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n510), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G860), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n849), .A2(new_n852), .ZN(new_n857));
  INV_X1    g432(.A(new_n554), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n552), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n546), .A2(new_n548), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n853), .A2(new_n860), .A3(new_n554), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n610), .A2(G559), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n610), .B2(G559), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n859), .A2(new_n862), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n854), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(new_n872), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n870), .B2(new_n866), .ZN(new_n876));
  OAI21_X1  g451(.A(KEYINPUT39), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT100), .B(KEYINPUT39), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n874), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI211_X1 g458(.A(KEYINPUT101), .B(new_n874), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n856), .B1(new_n883), .B2(new_n884), .ZN(G145));
  XNOR2_X1  g460(.A(new_n634), .B(new_n788), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(G162), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n778), .B(new_n824), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n758), .A2(new_n499), .A3(new_n761), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n499), .B1(new_n758), .B2(new_n761), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n477), .A2(G130), .ZN(new_n895));
  NOR2_X1   g470(.A1(G106), .A2(G2105), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G142), .B2(new_n484), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n736), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n625), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n891), .A2(new_n892), .A3(new_n889), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n894), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n905), .B2(new_n893), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n887), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  OAI211_X1 g483(.A(KEYINPUT102), .B(new_n902), .C1(new_n894), .C2(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n901), .A3(new_n893), .ZN(new_n910));
  INV_X1    g485(.A(new_n887), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n906), .A2(KEYINPUT102), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n907), .B(new_n908), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g490(.A(new_n619), .B(new_n863), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n609), .A2(new_n572), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n609), .A2(new_n572), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT41), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n920));
  OR3_X1    g495(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  XNOR2_X1  g497(.A(G303), .B(new_n595), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n706), .B(KEYINPUT103), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n924), .A2(G305), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(G305), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n924), .A2(G305), .ZN(new_n928));
  XNOR2_X1  g503(.A(G290), .B(G303), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(G305), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT42), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n922), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n921), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n933), .A2(new_n922), .A3(new_n934), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n857), .A2(new_n597), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(G331));
  NAND2_X1  g519(.A1(new_n917), .A2(new_n918), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n535), .A2(new_n543), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n535), .B2(new_n543), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n948), .A2(new_n949), .A3(G168), .ZN(new_n950));
  NAND2_X1  g525(.A1(G301), .A2(KEYINPUT105), .ZN(new_n951));
  AOI21_X1  g526(.A(G286), .B1(new_n951), .B2(new_n947), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n950), .A2(new_n952), .A3(new_n863), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(G286), .A3(new_n947), .ZN(new_n954));
  OAI21_X1  g529(.A(G168), .B1(new_n948), .B2(new_n949), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n871), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n945), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n863), .B1(new_n950), .B2(new_n952), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n955), .A2(new_n871), .A3(new_n954), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n958), .B(new_n959), .C1(new_n920), .C2(new_n919), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n932), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n932), .A2(new_n957), .A3(new_n960), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n963), .A2(new_n908), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(KEYINPUT106), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n963), .A2(new_n971), .A3(new_n908), .A4(new_n964), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT43), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n965), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n967), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n965), .B2(KEYINPUT106), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n970), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n968), .B1(new_n977), .B2(new_n979), .ZN(G397));
  INV_X1    g555(.A(G1384), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n486), .A2(new_n487), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n493), .A2(new_n498), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT108), .B(G40), .Z(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(G160), .A2(KEYINPUT109), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n473), .A2(G2105), .ZN(new_n990));
  INV_X1    g565(.A(new_n463), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n988), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n986), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n995), .A2(G1996), .A3(new_n778), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT110), .ZN(new_n997));
  INV_X1    g572(.A(G2067), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n824), .B(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(G1996), .B2(new_n778), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n997), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n995), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n736), .B(new_n743), .Z(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n595), .B(new_n690), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n995), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n499), .A2(new_n1008), .A3(new_n981), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT109), .B1(G160), .B2(new_n988), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n476), .B1(new_n471), .B2(new_n472), .ZN(new_n1011));
  NOR4_X1   g586(.A1(new_n1011), .A2(new_n993), .A3(new_n463), .A4(new_n987), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n1015));
  OAI211_X1 g590(.A(new_n986), .B(new_n1015), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT56), .B(G2072), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI22_X1  g593(.A1(new_n1014), .A2(G1956), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n565), .B2(new_n571), .ZN(new_n1024));
  INV_X1    g599(.A(G65), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n605), .B2(new_n606), .ZN(new_n1026));
  INV_X1    g601(.A(new_n564), .ZN(new_n1027));
  OAI21_X1  g602(.A(G651), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n571), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(KEYINPUT120), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n570), .A2(KEYINPUT119), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n568), .B2(new_n569), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1022), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n572), .A2(KEYINPUT57), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1020), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT121), .B(new_n1038), .C1(new_n1041), .C2(new_n1022), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1019), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1348), .ZN(new_n1044));
  INV_X1    g619(.A(new_n984), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(new_n998), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1044), .A2(new_n1013), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n610), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1040), .A2(new_n1042), .A3(new_n1019), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1040), .A2(new_n1042), .A3(new_n1019), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1055), .A2(new_n1043), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1019), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n565), .A2(new_n1023), .A3(new_n571), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1036), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1021), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT121), .B1(new_n1062), .B2(new_n1038), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1042), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT61), .B1(new_n1065), .B2(new_n1053), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1057), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1069));
  XOR2_X1   g644(.A(new_n1069), .B(KEYINPUT126), .Z(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n994), .A2(new_n989), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT4), .B(G138), .C1(new_n459), .C2(new_n460), .ZN(new_n1073));
  AOI21_X1  g648(.A(G2105), .B1(new_n1073), .B2(new_n491), .ZN(new_n1074));
  OAI21_X1  g649(.A(G126), .B1(new_n459), .B2(new_n460), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n487), .B1(G114), .B2(G2104), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n476), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  AOI211_X1 g653(.A(new_n985), .B(G1384), .C1(new_n1078), .C2(new_n488), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n499), .B2(new_n981), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT123), .B(G1996), .Z(new_n1082));
  NAND3_X1  g657(.A1(new_n1072), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1045), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(new_n1086), .A3(KEYINPUT124), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT124), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n618), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1071), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1090), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1088), .A2(new_n618), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1092), .B(new_n1070), .C1(new_n1093), .C2(new_n1087), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1050), .A2(KEYINPUT60), .A3(new_n610), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1048), .A2(KEYINPUT60), .A3(new_n1049), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT60), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(new_n1051), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1091), .A2(new_n1094), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1054), .B1(new_n1067), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1013), .A2(new_n813), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2078), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1072), .A2(new_n1081), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1072), .A2(new_n1081), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G2078), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1102), .B(new_n1105), .C1(new_n1109), .C2(KEYINPUT53), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1101), .B1(new_n1111), .B2(G301), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1081), .A2(G40), .A3(G160), .A4(new_n1104), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1102), .C1(new_n1109), .C2(KEYINPUT53), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1112), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1106), .A2(new_n705), .A3(new_n1108), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT112), .B(G2090), .Z(new_n1121));
  NAND2_X1  g696(.A1(new_n1014), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G303), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT55), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(G8), .A3(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n580), .A2(new_n583), .A3(G1981), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(G1981), .B1(new_n580), .B2(new_n583), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(KEYINPUT49), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1130), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1132), .B1(new_n1135), .B2(new_n1128), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1134), .A2(new_n1136), .A3(new_n1084), .A4(G8), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n706), .A2(G1976), .ZN(new_n1138));
  INV_X1    g713(.A(G1976), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT52), .B1(G288), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1084), .A2(G8), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1084), .A2(G8), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1138), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(KEYINPUT52), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1127), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1126), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1123), .A2(KEYINPUT115), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1120), .A2(new_n1149), .A3(new_n1122), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1148), .A2(G8), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1146), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1110), .A2(G171), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1114), .A2(G171), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1101), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT116), .B1(new_n1013), .B2(G2084), .ZN(new_n1156));
  AOI211_X1 g731(.A(KEYINPUT50), .B(G1384), .C1(new_n1078), .C2(new_n488), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1008), .B1(new_n499), .B2(new_n981), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1072), .A2(new_n1159), .A3(new_n1160), .A4(new_n796), .ZN(new_n1161));
  INV_X1    g736(.A(G1966), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1016), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1156), .A2(G168), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1072), .A2(new_n1159), .A3(new_n796), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1166), .A2(KEYINPUT116), .B1(new_n1162), .B2(new_n1016), .ZN(new_n1167));
  AOI21_X1  g742(.A(G168), .B1(new_n1167), .B2(new_n1161), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT51), .B1(new_n1164), .B2(G8), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1119), .A2(new_n1152), .A3(new_n1155), .A4(new_n1171), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1100), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1170), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1176), .B(KEYINPUT62), .C1(new_n1168), .C2(new_n1165), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1152), .A2(new_n1153), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1127), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G288), .A2(G1976), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT114), .Z(new_n1182));
  OAI21_X1  g757(.A(new_n1129), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  AOI22_X1  g758(.A1(new_n1179), .A2(new_n1145), .B1(new_n1143), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(G168), .A2(G8), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1185), .B1(new_n1167), .B2(new_n1161), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n1152), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1123), .A2(G8), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1189), .B2(new_n1147), .ZN(new_n1190));
  AOI211_X1 g765(.A(KEYINPUT117), .B(new_n1126), .C1(new_n1123), .C2(G8), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1145), .A2(KEYINPUT63), .A3(new_n1186), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1178), .B(new_n1184), .C1(new_n1187), .C2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1006), .B1(new_n1173), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1002), .A2(G1996), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT46), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n999), .A2(new_n779), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1196), .A2(new_n1197), .B1(new_n995), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1200));
  XOR2_X1   g775(.A(new_n1200), .B(KEYINPUT47), .Z(new_n1201));
  NAND3_X1  g776(.A1(new_n995), .A2(new_n690), .A3(new_n595), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1202), .B(KEYINPUT48), .Z(new_n1203));
  NOR2_X1   g778(.A1(new_n1004), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n736), .A2(new_n743), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1001), .A2(new_n1205), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n824), .A2(G2067), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1002), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g783(.A1(new_n1201), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1195), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g785(.A1(new_n654), .A2(G319), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n697), .B2(new_n698), .ZN(new_n1213));
  AND3_X1   g787(.A1(new_n673), .A2(new_n676), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n1214), .A2(new_n914), .A3(new_n966), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


