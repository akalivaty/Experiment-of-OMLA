

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(G2104), .A2(n523), .ZN(n890) );
  XNOR2_X1 U554 ( .A(n533), .B(KEYINPUT66), .ZN(n534) );
  AND2_X1 U555 ( .A1(n523), .A2(G2104), .ZN(n885) );
  NOR2_X1 U556 ( .A1(n539), .A2(n538), .ZN(G160) );
  BUF_X1 U557 ( .A(n703), .Z(n720) );
  XNOR2_X1 U558 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n685) );
  XNOR2_X1 U559 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U560 ( .A(n683), .B(KEYINPUT93), .ZN(n768) );
  NOR2_X1 U561 ( .A1(G1384), .A2(G164), .ZN(n682) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n533) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n636) );
  NOR2_X1 U564 ( .A1(G651), .A2(n636), .ZN(n645) );
  XOR2_X1 U565 ( .A(KEYINPUT15), .B(n589), .Z(n976) );
  XNOR2_X1 U566 ( .A(n535), .B(n534), .ZN(n537) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n520), .Z(n886) );
  NAND2_X1 U569 ( .A1(G138), .A2(n886), .ZN(n522) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U571 ( .A1(G114), .A2(n889), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n528) );
  INV_X1 U573 ( .A(G2105), .ZN(n523) );
  NAND2_X1 U574 ( .A1(n885), .A2(G102), .ZN(n526) );
  NAND2_X1 U575 ( .A1(G126), .A2(n890), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT87), .B(n524), .Z(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X2 U578 ( .A1(n528), .A2(n527), .ZN(G164) );
  NAND2_X1 U579 ( .A1(G125), .A2(n890), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT65), .B(n529), .Z(n532) );
  NAND2_X1 U581 ( .A1(G113), .A2(n889), .ZN(n530) );
  XOR2_X1 U582 ( .A(KEYINPUT67), .B(n530), .Z(n531) );
  NAND2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n539) );
  NAND2_X1 U584 ( .A1(G101), .A2(n885), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G137), .A2(n886), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n644) );
  NAND2_X1 U588 ( .A1(n644), .A2(G91), .ZN(n542) );
  INV_X1 U589 ( .A(G651), .ZN(n543) );
  OR2_X1 U590 ( .A1(n543), .A2(n636), .ZN(n540) );
  XOR2_X2 U591 ( .A(KEYINPUT68), .B(n540), .Z(n643) );
  NAND2_X1 U592 ( .A1(G78), .A2(n643), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n542), .A2(n541), .ZN(n548) );
  NOR2_X1 U594 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n544), .Z(n650) );
  NAND2_X1 U596 ( .A1(G65), .A2(n650), .ZN(n546) );
  NAND2_X1 U597 ( .A1(G53), .A2(n645), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  OR2_X1 U599 ( .A1(n548), .A2(n547), .ZN(G299) );
  NAND2_X1 U600 ( .A1(G64), .A2(n650), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G52), .A2(n645), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U603 ( .A1(n644), .A2(G90), .ZN(n552) );
  NAND2_X1 U604 ( .A1(G77), .A2(n643), .ZN(n551) );
  NAND2_X1 U605 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U606 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  XNOR2_X1 U607 ( .A(KEYINPUT69), .B(n554), .ZN(n555) );
  NOR2_X1 U608 ( .A1(n556), .A2(n555), .ZN(G171) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G132), .ZN(G219) );
  NAND2_X1 U612 ( .A1(G63), .A2(n650), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G51), .A2(n645), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(KEYINPUT6), .B(n559), .ZN(n565) );
  NAND2_X1 U616 ( .A1(n644), .A2(G89), .ZN(n560) );
  XNOR2_X1 U617 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G76), .A2(n643), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U620 ( .A(n563), .B(KEYINPUT5), .Z(n564) );
  NOR2_X1 U621 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U622 ( .A(KEYINPUT75), .B(n566), .Z(n567) );
  XOR2_X1 U623 ( .A(KEYINPUT7), .B(n567), .Z(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U626 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n833) );
  NAND2_X1 U628 ( .A1(n833), .A2(G567), .ZN(n569) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U630 ( .A1(n650), .A2(G56), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n570), .Z(n577) );
  NAND2_X1 U632 ( .A1(G68), .A2(n643), .ZN(n571) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n644), .A2(G81), .ZN(n572) );
  XOR2_X1 U635 ( .A(KEYINPUT12), .B(n572), .Z(n573) );
  NOR2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT13), .ZN(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT72), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G43), .A2(n645), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n974) );
  INV_X1 U642 ( .A(G860), .ZN(n595) );
  OR2_X1 U643 ( .A1(n974), .A2(n595), .ZN(G153) );
  INV_X1 U644 ( .A(G868), .ZN(n665) );
  NOR2_X1 U645 ( .A1(n665), .A2(G171), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT73), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n645), .A2(G54), .ZN(n588) );
  NAND2_X1 U648 ( .A1(G92), .A2(n644), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G66), .A2(n650), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n643), .A2(G79), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT74), .B(n584), .Z(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n665), .A2(n976), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(G284) );
  NOR2_X1 U657 ( .A1(G286), .A2(n665), .ZN(n593) );
  NOR2_X1 U658 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(KEYINPUT76), .B(n594), .ZN(G297) );
  NAND2_X1 U661 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U662 ( .A(n976), .ZN(n904) );
  NAND2_X1 U663 ( .A1(n596), .A2(n904), .ZN(n597) );
  XNOR2_X1 U664 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U665 ( .A1(G868), .A2(n974), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n904), .A2(G868), .ZN(n598) );
  NOR2_X1 U667 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U668 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U669 ( .A1(G99), .A2(n885), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G111), .A2(n889), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n603), .B(KEYINPUT77), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G135), .A2(n886), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n890), .A2(G123), .ZN(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT18), .B(n606), .Z(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n926) );
  XNOR2_X1 U678 ( .A(n926), .B(G2096), .ZN(n610) );
  INV_X1 U679 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U681 ( .A1(G559), .A2(n904), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(n974), .ZN(n661) );
  NOR2_X1 U683 ( .A1(n661), .A2(G860), .ZN(n621) );
  NAND2_X1 U684 ( .A1(G93), .A2(n644), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n612), .B(KEYINPUT78), .ZN(n619) );
  NAND2_X1 U686 ( .A1(G67), .A2(n650), .ZN(n614) );
  NAND2_X1 U687 ( .A1(G55), .A2(n645), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U689 ( .A1(G80), .A2(n643), .ZN(n615) );
  XNOR2_X1 U690 ( .A(KEYINPUT79), .B(n615), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n664) );
  XOR2_X1 U693 ( .A(n664), .B(KEYINPUT80), .Z(n620) );
  XNOR2_X1 U694 ( .A(n621), .B(n620), .ZN(G145) );
  NAND2_X1 U695 ( .A1(n644), .A2(G88), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G75), .A2(n643), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G62), .A2(n650), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G50), .A2(n645), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U701 ( .A1(n627), .A2(n626), .ZN(G166) );
  NAND2_X1 U702 ( .A1(n643), .A2(G73), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U704 ( .A1(G61), .A2(n650), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G48), .A2(n645), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U707 ( .A1(n644), .A2(G86), .ZN(n631) );
  XOR2_X1 U708 ( .A(KEYINPUT82), .B(n631), .Z(n632) );
  NOR2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U711 ( .A1(n636), .A2(G87), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G49), .A2(n645), .ZN(n638) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n650), .A2(n639), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U717 ( .A(KEYINPUT81), .B(n642), .Z(G288) );
  AND2_X1 U718 ( .A1(G72), .A2(n643), .ZN(n649) );
  NAND2_X1 U719 ( .A1(G85), .A2(n644), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G47), .A2(n645), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n650), .A2(G60), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n652), .A2(n651), .ZN(G290) );
  XOR2_X1 U725 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(G166), .B(n655), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(n664), .ZN(n658) );
  XOR2_X1 U730 ( .A(G305), .B(G288), .Z(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(G290), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G299), .ZN(n903) );
  XNOR2_X1 U734 ( .A(KEYINPUT86), .B(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n903), .B(n662), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U743 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U745 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n672) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U748 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U749 ( .A1(G96), .A2(n674), .ZN(n837) );
  NAND2_X1 U750 ( .A1(n837), .A2(G2106), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U752 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(G108), .A2(n676), .ZN(n838) );
  NAND2_X1 U754 ( .A1(n838), .A2(G567), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n839) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U757 ( .A1(n839), .A2(n679), .ZN(n836) );
  NAND2_X1 U758 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  NAND2_X1 U760 ( .A1(G288), .A2(G1976), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT102), .B(n680), .Z(n982) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n801) );
  INV_X1 U763 ( .A(KEYINPUT64), .ZN(n681) );
  XNOR2_X1 U764 ( .A(n682), .B(n681), .ZN(n799) );
  NOR2_X1 U765 ( .A1(n801), .A2(n799), .ZN(n703) );
  INV_X2 U766 ( .A(n703), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n719), .A2(G8), .ZN(n683) );
  INV_X1 U768 ( .A(n768), .ZN(n774) );
  NOR2_X1 U769 ( .A1(G1966), .A2(n774), .ZN(n748) );
  NOR2_X1 U770 ( .A1(G2084), .A2(n719), .ZN(n744) );
  NOR2_X1 U771 ( .A1(n748), .A2(n744), .ZN(n684) );
  NAND2_X1 U772 ( .A1(G8), .A2(n684), .ZN(n686) );
  NOR2_X1 U773 ( .A1(G168), .A2(n687), .ZN(n692) );
  AND2_X1 U774 ( .A1(n719), .A2(G1961), .ZN(n690) );
  XNOR2_X1 U775 ( .A(G2078), .B(KEYINPUT94), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n688), .B(KEYINPUT25), .ZN(n960) );
  NOR2_X1 U777 ( .A1(n960), .A2(n719), .ZN(n689) );
  NOR2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n733) );
  NOR2_X1 U779 ( .A1(G171), .A2(n733), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U781 ( .A(KEYINPUT31), .B(n693), .Z(n746) );
  INV_X1 U782 ( .A(G8), .ZN(n700) );
  NOR2_X1 U783 ( .A1(G1971), .A2(n774), .ZN(n694) );
  XOR2_X1 U784 ( .A(KEYINPUT99), .B(n694), .Z(n696) );
  NOR2_X1 U785 ( .A1(G2090), .A2(n719), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U787 ( .A(n697), .B(KEYINPUT100), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n698), .A2(G303), .ZN(n699) );
  OR2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n738) );
  XOR2_X1 U790 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n707) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n707), .ZN(n702) );
  NAND2_X1 U792 ( .A1(G2067), .A2(n976), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n704), .A2(n720), .ZN(n714) );
  INV_X1 U795 ( .A(G1341), .ZN(n1013) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n976), .ZN(n705) );
  NAND2_X1 U797 ( .A1(n1013), .A2(n705), .ZN(n706) );
  NAND2_X1 U798 ( .A1(n706), .A2(n719), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n720), .A2(G1996), .ZN(n709) );
  INV_X1 U800 ( .A(n707), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U803 ( .A1(n974), .A2(n712), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n727) );
  NAND2_X1 U805 ( .A1(n720), .A2(G2072), .ZN(n715) );
  XOR2_X1 U806 ( .A(KEYINPUT27), .B(n715), .Z(n717) );
  NAND2_X1 U807 ( .A1(G1956), .A2(n719), .ZN(n716) );
  NAND2_X1 U808 ( .A1(n717), .A2(n716), .ZN(n728) );
  NOR2_X1 U809 ( .A1(G299), .A2(n728), .ZN(n718) );
  XNOR2_X1 U810 ( .A(n718), .B(KEYINPUT96), .ZN(n725) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n719), .ZN(n722) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n720), .ZN(n721) );
  NAND2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n976), .A2(n723), .ZN(n724) );
  NOR2_X1 U815 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n731) );
  NAND2_X1 U817 ( .A1(G299), .A2(n728), .ZN(n729) );
  XNOR2_X1 U818 ( .A(n729), .B(KEYINPUT28), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U820 ( .A(n732), .B(KEYINPUT29), .ZN(n735) );
  AND2_X1 U821 ( .A1(G171), .A2(n733), .ZN(n734) );
  NOR2_X1 U822 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U823 ( .A(KEYINPUT97), .B(n736), .ZN(n745) );
  AND2_X1 U824 ( .A1(n738), .A2(n745), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n746), .A2(n737), .ZN(n742) );
  INV_X1 U826 ( .A(n738), .ZN(n740) );
  AND2_X1 U827 ( .A1(G286), .A2(G8), .ZN(n739) );
  OR2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U830 ( .A(KEYINPUT32), .B(n743), .ZN(n752) );
  NAND2_X1 U831 ( .A1(G8), .A2(n744), .ZN(n750) );
  AND2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U834 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U835 ( .A1(n752), .A2(n751), .ZN(n772) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U838 ( .A1(n756), .A2(n753), .ZN(n978) );
  NAND2_X1 U839 ( .A1(n772), .A2(n978), .ZN(n754) );
  XNOR2_X1 U840 ( .A(n754), .B(KEYINPUT101), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n982), .A2(n755), .ZN(n762) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n764) );
  NAND2_X1 U843 ( .A1(n768), .A2(n756), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n764), .A2(n757), .ZN(n758) );
  XNOR2_X1 U845 ( .A(n758), .B(KEYINPUT103), .ZN(n763) );
  AND2_X1 U846 ( .A1(n768), .A2(n763), .ZN(n760) );
  XNOR2_X1 U847 ( .A(G1981), .B(G305), .ZN(n996) );
  INV_X1 U848 ( .A(n996), .ZN(n759) );
  AND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n780) );
  INV_X1 U851 ( .A(n763), .ZN(n765) );
  OR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n996), .A2(n766), .ZN(n778) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XNOR2_X1 U855 ( .A(KEYINPUT24), .B(n767), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n776) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U863 ( .A1(n780), .A2(n779), .ZN(n806) );
  NAND2_X1 U864 ( .A1(G105), .A2(n885), .ZN(n781) );
  XNOR2_X1 U865 ( .A(n781), .B(KEYINPUT38), .ZN(n788) );
  NAND2_X1 U866 ( .A1(G117), .A2(n889), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G141), .A2(n886), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n890), .A2(G129), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT90), .B(n784), .Z(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n897) );
  NAND2_X1 U873 ( .A1(G1996), .A2(n897), .ZN(n789) );
  XOR2_X1 U874 ( .A(KEYINPUT91), .B(n789), .Z(n798) );
  NAND2_X1 U875 ( .A1(G95), .A2(n885), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G107), .A2(n889), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G119), .A2(n890), .ZN(n792) );
  XNOR2_X1 U879 ( .A(KEYINPUT89), .B(n792), .ZN(n793) );
  NOR2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U881 ( .A1(n886), .A2(G131), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n868) );
  NAND2_X1 U883 ( .A1(G1991), .A2(n868), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n927) );
  INV_X1 U885 ( .A(n799), .ZN(n800) );
  NOR2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n829) );
  NAND2_X1 U887 ( .A1(n927), .A2(n829), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n802), .B(KEYINPUT92), .ZN(n804) );
  XNOR2_X1 U889 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U890 ( .A1(n980), .A2(n829), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n817) );
  NAND2_X1 U893 ( .A1(n885), .A2(G104), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(KEYINPUT88), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G140), .A2(n886), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n810), .ZN(n815) );
  NAND2_X1 U898 ( .A1(G116), .A2(n889), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G128), .A2(n890), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n813), .Z(n814) );
  NOR2_X1 U902 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U903 ( .A(KEYINPUT36), .B(n816), .Z(n879) );
  XOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .Z(n825) );
  AND2_X1 U905 ( .A1(n879), .A2(n825), .ZN(n936) );
  NAND2_X1 U906 ( .A1(n829), .A2(n936), .ZN(n823) );
  NAND2_X1 U907 ( .A1(n817), .A2(n823), .ZN(n831) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n868), .ZN(n928) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U910 ( .A1(n928), .A2(n818), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n927), .A2(n819), .ZN(n821) );
  NOR2_X1 U912 ( .A1(n897), .A2(G1996), .ZN(n820) );
  XNOR2_X1 U913 ( .A(n820), .B(KEYINPUT104), .ZN(n938) );
  NOR2_X1 U914 ( .A1(n821), .A2(n938), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n879), .A2(n825), .ZN(n826) );
  XNOR2_X1 U918 ( .A(KEYINPUT105), .B(n826), .ZN(n944) );
  NAND2_X1 U919 ( .A1(n827), .A2(n944), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U922 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U925 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U929 ( .A(G120), .ZN(G236) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  INV_X1 U931 ( .A(G69), .ZN(G235) );
  NOR2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n839), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2090), .Z(n841) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U938 ( .A(n842), .B(G2100), .Z(n844) );
  XNOR2_X1 U939 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n846) );
  XNOR2_X1 U942 ( .A(KEYINPUT107), .B(G2678), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U945 ( .A(KEYINPUT109), .B(G1956), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U948 ( .A(n851), .B(KEYINPUT108), .Z(n853) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1971), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1961), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U955 ( .A(G2474), .B(KEYINPUT41), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U957 ( .A1(n886), .A2(G136), .ZN(n866) );
  NAND2_X1 U958 ( .A1(G100), .A2(n885), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G112), .A2(n889), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n890), .A2(G124), .ZN(n862) );
  XOR2_X1 U962 ( .A(KEYINPUT44), .B(n862), .Z(n863) );
  NOR2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT110), .B(n867), .Z(G162) );
  XNOR2_X1 U966 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n868), .B(KEYINPUT112), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n884) );
  NAND2_X1 U969 ( .A1(G106), .A2(n885), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G142), .A2(n886), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT45), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G118), .A2(n889), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G130), .A2(n890), .ZN(n876) );
  XNOR2_X1 U976 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  NOR2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n880) );
  XOR2_X1 U978 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U979 ( .A(G160), .B(G164), .ZN(n881) );
  XNOR2_X1 U980 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n884), .B(n883), .ZN(n899) );
  NAND2_X1 U982 ( .A1(G103), .A2(n885), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G139), .A2(n886), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U985 ( .A1(G115), .A2(n889), .ZN(n892) );
  NAND2_X1 U986 ( .A1(G127), .A2(n890), .ZN(n891) );
  NAND2_X1 U987 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U988 ( .A(KEYINPUT47), .B(n893), .ZN(n894) );
  XNOR2_X1 U989 ( .A(KEYINPUT113), .B(n894), .ZN(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n931) );
  XNOR2_X1 U991 ( .A(n897), .B(n931), .ZN(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n926), .B(n900), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(G162), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U996 ( .A(n903), .B(G286), .Z(n906) );
  XNOR2_X1 U997 ( .A(G171), .B(n904), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U999 ( .A(n907), .B(n974), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n908), .ZN(G397) );
  XOR2_X1 U1001 ( .A(KEYINPUT106), .B(G2446), .Z(n910) );
  XNOR2_X1 U1002 ( .A(G2443), .B(G2454), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1004 ( .A(n911), .B(G2451), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G1341), .B(G1348), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n917) );
  XOR2_X1 U1007 ( .A(G2435), .B(G2427), .Z(n915) );
  XNOR2_X1 U1008 ( .A(G2430), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1010 ( .A(n917), .B(n916), .Z(n918) );
  NAND2_X1 U1011 ( .A1(G14), .A2(n918), .ZN(n924) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n924), .ZN(n921) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1017 ( .A1(n923), .A2(n922), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  INV_X1 U1020 ( .A(n924), .ZN(G401) );
  INV_X1 U1021 ( .A(G171), .ZN(G301) );
  INV_X1 U1022 ( .A(KEYINPUT55), .ZN(n949) );
  XOR2_X1 U1023 ( .A(KEYINPUT52), .B(KEYINPUT114), .Z(n947) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n925) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n943) );
  XOR2_X1 U1028 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n941) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1039 ( .A(n947), .B(n946), .ZN(n948) );
  NAND2_X1 U1040 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1041 ( .A1(n950), .A2(G29), .ZN(n1006) );
  XNOR2_X1 U1042 ( .A(KEYINPUT115), .B(G2072), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(n951), .B(G33), .ZN(n959) );
  XNOR2_X1 U1044 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1045 ( .A(G25), .B(G1991), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(G28), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(KEYINPUT116), .B(G1996), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G32), .B(n955), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1052 ( .A(n960), .B(G27), .Z(n961) );
  NOR2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1054 ( .A(KEYINPUT53), .B(n963), .Z(n966) );
  XOR2_X1 U1055 ( .A(G34), .B(KEYINPUT54), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G2084), .B(n964), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G35), .B(G2090), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1060 ( .A(KEYINPUT55), .B(n969), .Z(n970) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n970), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(KEYINPUT117), .B(n971), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n973), .B(KEYINPUT118), .ZN(n1004) );
  XOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .Z(n1002) );
  XNOR2_X1 U1066 ( .A(G1341), .B(KEYINPUT122), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n993) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT120), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(n976), .ZN(n990) );
  INV_X1 U1070 ( .A(n978), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G299), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(G1971), .A2(G303), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G301), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n991), .B(KEYINPUT121), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G168), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n994), .B(KEYINPUT119), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n997), .Z(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(n1000), .B(KEYINPUT123), .ZN(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1034) );
  XOR2_X1 U1091 ( .A(G1986), .B(G24), .Z(n1010) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1012), .B(n1011), .ZN(n1028) );
  XNOR2_X1 U1098 ( .A(G19), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G1956), .B(G20), .ZN(n1015) );
  XNOR2_X1 U1100 ( .A(G6), .B(G1981), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT124), .B(n1018), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT59), .B(G1348), .Z(n1019) );
  XNOR2_X1 U1105 ( .A(G4), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT60), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1023), .B(KEYINPUT125), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(G21), .B(G1966), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(G5), .B(G1961), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1031), .Z(n1032) );
  NOR2_X1 U1116 ( .A1(G16), .A2(n1032), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1118 ( .A(n1035), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

