//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1161, new_n1162, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201, new_n1202, new_n1203;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n202), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n210), .B1(G97), .B2(G257), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n201), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G244), .Z(new_n220));
  OAI221_X1 g0020(.A(new_n217), .B1(new_n203), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n222), .A2(G13), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n224), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT65), .B(G107), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  XOR2_X1   g0053(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT74), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT74), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT77), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT74), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT74), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT77), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n259), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(G20), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n203), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n229), .A2(new_n261), .ZN(new_n275));
  INV_X1    g0075(.A(G159), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G58), .A2(G68), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n225), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(G20), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n255), .B1(new_n274), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n228), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n262), .A2(KEYINPUT3), .A3(new_n263), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n266), .A2(G33), .ZN(new_n286));
  AOI21_X1  g0086(.A(G20), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G68), .B1(new_n287), .B2(new_n271), .ZN(new_n288));
  AOI211_X1 g0088(.A(KEYINPUT7), .B(G20), .C1(new_n285), .C2(new_n286), .ZN(new_n289));
  OAI211_X1 g0089(.A(KEYINPUT16), .B(new_n280), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT75), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n286), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(new_n258), .B2(KEYINPUT3), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT7), .B1(new_n294), .B2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n287), .A2(new_n271), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G68), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n297), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n280), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n282), .A2(new_n284), .A3(new_n292), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n212), .A2(G1698), .ZN(new_n300));
  OR2_X1    g0100(.A1(G223), .A2(G1698), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n294), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n261), .B2(new_n208), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G1), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G41), .B2(G45), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G41), .ZN(new_n310));
  OAI211_X1 g0110(.A(G1), .B(G13), .C1(new_n261), .C2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n311), .A2(G232), .A3(new_n307), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT78), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n305), .A2(new_n309), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G190), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT8), .B(G58), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n306), .A2(G13), .A3(G20), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n284), .B1(new_n306), .B2(G20), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n314), .A2(G200), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n299), .A2(new_n316), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT17), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n292), .A2(new_n284), .A3(new_n298), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n324), .B1(new_n330), .B2(new_n282), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT17), .A3(new_n316), .A4(new_n326), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n270), .A2(new_n273), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G68), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n254), .B1(new_n334), .B2(new_n280), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n292), .A2(new_n284), .A3(new_n298), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n314), .A2(G169), .ZN(new_n338));
  INV_X1    g0138(.A(G179), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(new_n314), .ZN(new_n340));
  AND3_X1   g0140(.A1(new_n337), .A2(new_n340), .A3(KEYINPUT18), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT18), .B1(new_n337), .B2(new_n340), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n329), .B(new_n332), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT79), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G223), .A2(G1698), .ZN(new_n345));
  INV_X1    g0145(.A(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G222), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n272), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n304), .C1(G77), .C2(new_n272), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n311), .A2(new_n307), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n349), .B(new_n309), .C1(new_n212), .C2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n351), .B(KEYINPUT66), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G190), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n204), .A2(G20), .ZN(new_n355));
  INV_X1    g0155(.A(G150), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n229), .A2(G33), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n355), .B1(new_n356), .B2(new_n275), .C1(new_n317), .C2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n284), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n201), .B1(new_n306), .B2(G20), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT67), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n320), .A2(new_n284), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n359), .B(new_n363), .C1(G50), .C2(new_n319), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT9), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n352), .A2(G200), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n354), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  OR3_X1    g0169(.A1(new_n369), .A2(KEYINPUT71), .A3(KEYINPUT10), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT71), .B1(new_n369), .B2(KEYINPUT10), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT72), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT72), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n375), .A3(KEYINPUT10), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n309), .B1(new_n350), .B2(new_n220), .ZN(new_n379));
  XNOR2_X1  g0179(.A(new_n379), .B(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G238), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n272), .B(new_n381), .C1(new_n207), .C2(G1698), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT70), .B(G107), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n304), .C1(new_n272), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(G200), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G20), .A2(G77), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT15), .B(G87), .Z(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI221_X1 g0190(.A(new_n388), .B1(new_n275), .B2(new_n317), .C1(new_n390), .C2(new_n357), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n391), .A2(new_n284), .B1(new_n219), .B2(new_n320), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n322), .A2(G77), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n387), .B(new_n394), .C1(new_n315), .C2(new_n386), .ZN(new_n395));
  INV_X1    g0195(.A(G169), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n352), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n364), .C1(G179), .C2(new_n352), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT68), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n394), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n386), .A2(new_n396), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n401), .B(new_n402), .C1(G179), .C2(new_n386), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n378), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n207), .A2(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(G226), .B2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n286), .A2(new_n268), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n304), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(new_n309), .C1(new_n218), .C2(new_n350), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT13), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n412), .B(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G190), .ZN(new_n417));
  OAI22_X1  g0217(.A1(new_n275), .A2(new_n201), .B1(new_n357), .B2(new_n219), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n229), .A2(G68), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n284), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT11), .ZN(new_n421));
  OAI22_X1  g0221(.A1(new_n420), .A2(new_n421), .B1(new_n323), .B2(new_n203), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n306), .A3(G13), .ZN(new_n424));
  XOR2_X1   g0224(.A(new_n424), .B(KEYINPUT12), .Z(new_n425));
  NOR3_X1   g0225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n414), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(G169), .ZN(new_n429));
  XOR2_X1   g0229(.A(new_n429), .B(KEYINPUT14), .Z(new_n430));
  INV_X1    g0230(.A(new_n416), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n430), .B1(new_n339), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n426), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n343), .A2(KEYINPUT79), .ZN(new_n435));
  AND4_X1   g0235(.A1(new_n344), .A2(new_n405), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n285), .A2(new_n229), .A3(G68), .A4(new_n286), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT19), .ZN(new_n438));
  NOR2_X1   g0238(.A1(G87), .A2(G97), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n383), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n406), .A2(new_n229), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n406), .A2(KEYINPUT19), .A3(G20), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n284), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n389), .A2(new_n319), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n306), .A2(G33), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n362), .A2(G87), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G200), .ZN(new_n452));
  MUX2_X1   g0252(.A(G238), .B(G244), .S(G1698), .Z(new_n453));
  NAND2_X1  g0253(.A1(new_n294), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n246), .B1(new_n262), .B2(new_n263), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n304), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT82), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n308), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n304), .A2(new_n209), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n459), .B(new_n462), .C1(new_n463), .C2(new_n461), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n461), .B1(new_n311), .B2(G250), .ZN(new_n465));
  INV_X1    g0265(.A(new_n462), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT82), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n452), .B1(new_n458), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT84), .B1(new_n451), .B2(new_n469), .ZN(new_n470));
  AOI211_X1 g0270(.A(new_n446), .B(new_n449), .C1(new_n444), .C2(new_n284), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n464), .A2(new_n467), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n311), .B1(new_n454), .B2(new_n456), .ZN(new_n473));
  OAI21_X1  g0273(.A(G200), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT84), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n471), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n472), .A2(new_n473), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n458), .A2(new_n468), .A3(G179), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n477), .B2(new_n396), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n362), .A2(new_n448), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n389), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n445), .A2(new_n447), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n445), .A2(new_n486), .A3(new_n447), .A4(new_n483), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT85), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n479), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(new_n479), .B2(new_n488), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n310), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT5), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G41), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n461), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n311), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n214), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n308), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n294), .A2(KEYINPUT89), .A3(G257), .A4(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n285), .A2(G257), .A3(G1698), .A4(new_n286), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n294), .A2(G250), .A3(new_n346), .ZN(new_n504));
  XOR2_X1   g0304(.A(KEYINPUT90), .B(G294), .Z(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n264), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n500), .A2(new_n503), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n498), .B(new_n499), .C1(new_n507), .C2(new_n304), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G190), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n304), .ZN(new_n510));
  INV_X1    g0310(.A(new_n498), .ZN(new_n511));
  INV_X1    g0311(.A(new_n499), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n229), .B1(new_n455), .B2(KEYINPUT23), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n229), .A2(KEYINPUT23), .A3(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n208), .A2(G20), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n286), .A3(new_n268), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT22), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n285), .A2(KEYINPUT22), .A3(new_n286), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n384), .A2(KEYINPUT23), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n515), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT24), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n306), .A2(new_n213), .A3(G13), .A4(G20), .ZN(new_n525));
  OR2_X1    g0325(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT25), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n362), .A2(G107), .A3(new_n448), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(KEYINPUT25), .A3(new_n527), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT88), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n530), .A2(new_n535), .A3(new_n531), .A4(new_n532), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n524), .A2(new_n284), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n509), .A2(new_n514), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n513), .A2(new_n396), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n536), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n523), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n523), .A2(new_n541), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n284), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n510), .A2(new_n339), .A3(new_n511), .A4(new_n512), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n539), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT91), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n547), .A3(KEYINPUT91), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n383), .B1(new_n270), .B2(new_n273), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n275), .A2(new_n219), .ZN(new_n554));
  XNOR2_X1  g0354(.A(G97), .B(G107), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n556), .A2(KEYINPUT80), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(G97), .ZN(new_n558));
  OR3_X1    g0358(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n555), .A2(new_n557), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n229), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n553), .A2(new_n554), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n284), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n285), .A2(G244), .A3(new_n346), .A4(new_n286), .ZN(new_n565));
  XOR2_X1   g0365(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n566));
  AOI22_X1  g0366(.A1(new_n565), .A2(new_n566), .B1(G33), .B2(G283), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n346), .A2(KEYINPUT4), .A3(G244), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n568), .B1(new_n209), .B2(new_n346), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n272), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n499), .B1(new_n571), .B2(new_n304), .ZN(new_n572));
  INV_X1    g0372(.A(G257), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n497), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n452), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n311), .B1(new_n567), .B2(new_n570), .ZN(new_n577));
  NOR4_X1   g0377(.A1(new_n577), .A2(new_n315), .A3(new_n499), .A4(new_n574), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n320), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n482), .A2(G97), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n564), .A2(new_n579), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n214), .A2(G1698), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n573), .A2(new_n346), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n285), .A2(new_n286), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n409), .A2(G303), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n311), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n496), .A2(G270), .A3(new_n311), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n588), .A2(new_n499), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n362), .A2(G116), .A3(new_n448), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n306), .A2(new_n246), .A3(G13), .A4(G20), .ZN(new_n592));
  XNOR2_X1  g0392(.A(new_n592), .B(KEYINPUT86), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n283), .A2(new_n228), .B1(G20), .B2(new_n246), .ZN(new_n594));
  AOI21_X1  g0394(.A(G20), .B1(G33), .B2(G283), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G33), .B2(new_n580), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n596), .A3(KEYINPUT20), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT20), .B1(new_n594), .B2(new_n596), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n591), .B(new_n593), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n590), .A2(G179), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n590), .A2(G190), .ZN(new_n601));
  INV_X1    g0401(.A(new_n599), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n452), .C2(new_n590), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT21), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n590), .A2(new_n396), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n599), .ZN(new_n606));
  NOR4_X1   g0406(.A1(new_n590), .A2(new_n602), .A3(KEYINPUT21), .A4(new_n396), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n600), .B(new_n603), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n581), .B(new_n582), .C1(new_n562), .C2(new_n563), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n577), .A2(new_n499), .A3(new_n574), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n339), .ZN(new_n612));
  INV_X1    g0412(.A(new_n611), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n396), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n583), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  AND4_X1   g0416(.A1(new_n436), .A2(new_n492), .A3(new_n552), .A4(new_n616), .ZN(G372));
  INV_X1    g0417(.A(new_n400), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n432), .A2(new_n433), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n428), .B1(new_n619), .B2(new_n403), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n329), .A3(new_n332), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n341), .A2(new_n342), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n623), .B2(new_n378), .ZN(new_n624));
  INV_X1    g0424(.A(new_n436), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n481), .A2(new_n484), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n478), .A2(new_n474), .A3(new_n471), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n630), .B2(new_n547), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n538), .A3(new_n615), .A4(new_n583), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n626), .B(KEYINPUT92), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n615), .A2(new_n628), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT26), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n490), .A2(new_n491), .A3(new_n615), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n632), .B(new_n636), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n624), .B1(new_n625), .B2(new_n639), .ZN(G369));
  NAND3_X1  g0440(.A1(new_n550), .A2(new_n547), .A3(new_n551), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n630), .A2(new_n547), .ZN(new_n642));
  INV_X1    g0442(.A(G13), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G20), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n306), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT27), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(G343), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n641), .A2(new_n642), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n552), .B1(new_n537), .B2(new_n651), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n547), .A2(new_n651), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n651), .A2(new_n602), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n629), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT93), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n608), .B(KEYINPUT94), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n652), .B1(new_n656), .B2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n232), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n383), .A2(new_n246), .A3(new_n439), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n665), .A2(new_n666), .A3(new_n306), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n227), .B2(new_n665), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT28), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n637), .A2(new_n635), .ZN(new_n670));
  INV_X1    g0470(.A(new_n633), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n615), .B2(new_n628), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n632), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n651), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n639), .A2(KEYINPUT29), .A3(new_n650), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n616), .A2(new_n552), .A3(new_n492), .A4(new_n651), .ZN(new_n679));
  INV_X1    g0479(.A(new_n480), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n588), .A2(new_n589), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n508), .A2(new_n680), .A3(new_n611), .A4(new_n681), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT30), .Z(new_n683));
  XOR2_X1   g0483(.A(new_n477), .B(KEYINPUT95), .Z(new_n684));
  NOR3_X1   g0484(.A1(new_n508), .A2(G179), .A3(new_n590), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n684), .A2(new_n613), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n650), .B1(new_n683), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n679), .A2(KEYINPUT31), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(KEYINPUT31), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n678), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n669), .B1(new_n693), .B2(G1), .ZN(G364));
  INV_X1    g0494(.A(new_n665), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n644), .A2(G45), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n229), .A2(new_n339), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(new_n315), .A3(new_n452), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n229), .A2(G179), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(G190), .A3(G200), .ZN(new_n702));
  OAI22_X1  g0502(.A1(new_n700), .A2(new_n219), .B1(new_n702), .B2(new_n208), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(G190), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n452), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n272), .B1(new_n706), .B2(new_n201), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n699), .A2(new_n315), .A3(G200), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n703), .B(new_n707), .C1(G68), .C2(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n315), .A2(G179), .A3(G200), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n229), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n580), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n701), .A2(new_n315), .A3(G200), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT98), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n704), .A2(G200), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n717), .A2(G107), .B1(G58), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n701), .A2(new_n315), .A3(new_n452), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n276), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT32), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n710), .A2(new_n714), .A3(new_n719), .A4(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n712), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n505), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n718), .A2(G322), .B1(new_n705), .B2(G326), .ZN(new_n726));
  INV_X1    g0526(.A(new_n700), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G311), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n717), .A2(G283), .ZN(new_n730));
  XOR2_X1   g0530(.A(KEYINPUT99), .B(G317), .Z(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT33), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n709), .ZN(new_n733));
  INV_X1    g0533(.A(G303), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n409), .B1(new_n702), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n720), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(G329), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n729), .A2(new_n730), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n723), .B1(new_n725), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n228), .B1(G20), .B2(new_n396), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n643), .A2(new_n261), .A3(KEYINPUT97), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT97), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(G13), .B2(G33), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n272), .A2(G355), .A3(new_n232), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G116), .B2(new_n232), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT96), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n294), .A2(new_n664), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n227), .A2(new_n460), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n751), .B(new_n752), .C1(new_n252), .C2(new_n460), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(new_n739), .A2(new_n740), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n746), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n698), .B(new_n755), .C1(new_n661), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n662), .A2(new_n697), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n661), .A2(G330), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(G396));
  OAI21_X1  g0560(.A(new_n395), .B1(new_n394), .B2(new_n651), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n403), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n403), .A2(new_n650), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n639), .B2(new_n650), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n638), .A2(new_n651), .A3(new_n764), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(new_n691), .Z(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n697), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n716), .A2(new_n203), .ZN(new_n771));
  INV_X1    g0571(.A(G132), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n294), .B1(new_n201), .B2(new_n702), .C1(new_n772), .C2(new_n720), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G143), .A2(new_n718), .B1(new_n709), .B2(G150), .ZN(new_n774));
  INV_X1    g0574(.A(G137), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n774), .B1(new_n775), .B2(new_n706), .C1(new_n276), .C2(new_n700), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT34), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n771), .B(new_n773), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n778), .B1(new_n777), .B2(new_n776), .C1(new_n202), .C2(new_n712), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n706), .A2(new_n734), .B1(new_n246), .B2(new_n700), .ZN(new_n780));
  INV_X1    g0580(.A(new_n702), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n713), .B(new_n780), .C1(G107), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n717), .A2(G87), .ZN(new_n783));
  INV_X1    g0583(.A(new_n718), .ZN(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n785), .B1(new_n786), .B2(new_n708), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G311), .B2(new_n736), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n782), .A2(new_n409), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n779), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n744), .A2(new_n740), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n790), .A2(new_n740), .B1(new_n219), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n792), .B(new_n698), .C1(new_n764), .C2(new_n745), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n770), .A2(new_n793), .ZN(G384));
  OAI21_X1  g0594(.A(new_n434), .B1(new_n426), .B2(new_n651), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n433), .B(new_n650), .C1(new_n432), .C2(new_n428), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n690), .A2(new_n764), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT102), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT38), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT101), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n331), .B2(new_n648), .ZN(new_n802));
  INV_X1    g0602(.A(new_n648), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n337), .A2(KEYINPUT101), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n337), .A2(new_n340), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n806), .A2(new_n327), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT37), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n805), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n255), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n292), .A2(new_n811), .A3(new_n298), .A4(new_n284), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n325), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n803), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(KEYINPUT100), .A3(new_n803), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n340), .A2(new_n813), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n816), .A2(new_n327), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(KEYINPUT37), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n809), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n816), .A2(new_n817), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n343), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n799), .B(new_n800), .C1(new_n821), .C2(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n809), .A2(new_n820), .B1(new_n343), .B2(new_n822), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT102), .B1(new_n825), .B2(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT38), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n798), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT40), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n805), .A2(new_n807), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n833));
  INV_X1    g0633(.A(new_n805), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n833), .A2(new_n809), .B1(new_n343), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n827), .B1(new_n835), .B2(KEYINPUT38), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n798), .A2(KEYINPUT40), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n436), .A2(new_n690), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n838), .B(new_n839), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G330), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT104), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n436), .B1(new_n676), .B2(new_n677), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n624), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n842), .B(new_n844), .Z(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT39), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n827), .B(new_n848), .C1(new_n835), .C2(KEYINPUT38), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n847), .A2(new_n846), .A3(new_n849), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n619), .A2(new_n650), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n767), .A2(new_n763), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n795), .A2(new_n796), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n853), .A2(new_n854), .B1(new_n828), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n622), .B2(new_n803), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n845), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n860), .B1(new_n306), .B2(new_n644), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n559), .A2(new_n560), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n246), .B1(new_n862), .B2(KEYINPUT35), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n230), .C1(KEYINPUT35), .C2(new_n862), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT36), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n278), .A2(G77), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n226), .A2(new_n866), .B1(G50), .B2(new_n203), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n867), .A2(G1), .A3(new_n643), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n861), .A2(new_n865), .A3(new_n868), .ZN(G367));
  NOR2_X1   g0669(.A1(new_n630), .A2(new_n650), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n552), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n583), .A2(new_n615), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n610), .A2(new_n650), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n615), .A2(new_n651), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT42), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n615), .B1(new_n874), .B2(new_n547), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n651), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n451), .A2(new_n650), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n628), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n633), .B2(new_n880), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT105), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n877), .A2(new_n879), .B1(KEYINPUT43), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n656), .A2(new_n662), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n874), .A2(new_n875), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n885), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n884), .A2(KEYINPUT43), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n665), .B(new_n892), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n652), .A2(new_n872), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT44), .Z(new_n896));
  NAND2_X1  g0696(.A1(new_n887), .A2(new_n652), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT45), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(new_n886), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n871), .B1(new_n655), .B2(new_n870), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n661), .A2(KEYINPUT107), .A3(G330), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT107), .B1(new_n661), .B2(G330), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n901), .A2(new_n903), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n900), .A2(new_n693), .A3(new_n904), .A4(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n894), .B1(new_n906), .B2(new_n693), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n696), .A2(G1), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n891), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n751), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n747), .B1(new_n232), .B2(new_n390), .C1(new_n910), .C2(new_n243), .ZN(new_n911));
  INV_X1    g0711(.A(new_n715), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n781), .A2(G58), .B1(new_n912), .B2(G77), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n272), .C1(new_n276), .C2(new_n708), .ZN(new_n914));
  AOI22_X1  g0714(.A1(G68), .A2(new_n724), .B1(new_n727), .B2(G50), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n705), .A2(G143), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(new_n356), .C2(new_n784), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n914), .B(new_n917), .C1(G137), .C2(new_n736), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(G97), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT108), .B(G311), .Z(new_n920));
  AOI22_X1  g0720(.A1(new_n705), .A2(new_n920), .B1(new_n709), .B2(new_n505), .ZN(new_n921));
  OAI221_X1 g0721(.A(new_n921), .B1(new_n786), .B2(new_n700), .C1(new_n734), .C2(new_n784), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n702), .A2(new_n246), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT46), .ZN(new_n924));
  INV_X1    g0724(.A(new_n294), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n925), .B1(new_n926), .B2(new_n720), .C1(new_n383), .C2(new_n712), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n922), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n918), .B1(new_n919), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT47), .Z(new_n930));
  AOI21_X1  g0730(.A(new_n697), .B1(new_n930), .B2(new_n740), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n911), .B(new_n931), .C1(new_n884), .C2(new_n756), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n909), .A2(new_n932), .ZN(G387));
  NAND2_X1  g0733(.A1(new_n905), .A2(new_n904), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n692), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n695), .B1(new_n692), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n666), .A2(new_n232), .A3(new_n272), .ZN(new_n938));
  AOI211_X1 g0738(.A(G45), .B(new_n666), .C1(G68), .C2(G77), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT50), .B1(new_n317), .B2(G50), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n317), .A2(KEYINPUT50), .A3(G50), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n944), .A2(new_n945), .B1(new_n460), .B2(new_n240), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n938), .B1(G107), .B2(new_n232), .C1(new_n946), .C2(new_n910), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n747), .B1(new_n947), .B2(KEYINPUT110), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(KEYINPUT110), .B2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n781), .A2(new_n505), .ZN(new_n950));
  AOI22_X1  g0750(.A1(G322), .A2(new_n705), .B1(new_n727), .B2(G303), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n709), .A2(new_n920), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n926), .C2(new_n784), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT48), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n950), .B1(new_n786), .B2(new_n712), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT112), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT49), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n736), .A2(G326), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT49), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n294), .B1(G116), .B2(new_n912), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n959), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT111), .B(G150), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n925), .B1(new_n736), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n201), .B2(new_n784), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n724), .A2(new_n389), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n203), .B2(new_n700), .C1(new_n706), .C2(new_n276), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n318), .C2(new_n709), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n219), .B2(new_n702), .C1(new_n580), .C2(new_n716), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n971), .B2(new_n740), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n698), .C1(new_n655), .C2(new_n756), .ZN(new_n973));
  INV_X1    g0773(.A(new_n908), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n937), .B(new_n973), .C1(new_n974), .C2(new_n934), .ZN(G393));
  XNOR2_X1  g0775(.A(new_n900), .B(new_n935), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n665), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n900), .A2(new_n908), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n718), .A2(G311), .B1(new_n705), .B2(G317), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT52), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n717), .A2(G107), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n781), .A2(G283), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n409), .B1(new_n712), .B2(new_n246), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n700), .A2(new_n785), .B1(new_n708), .B2(new_n734), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(G322), .C2(new_n736), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n718), .A2(G159), .B1(new_n705), .B2(G150), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT51), .Z(new_n988));
  AOI22_X1  g0788(.A1(new_n717), .A2(G87), .B1(G68), .B2(new_n781), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n712), .A2(new_n219), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n318), .B2(new_n727), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n201), .B2(new_n708), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n925), .B1(G143), .B2(new_n736), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n988), .A2(new_n989), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n992), .A2(KEYINPUT113), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n986), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n740), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n249), .A2(new_n751), .B1(G97), .B2(new_n664), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n747), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(new_n698), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT114), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n887), .B2(new_n756), .ZN(new_n1003));
  AND3_X1   g0803(.A1(new_n977), .A2(new_n978), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(G390));
  OAI22_X1  g0805(.A1(new_n784), .A2(new_n246), .B1(new_n706), .B2(new_n786), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G97), .B2(new_n727), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n208), .B2(new_n702), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n990), .B1(new_n384), .B2(new_n709), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n785), .B2(new_n720), .ZN(new_n1010));
  OR4_X1    g0810(.A1(new_n272), .A2(new_n1008), .A3(new_n771), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n715), .A2(new_n201), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n784), .A2(new_n772), .B1(new_n775), .B2(new_n708), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G128), .C2(new_n705), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n781), .A2(new_n964), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT53), .Z(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT54), .B(G143), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT119), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n727), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n409), .B1(new_n724), .B2(G159), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n736), .A2(G125), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n1023), .A2(new_n740), .B1(new_n317), .B2(new_n791), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n698), .B(new_n1024), .C1(new_n853), .C2(new_n745), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT120), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n690), .A2(G330), .A3(new_n764), .A4(new_n797), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n847), .A2(new_n846), .A3(new_n849), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n857), .A2(new_n854), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1030), .A2(new_n850), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n674), .A2(new_n762), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n763), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n797), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n854), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n1036), .A3(new_n836), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1029), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1031), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n851), .A2(new_n852), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1041), .A2(new_n1037), .A3(new_n1028), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n908), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1027), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(G330), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n843), .B(new_n624), .C1(new_n1046), .C2(new_n839), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT115), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n688), .A2(G330), .A3(new_n689), .A4(new_n764), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n856), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1028), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n855), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI211_X1 g0853(.A(KEYINPUT115), .B(new_n855), .C1(new_n1028), .C2(new_n1050), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1051), .A2(new_n1034), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1047), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1039), .A2(new_n1042), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT116), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT116), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1039), .A2(new_n1057), .A3(new_n1042), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n665), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT117), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1057), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1062), .A2(KEYINPUT117), .A3(new_n665), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(KEYINPUT118), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT118), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1065), .A2(new_n1072), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1045), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G378));
  NAND2_X1  g0875(.A1(new_n364), .A2(new_n803), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n378), .A2(new_n398), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1078), .A2(KEYINPUT121), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1077), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1081), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n1079), .A3(new_n1076), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1090), .A2(G330), .A3(new_n831), .A4(new_n837), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1088), .C1(new_n838), .C2(new_n1046), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n859), .B(new_n1093), .Z(new_n1094));
  INV_X1    g0894(.A(new_n1047), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1062), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1096), .A3(KEYINPUT57), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT122), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1091), .A2(new_n1092), .A3(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n859), .B(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1095), .B2(new_n1062), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1097), .B(new_n665), .C1(new_n1101), .C2(KEYINPUT57), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1100), .A2(new_n974), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1090), .A2(new_n744), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n791), .A2(new_n201), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n724), .A2(G68), .B1(new_n781), .B2(G77), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n390), .B2(new_n700), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n706), .A2(new_n246), .B1(new_n580), .B2(new_n708), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n925), .B(new_n310), .C1(new_n786), .C2(new_n720), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n715), .A2(new_n202), .ZN(new_n1110));
  NOR4_X1   g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n213), .B2(new_n784), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT58), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1018), .A2(new_n781), .B1(G132), .B2(new_n709), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n724), .A2(G150), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n718), .A2(G128), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G125), .A2(new_n705), .B1(new_n727), .B2(G137), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT59), .Z(new_n1119));
  AOI21_X1  g0919(.A(G41), .B1(new_n912), .B2(G159), .ZN(new_n1120));
  AOI21_X1  g0920(.A(G33), .B1(new_n736), .B2(G124), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(G41), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1113), .B(new_n1122), .C1(G50), .C2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n697), .B1(new_n1124), .B2(new_n740), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1104), .A2(new_n1105), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1102), .A2(new_n1103), .A3(new_n1126), .ZN(G375));
  NAND3_X1  g0927(.A1(new_n1055), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1067), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n894), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT123), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n974), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n856), .A2(new_n744), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n409), .B1(new_n716), .B2(new_n219), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT124), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n706), .A2(new_n785), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n784), .A2(new_n786), .B1(new_n246), .B2(new_n708), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n967), .B1(new_n580), .B2(new_n702), .C1(new_n734), .C2(new_n720), .ZN(new_n1139));
  NOR4_X1   g0939(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n1135), .B2(new_n1134), .C1(new_n383), .C2(new_n700), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n700), .A2(new_n356), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n712), .A2(new_n201), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n784), .A2(new_n775), .B1(new_n276), .B2(new_n702), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G132), .C2(new_n705), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1018), .A2(new_n709), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1110), .B(new_n925), .C1(G128), .C2(new_n736), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1141), .B1(new_n1142), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1149), .A2(new_n740), .B1(new_n203), .B2(new_n791), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1133), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1132), .B1(new_n698), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1131), .A2(new_n1152), .ZN(G381));
  INV_X1    g0953(.A(new_n1045), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1070), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1156), .A2(G375), .ZN(new_n1157));
  NOR4_X1   g0957(.A1(G390), .A2(G387), .A3(G396), .A4(G393), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(G381), .A2(G384), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(G407));
  INV_X1    g0960(.A(G213), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n1157), .B2(new_n649), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(G407), .ZN(G409));
  XNOR2_X1  g0963(.A(G387), .B(new_n1004), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(G393), .B(G396), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1101), .A2(new_n893), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1094), .A2(new_n908), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n1126), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1155), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1074), .B2(G375), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1129), .A2(KEYINPUT60), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1128), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n665), .C1(KEYINPUT60), .C2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1174), .A2(G384), .A3(new_n1152), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G384), .B1(new_n1174), .B2(new_n1152), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1161), .A2(G343), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1171), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(G2897), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1177), .B(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1171), .B2(new_n1179), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1180), .B1(new_n1183), .B2(KEYINPUT62), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT125), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1171), .A2(KEYINPUT125), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT62), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1166), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT61), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT63), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1180), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(new_n1183), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1188), .A2(new_n1189), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1166), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1191), .A2(new_n1199), .ZN(G405));
  NAND2_X1  g1000(.A1(G375), .A2(new_n1155), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1074), .B2(G375), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(new_n1166), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(new_n1177), .ZN(G402));
endmodule


