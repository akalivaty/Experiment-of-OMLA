//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n212, new_n213, new_n214, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1293, new_n1294, new_n1295, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351;
  INV_X1    g0000(.A(KEYINPUT65), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(KEYINPUT64), .ZN(new_n205));
  OAI21_X1  g0005(.A(new_n205), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n201), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI211_X1 g0009(.A(KEYINPUT65), .B(G50), .C1(new_n204), .C2(new_n206), .ZN(new_n210));
  NOR3_X1   g0010(.A1(new_n209), .A2(new_n210), .A3(G77), .ZN(G353));
  INV_X1    g0011(.A(G97), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G87), .ZN(G355));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT0), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n207), .A2(new_n208), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n217), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n203), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n234));
  AOI22_X1  g0034(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n231), .A2(new_n232), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n219), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI211_X1 g0038(.A(new_n222), .B(new_n226), .C1(new_n238), .C2(KEYINPUT1), .ZN(new_n239));
  AOI21_X1  g0039(.A(new_n239), .B1(KEYINPUT1), .B2(new_n238), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G250), .B(G257), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G264), .B(G270), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G358));
  NAND2_X1  g0049(.A1(new_n208), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n203), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n224), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT8), .B(G58), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n263), .A2(new_n264), .B1(G20), .B2(G77), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT15), .B(G87), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n261), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n260), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n216), .A2(G20), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G77), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n275), .A2(new_n277), .B1(G77), .B2(new_n272), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT70), .B1(new_n271), .B2(new_n278), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n268), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(G1698), .ZN(new_n290));
  OAI221_X1 g0090(.A(new_n289), .B1(new_n213), .B2(new_n287), .C1(new_n290), .C2(new_n228), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  OAI211_X1 g0099(.A(G1), .B(G13), .C1(new_n268), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n296), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n230), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n293), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n283), .B1(G200), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(new_n292), .B2(new_n291), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G190), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n305), .A2(new_n307), .B1(new_n283), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n298), .B1(new_n312), .B2(new_n301), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n287), .A2(G222), .A3(new_n288), .ZN(new_n314));
  XOR2_X1   g0114(.A(KEYINPUT68), .B(G223), .Z(new_n315));
  OAI221_X1 g0115(.A(new_n314), .B1(new_n229), .B2(new_n287), .C1(new_n290), .C2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n313), .B1(new_n316), .B2(new_n292), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G169), .B2(new_n317), .ZN(new_n320));
  INV_X1    g0120(.A(new_n269), .ZN(new_n321));
  INV_X1    g0121(.A(G150), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n217), .A2(new_n268), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n262), .A2(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT69), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(G20), .B1(new_n209), .B2(new_n210), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n261), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n276), .A2(G50), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n275), .A2(new_n329), .B1(G50), .B2(new_n272), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n320), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT9), .ZN(new_n333));
  INV_X1    g0133(.A(new_n330), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n326), .A2(new_n327), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n261), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT9), .B1(new_n328), .B2(new_n330), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G200), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n317), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT71), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT10), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(G190), .B2(new_n317), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n338), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n338), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n311), .B(new_n332), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n287), .A2(G226), .A3(new_n288), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n287), .A2(G232), .A3(G1698), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n292), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n352));
  INV_X1    g0152(.A(new_n301), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(G238), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT13), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G190), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT72), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n351), .A2(new_n357), .A3(new_n354), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n357), .B1(new_n351), .B2(new_n354), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT72), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n365), .A3(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n264), .A2(G50), .ZN(new_n368));
  XOR2_X1   g0168(.A(new_n368), .B(KEYINPUT73), .Z(new_n369));
  OAI22_X1  g0169(.A1(new_n321), .A2(new_n229), .B1(new_n217), .B2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n260), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT11), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g0173(.A(KEYINPUT11), .B(new_n260), .C1(new_n369), .C2(new_n370), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT12), .B1(new_n272), .B2(G68), .ZN(new_n375));
  OR3_X1    g0175(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n203), .B1(new_n216), .B2(G20), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n375), .A2(new_n376), .B1(new_n274), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n364), .B2(new_n339), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n367), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G169), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n356), .B2(new_n358), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(new_n359), .B2(new_n318), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(G169), .C1(new_n362), .C2(new_n363), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(KEYINPUT74), .A3(new_n385), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n382), .B1(new_n391), .B2(new_n379), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n262), .B1(new_n216), .B2(G20), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n274), .B1(new_n273), .B2(new_n262), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT75), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G33), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n398), .A3(new_n284), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n285), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n203), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n204), .A2(new_n206), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n323), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n395), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n260), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n408), .B2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n284), .B1(new_n396), .B2(new_n398), .ZN(new_n418));
  INV_X1    g0218(.A(new_n285), .ZN(new_n419));
  NOR3_X1   g0219(.A1(new_n418), .A2(G20), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n203), .B1(new_n420), .B2(new_n404), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT75), .B(G33), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n217), .B(new_n285), .C1(new_n422), .C2(new_n284), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT7), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n417), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n394), .B1(new_n415), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n394), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n399), .A2(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n416), .B1(new_n430), .B2(new_n203), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n261), .B1(new_n431), .B2(new_n395), .ZN(new_n432));
  AOI211_X1 g0232(.A(new_n395), .B(new_n411), .C1(new_n408), .C2(G20), .ZN(new_n433));
  OAI21_X1  g0233(.A(G68), .B1(new_n423), .B2(KEYINPUT7), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n396), .A2(new_n398), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n419), .B1(new_n435), .B2(KEYINPUT3), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n404), .B1(new_n436), .B2(new_n217), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n433), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n429), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  INV_X1    g0240(.A(G232), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n298), .B1(new_n441), .B2(new_n301), .ZN(new_n442));
  NOR2_X1   g0242(.A1(G223), .A2(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n312), .B2(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n418), .B2(new_n419), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G87), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n300), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G169), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n352), .B1(G232), .B2(new_n353), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n285), .B1(new_n422), .B2(new_n284), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n444), .B1(G33), .B2(G87), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(G179), .C1(new_n300), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n428), .A2(new_n440), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT18), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n428), .A2(new_n453), .A3(new_n456), .A4(new_n440), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n442), .B2(new_n447), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n449), .B(G190), .C1(new_n300), .C2(new_n451), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n460), .A2(KEYINPUT17), .A3(new_n439), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT17), .B1(new_n460), .B2(new_n439), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n457), .A3(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n346), .A2(new_n392), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n217), .B(G87), .C1(new_n418), .C2(new_n419), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(KEYINPUT80), .A3(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(new_n287), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n474));
  INV_X1    g0274(.A(G87), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n473), .A2(new_n474), .A3(G20), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n435), .A2(new_n217), .A3(G116), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT23), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(G20), .B2(new_n213), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n217), .A2(KEYINPUT23), .A3(G107), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n479), .A2(KEYINPUT83), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT83), .B1(new_n479), .B2(new_n483), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n467), .B1(new_n478), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n476), .B1(new_n469), .B2(new_n470), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n472), .ZN(new_n489));
  INV_X1    g0289(.A(new_n486), .ZN(new_n490));
  INV_X1    g0290(.A(new_n467), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n261), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT25), .B1(new_n273), .B2(new_n213), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n216), .A2(G33), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n272), .A2(new_n497), .A3(new_n224), .A4(new_n259), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n495), .A2(new_n496), .B1(G107), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(G250), .A2(G1698), .ZN(new_n502));
  INV_X1    g0302(.A(G257), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G1698), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n450), .A2(new_n504), .B1(G294), .B2(new_n435), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT84), .B1(new_n505), .B2(new_n300), .ZN(new_n506));
  INV_X1    g0306(.A(new_n504), .ZN(new_n507));
  INV_X1    g0307(.A(G294), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n436), .A2(new_n507), .B1(new_n508), .B2(new_n422), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT84), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n510), .A3(new_n292), .ZN(new_n511));
  OR2_X1    g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NAND2_X1  g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n216), .A2(G45), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AND4_X1   g0316(.A1(G274), .A2(new_n514), .A3(new_n300), .A4(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n515), .B1(new_n512), .B2(new_n513), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n292), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(G264), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n506), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT85), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n506), .A2(new_n511), .A3(new_n523), .A4(new_n520), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n383), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n519), .A2(G264), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n295), .A2(new_n518), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n505), .C2(new_n300), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(new_n318), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n493), .A2(new_n501), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n522), .A2(new_n360), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n339), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n491), .B1(new_n489), .B2(new_n490), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n467), .B(new_n486), .C1(new_n488), .C2(new_n472), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n260), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n536), .A3(new_n500), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n519), .A2(G257), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n527), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n230), .A2(G1698), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n287), .A2(G250), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G283), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT77), .B(new_n540), .C1(new_n418), .C2(new_n419), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT77), .B1(new_n450), .B2(new_n540), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n544), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n539), .B1(new_n549), .B2(new_n292), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n318), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT77), .ZN(new_n552));
  INV_X1    g0352(.A(new_n540), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n436), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n554), .A2(new_n546), .A3(new_n545), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n300), .B1(new_n555), .B2(new_n544), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n383), .B1(new_n556), .B2(new_n539), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n273), .A2(new_n212), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n498), .B2(new_n212), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n264), .A2(G77), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT6), .B1(new_n214), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n560), .B1(new_n564), .B2(new_n217), .C1(new_n430), .C2(new_n213), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n559), .B1(new_n565), .B2(new_n260), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n551), .A2(new_n557), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n550), .A2(G190), .ZN(new_n569));
  OAI21_X1  g0369(.A(G200), .B1(new_n556), .B2(new_n539), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n566), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G238), .A2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n230), .B2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n418), .B2(new_n419), .ZN(new_n575));
  INV_X1    g0375(.A(G116), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n422), .A2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n300), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n300), .A2(G274), .A3(new_n516), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n300), .A2(G250), .A3(new_n515), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n383), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT78), .ZN(new_n584));
  INV_X1    g0384(.A(new_n582), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n577), .B1(new_n450), .B2(new_n574), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n318), .C1(new_n586), .C2(new_n300), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n583), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n584), .B1(new_n583), .B2(new_n587), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n450), .A2(new_n217), .A3(G68), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT19), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n269), .A2(new_n591), .A3(G97), .ZN(new_n592));
  NOR2_X1   g0392(.A1(G97), .A2(G107), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n475), .B1(new_n349), .B2(new_n217), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n592), .B1(new_n594), .B2(new_n591), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n261), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n267), .A2(new_n272), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n498), .A2(new_n266), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n588), .A2(new_n589), .A3(new_n599), .ZN(new_n600));
  MUX2_X1   g0400(.A(G257), .B(G264), .S(G1698), .Z(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n418), .B2(new_n419), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n473), .A2(G303), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n300), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n514), .A2(new_n516), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(G270), .A3(new_n300), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n527), .ZN(new_n607));
  OAI21_X1  g0407(.A(G200), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n272), .A2(new_n576), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n499), .B2(new_n576), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n543), .B(new_n217), .C1(G33), .C2(new_n212), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  AOI22_X1  g0412(.A1(KEYINPUT79), .A2(new_n612), .B1(new_n576), .B2(G20), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT79), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT20), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n611), .A2(new_n613), .A3(new_n260), .A4(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n613), .A3(new_n260), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n614), .A3(KEYINPUT20), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n610), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n450), .A2(new_n601), .B1(G303), .B2(new_n473), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n527), .B(new_n606), .C1(new_n621), .C2(new_n300), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n608), .B(new_n620), .C1(new_n622), .C2(new_n360), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  OAI21_X1  g0424(.A(G169), .B1(new_n604), .B2(new_n607), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n620), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n604), .A2(new_n607), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(G179), .A3(new_n619), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n622), .A2(KEYINPUT21), .A3(G169), .A4(new_n619), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n623), .A2(new_n626), .A3(new_n628), .A4(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n498), .A2(new_n475), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n596), .A2(new_n597), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n579), .A2(new_n582), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G190), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n633), .A2(new_n339), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n600), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n530), .A2(new_n537), .A3(new_n572), .A4(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n466), .A2(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n332), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n391), .A2(new_n379), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n380), .B1(new_n366), .B2(new_n361), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n310), .A2(new_n283), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n463), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n426), .A2(new_n453), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n344), .A2(new_n345), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n641), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT86), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT86), .B1(new_n580), .B2(new_n581), .ZN(new_n655));
  OAI22_X1  g0455(.A1(new_n654), .A2(new_n655), .B1(new_n586), .B2(new_n300), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G200), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n632), .A2(new_n657), .A3(new_n634), .ZN(new_n658));
  INV_X1    g0458(.A(new_n597), .ZN(new_n659));
  INV_X1    g0459(.A(new_n598), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n590), .A2(new_n595), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n659), .B(new_n660), .C1(new_n661), .C2(new_n261), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n383), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(new_n587), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(new_n568), .A3(new_n571), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n537), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n536), .A2(new_n500), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n522), .A2(new_n524), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G169), .ZN(new_n671));
  INV_X1    g0471(.A(new_n529), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n668), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n653), .B1(new_n667), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n530), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n677), .A2(KEYINPUT87), .A3(new_n537), .A4(new_n666), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n664), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n658), .A2(new_n664), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT88), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n568), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n682), .B2(new_n568), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT26), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n568), .A2(new_n600), .A3(new_n637), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n680), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n679), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n652), .B1(new_n691), .B2(new_n466), .ZN(G369));
  AND2_X1   g0492(.A1(new_n530), .A2(new_n537), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n216), .A2(new_n217), .A3(G13), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT89), .Z(new_n698));
  INV_X1    g0498(.A(KEYINPUT90), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(G343), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(G343), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n669), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n693), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n703), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(new_n530), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n620), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n668), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n630), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n676), .A2(new_n703), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n536), .A2(new_n500), .B1(new_n671), .B2(new_n672), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n693), .A2(new_n714), .B1(new_n715), .B2(new_n706), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n713), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n220), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n214), .A2(G87), .A3(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n223), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n720), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT28), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT29), .B(new_n703), .C1(new_n679), .C2(new_n689), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n537), .B(new_n666), .C1(new_n715), .C2(new_n668), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n684), .A2(KEYINPUT26), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n680), .B1(new_n687), .B2(new_n685), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n727), .B1(new_n731), .B2(new_n706), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n509), .A2(new_n292), .B1(G264), .B2(new_n519), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n633), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n622), .A2(new_n318), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n550), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  AND4_X1   g0537(.A1(new_n318), .A2(new_n622), .A3(new_n656), .A4(new_n528), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n549), .A2(new_n292), .ZN(new_n739));
  INV_X1    g0539(.A(new_n539), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n736), .A2(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n734), .A2(new_n550), .A3(KEYINPUT30), .A4(new_n735), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n706), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT31), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n639), .B2(new_n703), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT91), .B1(new_n744), .B2(KEYINPUT31), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n633), .A2(new_n627), .A3(new_n733), .A4(G179), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n737), .B1(new_n741), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n738), .A2(new_n741), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(new_n750), .A3(new_n743), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n703), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT91), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n747), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(G330), .B1(new_n746), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n726), .A2(new_n732), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n725), .B1(new_n759), .B2(G1), .ZN(G364));
  INV_X1    g0560(.A(G13), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n216), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n719), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n712), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n766), .B1(G330), .B2(new_n710), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n224), .B1(G20), .B2(new_n383), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n360), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n217), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n212), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n217), .A2(new_n318), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n360), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n217), .A2(G179), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n360), .A3(G200), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n776), .A2(new_n208), .B1(new_n778), .B2(new_n213), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n774), .A2(G190), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n772), .B(new_n779), .C1(G68), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G159), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT32), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n777), .A2(G190), .A3(G200), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n785), .A2(KEYINPUT32), .B1(new_n788), .B2(G87), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n773), .A2(new_n782), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n287), .B1(new_n790), .B2(new_n229), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n773), .A2(G190), .A3(new_n339), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n791), .B1(G58), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n781), .A2(new_n786), .A3(new_n789), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n473), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(G329), .C2(new_n784), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n775), .A2(G326), .ZN(new_n801));
  XNOR2_X1  g0601(.A(KEYINPUT33), .B(G317), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n780), .A2(new_n802), .B1(new_n788), .B2(G303), .ZN(new_n803));
  INV_X1    g0603(.A(new_n771), .ZN(new_n804));
  INV_X1    g0604(.A(new_n778), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n804), .A2(G294), .B1(new_n805), .B2(G283), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n800), .A2(new_n801), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n769), .B1(new_n795), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G13), .A2(G33), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n768), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  MUX2_X1   g0613(.A(new_n723), .B(new_n254), .S(G45), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n436), .A2(new_n220), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n718), .A2(new_n473), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n818), .A2(G355), .B1(new_n576), .B2(new_n718), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n813), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n765), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n808), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n811), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n710), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n767), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  NAND2_X1  g0626(.A1(new_n703), .A2(new_n283), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT94), .B1(new_n644), .B2(new_n706), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT94), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n310), .A2(new_n829), .A3(new_n283), .A4(new_n703), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n311), .A2(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n691), .B2(new_n703), .ZN(new_n832));
  INV_X1    g0632(.A(new_n831), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n690), .A2(new_n706), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n757), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n765), .B1(new_n835), .B2(new_n757), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n831), .A2(new_n809), .ZN(new_n839));
  INV_X1    g0639(.A(new_n790), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n793), .A2(G143), .B1(new_n840), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  INV_X1    g0642(.A(new_n780), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n841), .B1(new_n776), .B2(new_n842), .C1(new_n322), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G132), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n450), .B1(new_n847), .B2(new_n783), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n778), .A2(new_n203), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G58), .B2(new_n804), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n208), .B2(new_n787), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n846), .A2(new_n848), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n845), .B2(new_n844), .ZN(new_n853));
  INV_X1    g0653(.A(G283), .ZN(new_n854));
  INV_X1    g0654(.A(G303), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n843), .A2(new_n854), .B1(new_n776), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G107), .B2(new_n788), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n792), .A2(new_n508), .B1(new_n783), .B2(new_n798), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n287), .B(new_n858), .C1(G116), .C2(new_n840), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n772), .B1(G87), .B2(new_n805), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n769), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n768), .A2(new_n809), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n821), .B(new_n862), .C1(new_n229), .C2(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT93), .Z(new_n865));
  AOI22_X1  g0665(.A1(new_n837), .A2(new_n838), .B1(new_n839), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n762), .A2(new_n216), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n373), .A2(new_n374), .A3(new_n378), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n703), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n382), .B(new_n870), .C1(new_n391), .C2(new_n379), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n390), .A2(new_n389), .ZN(new_n872));
  OAI21_X1  g0672(.A(G169), .B1(new_n362), .B2(new_n363), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n873), .A2(KEYINPUT14), .B1(new_n364), .B2(G179), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n869), .B(new_n703), .C1(new_n875), .C2(new_n643), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n831), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT40), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n752), .A2(KEYINPUT99), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT99), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n751), .A2(new_n880), .A3(new_n703), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n879), .A2(new_n754), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n877), .B(new_n878), .C1(new_n746), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n460), .A2(new_n439), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n432), .A2(new_n438), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT76), .B1(new_n887), .B2(new_n394), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n427), .B(new_n429), .C1(new_n432), .C2(new_n438), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n890), .B2(new_n453), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT97), .B1(new_n890), .B2(new_n698), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT97), .ZN(new_n893));
  INV_X1    g0693(.A(new_n698), .ZN(new_n894));
  NOR4_X1   g0694(.A1(new_n888), .A2(new_n889), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n891), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n413), .B1(new_n421), .B2(new_n424), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT95), .B(new_n260), .C1(new_n897), .C2(KEYINPUT16), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT95), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n397), .A2(G33), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT3), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n902), .A2(new_n404), .A3(new_n217), .A4(new_n285), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n424), .A2(G68), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n904), .B2(new_n416), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n899), .B1(new_n905), .B2(new_n261), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n898), .A2(new_n906), .A3(new_n438), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n907), .A2(new_n394), .B1(new_n448), .B2(new_n452), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n894), .B1(new_n907), .B2(new_n394), .ZN(new_n909));
  INV_X1    g0709(.A(new_n884), .ZN(new_n910));
  NOR3_X1   g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n896), .B1(new_n911), .B2(new_n885), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n464), .A2(KEYINPUT96), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT96), .B1(new_n464), .B2(new_n909), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n912), .B(KEYINPUT38), .C1(new_n913), .C2(new_n914), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n883), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n879), .A2(new_n754), .A3(new_n881), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(new_n745), .C1(new_n639), .C2(new_n703), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n877), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT98), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n647), .A2(new_n884), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n428), .A2(new_n440), .A3(new_n698), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n893), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n428), .A2(KEYINPUT97), .A3(new_n440), .A4(new_n698), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n924), .B1(new_n929), .B2(new_n885), .ZN(new_n930));
  INV_X1    g0730(.A(new_n925), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n892), .B2(new_n895), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(KEYINPUT98), .A3(KEYINPUT37), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n933), .A3(new_n896), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n649), .A2(new_n463), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n927), .A3(new_n928), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n916), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n923), .B1(new_n938), .B2(new_n918), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n920), .B1(new_n939), .B2(new_n878), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n922), .A2(new_n465), .ZN(new_n941));
  OAI21_X1  g0741(.A(G330), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n942), .A2(KEYINPUT100), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(KEYINPUT100), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT39), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n934), .B2(new_n936), .ZN(new_n948));
  INV_X1    g0748(.A(new_n918), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n642), .A2(new_n706), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n918), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n917), .A2(new_n918), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n871), .A2(new_n876), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n703), .B(new_n831), .C1(new_n679), .C2(new_n689), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n644), .A2(new_n703), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n648), .A2(new_n894), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n465), .B1(new_n726), .B2(new_n732), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n652), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n961), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n868), .B1(new_n946), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n964), .B2(new_n946), .ZN(new_n966));
  INV_X1    g0766(.A(new_n564), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT35), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n968), .A2(G116), .A3(new_n225), .A4(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT36), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n407), .A2(G77), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n250), .B1(new_n723), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(G1), .A3(new_n761), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n966), .A2(new_n971), .A3(new_n974), .ZN(G367));
  OR2_X1    g0775(.A1(new_n706), .A2(new_n632), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n664), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n978), .A2(KEYINPUT101), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n665), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n978), .A2(KEYINPUT101), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n811), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n816), .A2(new_n248), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n812), .C1(new_n220), .C2(new_n266), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n765), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n986), .B(KEYINPUT106), .Z(new_n987));
  OAI22_X1  g0787(.A1(new_n843), .A2(new_n410), .B1(new_n787), .B2(new_n202), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G68), .B2(new_n804), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n792), .A2(new_n322), .B1(new_n783), .B2(new_n842), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n473), .B(new_n990), .C1(G50), .C2(new_n840), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n775), .A2(G143), .B1(new_n805), .B2(G77), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n776), .A2(new_n798), .B1(new_n213), .B2(new_n771), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n450), .B(new_n994), .C1(G97), .C2(new_n805), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n792), .A2(new_n855), .B1(new_n783), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G283), .B2(new_n840), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n787), .A2(new_n576), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n843), .A2(new_n508), .B1(KEYINPUT46), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT46), .B2(new_n1000), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n995), .B(new_n998), .C1(new_n999), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n993), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT47), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n768), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n983), .B(new_n987), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n572), .B1(new_n566), .B2(new_n706), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n568), .B2(new_n706), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n716), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT44), .Z(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n716), .A2(new_n1013), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT103), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n693), .A2(new_n714), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(new_n707), .C2(new_n714), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n711), .A2(KEYINPUT105), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n759), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1023), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n759), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n719), .B(KEYINPUT41), .Z(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n764), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1013), .A2(new_n693), .A3(new_n714), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n568), .B1(new_n1012), .B2(new_n530), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(KEYINPUT42), .B1(new_n706), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(KEYINPUT42), .B2(new_n1036), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT43), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n982), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n982), .A2(new_n1040), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n713), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1044), .A2(new_n1013), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1043), .B1(KEYINPUT102), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1045), .B(KEYINPUT102), .Z(new_n1047));
  OAI21_X1  g0847(.A(new_n1046), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1011), .B1(new_n1035), .B2(new_n1048), .ZN(G387));
  AOI21_X1  g0849(.A(new_n720), .B1(new_n1028), .B2(new_n759), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n759), .B2(new_n1028), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n707), .A2(new_n823), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n721), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n818), .A2(new_n1053), .B1(new_n213), .B2(new_n718), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n245), .A2(G45), .ZN(new_n1055));
  AOI21_X1  g0855(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n263), .A2(KEYINPUT50), .A3(new_n208), .ZN(new_n1057));
  AOI21_X1  g0857(.A(KEYINPUT50), .B1(new_n263), .B2(new_n208), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n721), .B(new_n1056), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n816), .A2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1054), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT108), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n812), .A3(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n793), .A2(G317), .B1(new_n840), .B2(G303), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n776), .B2(new_n796), .C1(new_n798), .C2(new_n843), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n804), .A2(G283), .B1(new_n788), .B2(G294), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(KEYINPUT49), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n778), .A2(new_n576), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n450), .B(new_n1076), .C1(G326), .C2(new_n784), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n776), .A2(new_n410), .B1(new_n778), .B2(new_n212), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n843), .A2(new_n262), .B1(new_n266), .B2(new_n771), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n787), .A2(new_n229), .B1(new_n783), .B2(new_n322), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT109), .Z(new_n1083));
  AOI22_X1  g0883(.A1(new_n793), .A2(G50), .B1(new_n840), .B2(G68), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1081), .A2(new_n1083), .A3(new_n450), .A4(new_n1084), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1078), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n765), .B(new_n1065), .C1(new_n1086), .C2(new_n769), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT110), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1028), .A2(new_n764), .B1(new_n1052), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1051), .A2(new_n1089), .ZN(G393));
  NAND2_X1  g0890(.A1(new_n1021), .A2(new_n1044), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1021), .A2(new_n1044), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1029), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n719), .A3(new_n1031), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n1092), .A2(new_n763), .A3(new_n1093), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G317), .A2(new_n775), .B1(new_n793), .B2(G311), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n473), .B1(new_n783), .B2(new_n796), .C1(new_n508), .C2(new_n790), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n843), .A2(new_n855), .B1(new_n778), .B2(new_n213), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n771), .A2(new_n576), .B1(new_n787), .B2(new_n854), .ZN(new_n1101));
  OR4_X1    g0901(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n776), .A2(new_n322), .B1(new_n410), .B2(new_n792), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT51), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n263), .A2(new_n840), .B1(new_n784), .B2(G143), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n771), .A2(new_n229), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n203), .A2(new_n787), .B1(new_n778), .B2(new_n475), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G50), .C2(new_n780), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n450), .A3(new_n1105), .A4(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n769), .B1(new_n1102), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n816), .A2(new_n257), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n813), .B1(G97), .B2(new_n718), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n821), .B(new_n1110), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1013), .B2(new_n823), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1095), .A2(new_n1096), .A3(new_n1114), .ZN(G390));
  INV_X1    g0915(.A(G330), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n831), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n922), .A2(new_n956), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1120), .A2(new_n951), .B1(new_n950), .B2(new_n953), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n948), .A2(new_n949), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n956), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n731), .A2(new_n706), .A3(new_n833), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n958), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1122), .A2(new_n1126), .A3(new_n952), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1122), .A2(new_n952), .A3(new_n1126), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1117), .B1(new_n746), .B2(new_n756), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(new_n1123), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n950), .A2(new_n953), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n834), .A2(new_n1125), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n952), .B1(new_n1134), .B2(new_n956), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1129), .B(new_n1132), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n956), .B1(new_n922), .B2(new_n1117), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1131), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1130), .A2(new_n1123), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT112), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT112), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1130), .A2(new_n1123), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1142), .A2(new_n1118), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1140), .B1(new_n1145), .B2(new_n1134), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n922), .A2(G330), .A3(new_n465), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT111), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n962), .A3(new_n652), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n720), .B1(new_n1137), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1128), .A2(new_n1154), .A3(new_n1136), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT113), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1137), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1133), .A2(new_n810), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n863), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n765), .B1(new_n263), .B2(new_n1161), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n792), .A2(new_n576), .B1(new_n783), .B2(new_n508), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n287), .B(new_n1163), .C1(G97), .C2(new_n840), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n780), .A2(G107), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1106), .B1(G283), .B2(new_n775), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n849), .B1(G87), .B2(new_n788), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(G125), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n287), .B1(new_n783), .B2(new_n1169), .C1(new_n208), .C2(new_n778), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT114), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n775), .A2(G128), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT54), .B(G143), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1172), .B1(new_n847), .B2(new_n792), .C1(new_n790), .C2(new_n1173), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n843), .A2(new_n842), .B1(new_n410), .B2(new_n771), .ZN(new_n1175));
  OR3_X1    g0975(.A1(new_n1171), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n787), .A2(new_n322), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT115), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT53), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1168), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1162), .B1(new_n1180), .B2(new_n768), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1159), .A2(new_n764), .B1(new_n1160), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1158), .A2(new_n1182), .ZN(G378));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n961), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n651), .A2(new_n332), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n331), .A2(new_n894), .ZN(new_n1187));
  AND2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OR3_X1    g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1191), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n940), .B2(G330), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n922), .A2(new_n877), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n948), .B2(new_n949), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n919), .B1(new_n1198), .B2(KEYINPUT40), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(new_n1116), .A3(new_n1194), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1185), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT118), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT117), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n940), .A2(G330), .A3(new_n1195), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1194), .B1(new_n1199), .B2(new_n1116), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n961), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT118), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n1208), .A3(new_n1185), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1202), .A2(new_n1203), .A3(new_n1206), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n1203), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1208), .B1(new_n1207), .B2(new_n1185), .ZN(new_n1212));
  AOI211_X1 g1012(.A(KEYINPUT118), .B(new_n961), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT120), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1155), .A2(new_n1216), .A3(new_n1151), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1155), .B2(new_n1151), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1184), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(KEYINPUT121), .B(new_n1184), .C1(new_n1215), .C2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1224));
  OAI211_X1 g1024(.A(KEYINPUT57), .B(new_n1224), .C1(new_n1217), .C2(new_n1218), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n719), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1222), .A2(new_n1223), .A3(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1210), .A2(new_n1214), .A3(new_n764), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1195), .A2(new_n809), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n765), .B1(G50), .B2(new_n1161), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n790), .A2(new_n266), .B1(new_n783), .B2(new_n854), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n792), .A2(new_n213), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1233), .A2(KEYINPUT116), .B1(new_n229), .B2(new_n787), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1234), .C1(G68), .C2(new_n804), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n778), .A2(new_n202), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G97), .B2(new_n780), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1233), .A2(KEYINPUT116), .B1(new_n775), .B2(G116), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n450), .A2(G41), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1243));
  AOI211_X1 g1043(.A(G50), .B(new_n1239), .C1(new_n268), .C2(new_n299), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n843), .A2(new_n847), .B1(new_n776), .B2(new_n1169), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n793), .A2(G128), .B1(new_n840), .B2(G137), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n787), .B2(new_n1173), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1246), .B(new_n1248), .C1(G150), .C2(new_n804), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n805), .A2(G159), .ZN(new_n1252));
  AOI211_X1 g1052(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1250), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1242), .B(new_n1245), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1231), .B1(new_n1256), .B2(new_n768), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1230), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1229), .A2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT119), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT119), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1229), .A2(new_n1261), .A3(new_n1258), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1228), .A2(new_n1263), .ZN(G375));
  NAND2_X1  g1064(.A1(new_n1123), .A2(new_n809), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n765), .B1(G68), .B2(new_n1161), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G50), .A2(new_n804), .B1(new_n775), .B2(G132), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n410), .B2(new_n787), .C1(new_n843), .C2(new_n1173), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n793), .A2(G137), .B1(new_n840), .B2(G150), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1236), .A2(new_n436), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n784), .A2(G128), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n790), .A2(new_n213), .B1(new_n783), .B2(new_n855), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G283), .B2(new_n793), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n267), .A2(new_n804), .B1(new_n780), .B2(G116), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n775), .A2(G294), .B1(new_n788), .B2(G97), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n287), .B1(new_n805), .B2(G77), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(KEYINPUT122), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n1268), .A2(new_n1272), .B1(new_n1277), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1266), .B1(new_n1280), .B2(new_n768), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1147), .A2(new_n764), .B1(new_n1265), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1152), .A2(new_n1034), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1283), .B2(new_n1284), .ZN(G381));
  AOI21_X1  g1085(.A(new_n1226), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1286));
  AOI22_X1  g1086(.A1(new_n1286), .A2(new_n1223), .B1(new_n1262), .B2(new_n1260), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1156), .A2(new_n1182), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n866), .A2(new_n825), .A3(new_n1051), .A4(new_n1089), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1291), .ZN(G407));
  NAND3_X1  g1092(.A1(new_n700), .A2(new_n701), .A3(G213), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1287), .A2(new_n1289), .A3(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G407), .A2(new_n1295), .A3(G213), .ZN(G409));
  OAI211_X1 g1096(.A(G390), .B(new_n1011), .C1(new_n1035), .C2(new_n1048), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT125), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(G396), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(G387), .A2(new_n1095), .A3(new_n1096), .A4(new_n1114), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1297), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1298), .A2(new_n1301), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1304));
  AND3_X1   g1104(.A1(new_n1303), .A2(KEYINPUT127), .A3(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1284), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n719), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1308), .A2(new_n1284), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1282), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n866), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G384), .B(new_n1282), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1313), .B(new_n1314), .C1(KEYINPUT124), .C2(new_n1293), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1294), .A2(G2897), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n1315), .B(new_n1316), .ZN(new_n1317));
  OR3_X1    g1117(.A1(new_n1215), .A2(new_n1219), .A3(new_n1033), .ZN(new_n1318));
  OR2_X1    g1118(.A1(new_n1224), .A2(KEYINPUT123), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n763), .B1(new_n1224), .B2(KEYINPUT123), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1319), .A2(new_n1320), .B1(new_n1230), .B2(new_n1257), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1288), .B1(new_n1318), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1287), .B2(G378), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1317), .B1(new_n1323), .B2(new_n1294), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1228), .A2(G378), .A3(new_n1263), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT62), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1327), .A2(new_n1328), .A3(new_n1293), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT61), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1324), .A2(new_n1331), .A3(new_n1332), .ZN(new_n1333));
  XOR2_X1   g1133(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1334));
  AOI21_X1  g1134(.A(new_n1294), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1334), .B1(new_n1335), .B2(new_n1330), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1307), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1327), .A2(new_n1293), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1338), .B1(new_n1339), .B2(new_n1329), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1339), .B2(new_n1317), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1335), .A2(KEYINPUT63), .A3(new_n1330), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1340), .A2(new_n1341), .A3(new_n1342), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1337), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1289), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1325), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1330), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1329), .A3(new_n1325), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1342), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1350), .B(new_n1351), .ZN(G402));
endmodule


