

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782;

  AND2_X1 U372 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U373 ( .A(n400), .B(n411), .ZN(n692) );
  XNOR2_X1 U374 ( .A(n509), .B(n396), .ZN(n523) );
  XNOR2_X1 U375 ( .A(n381), .B(n492), .ZN(n387) );
  INV_X1 U376 ( .A(KEYINPUT64), .ZN(n465) );
  BUF_X1 U377 ( .A(n735), .Z(n746) );
  OR2_X2 U378 ( .A1(n747), .A2(G902), .ZN(n537) );
  XNOR2_X2 U379 ( .A(G113), .B(KEYINPUT88), .ZN(n458) );
  XNOR2_X2 U380 ( .A(n350), .B(n351), .ZN(n412) );
  NOR2_X2 U381 ( .A1(n586), .A2(n518), .ZN(n350) );
  XNOR2_X2 U382 ( .A(n554), .B(n526), .ZN(n698) );
  XNOR2_X2 U383 ( .A(n525), .B(G469), .ZN(n554) );
  XNOR2_X1 U384 ( .A(n588), .B(n587), .ZN(n685) );
  NOR2_X1 U385 ( .A1(n606), .A2(n584), .ZN(n572) );
  INV_X2 U386 ( .A(G143), .ZN(n493) );
  AND2_X1 U387 ( .A1(n756), .A2(n649), .ZN(n650) );
  AND2_X1 U388 ( .A1(n373), .A2(n372), .ZN(n371) );
  AND2_X1 U389 ( .A1(n407), .A2(n406), .ZN(n401) );
  AND2_X1 U390 ( .A1(n390), .A2(n604), .ZN(n360) );
  NOR2_X1 U391 ( .A1(n634), .A2(n629), .ZN(n626) );
  OR2_X1 U392 ( .A1(n609), .A2(n608), .ZN(n639) );
  XNOR2_X1 U393 ( .A(n572), .B(n571), .ZN(n727) );
  XNOR2_X1 U394 ( .A(n585), .B(n391), .ZN(n606) );
  XNOR2_X1 U395 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U396 ( .A(n500), .B(n353), .ZN(n559) );
  XNOR2_X1 U397 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U398 ( .A(n395), .B(G131), .ZN(n522) );
  XNOR2_X1 U399 ( .A(KEYINPUT16), .B(G122), .ZN(n459) );
  INV_X1 U400 ( .A(n692), .ZN(n756) );
  XOR2_X1 U401 ( .A(KEYINPUT71), .B(KEYINPUT22), .Z(n351) );
  XNOR2_X2 U402 ( .A(n546), .B(G472), .ZN(n615) );
  NOR2_X1 U403 ( .A1(n727), .A2(n586), .ZN(n573) );
  NOR2_X2 U404 ( .A1(n556), .A2(n555), .ZN(n683) );
  XNOR2_X2 U405 ( .A(n493), .B(G128), .ZN(n509) );
  XNOR2_X1 U406 ( .A(n392), .B(n523), .ZN(n769) );
  XNOR2_X1 U407 ( .A(n522), .B(n393), .ZN(n392) );
  XNOR2_X1 U408 ( .A(n394), .B(KEYINPUT4), .ZN(n393) );
  INV_X1 U409 ( .A(G137), .ZN(n394) );
  NOR2_X1 U410 ( .A1(n739), .A2(G902), .ZN(n525) );
  AND2_X1 U411 ( .A1(n638), .A2(n680), .ZN(n421) );
  NAND2_X1 U412 ( .A1(n360), .A2(n389), .ZN(n388) );
  INV_X1 U413 ( .A(n717), .ZN(n389) );
  XNOR2_X1 U414 ( .A(n616), .B(KEYINPUT110), .ZN(n617) );
  OR2_X1 U415 ( .A1(n483), .A2(n482), .ZN(n713) );
  INV_X1 U416 ( .A(KEYINPUT6), .ZN(n391) );
  XNOR2_X1 U417 ( .A(G119), .B(G116), .ZN(n447) );
  XNOR2_X1 U418 ( .A(n458), .B(n449), .ZN(n448) );
  INV_X1 U419 ( .A(KEYINPUT3), .ZN(n449) );
  INV_X1 U420 ( .A(KEYINPUT5), .ZN(n364) );
  XNOR2_X1 U421 ( .A(G104), .B(G110), .ZN(n462) );
  XNOR2_X1 U422 ( .A(G128), .B(G119), .ZN(n530) );
  XNOR2_X1 U423 ( .A(n529), .B(n531), .ZN(n385) );
  XNOR2_X1 U424 ( .A(G137), .B(G110), .ZN(n527) );
  INV_X1 U425 ( .A(KEYINPUT8), .ZN(n443) );
  XOR2_X1 U426 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n492) );
  XNOR2_X1 U427 ( .A(n491), .B(n382), .ZN(n381) );
  XOR2_X1 U428 ( .A(G122), .B(KEYINPUT12), .Z(n496) );
  INV_X1 U429 ( .A(KEYINPUT70), .ZN(n395) );
  XNOR2_X1 U430 ( .A(G143), .B(G104), .ZN(n417) );
  XNOR2_X1 U431 ( .A(n769), .B(G146), .ZN(n544) );
  XNOR2_X1 U432 ( .A(n639), .B(n399), .ZN(n398) );
  INV_X1 U433 ( .A(KEYINPUT108), .ZN(n399) );
  AND2_X1 U434 ( .A1(n605), .A2(n705), .ZN(n600) );
  XNOR2_X1 U435 ( .A(n535), .B(KEYINPUT96), .ZN(n536) );
  XNOR2_X1 U436 ( .A(n534), .B(KEYINPUT25), .ZN(n535) );
  OR2_X1 U437 ( .A1(n586), .A2(n426), .ZN(n425) );
  NAND2_X1 U438 ( .A1(n623), .A2(n427), .ZN(n426) );
  INV_X1 U439 ( .A(KEYINPUT73), .ZN(n413) );
  XNOR2_X1 U440 ( .A(n633), .B(KEYINPUT46), .ZN(n429) );
  INV_X1 U441 ( .A(KEYINPUT48), .ZN(n379) );
  NOR2_X1 U442 ( .A1(n685), .A2(n457), .ZN(n454) );
  OR2_X1 U443 ( .A1(n430), .A2(n379), .ZN(n377) );
  INV_X1 U444 ( .A(KEYINPUT84), .ZN(n380) );
  NOR2_X1 U445 ( .A1(n779), .A2(n578), .ZN(n418) );
  BUF_X1 U446 ( .A(n714), .Z(n414) );
  NOR2_X1 U447 ( .A1(n643), .A2(n683), .ZN(n717) );
  NAND2_X1 U448 ( .A1(n414), .A2(n713), .ZN(n434) );
  INV_X1 U449 ( .A(KEYINPUT15), .ZN(n475) );
  NOR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n476) );
  XOR2_X1 U451 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n503) );
  INV_X1 U452 ( .A(G902), .ZN(n545) );
  INV_X1 U453 ( .A(G953), .ZN(n755) );
  INV_X1 U454 ( .A(G134), .ZN(n396) );
  INV_X1 U455 ( .A(KEYINPUT45), .ZN(n411) );
  XNOR2_X1 U456 ( .A(KEYINPUT41), .B(n630), .ZN(n726) );
  AND2_X1 U457 ( .A1(n714), .A2(n432), .ZN(n630) );
  NOR2_X1 U458 ( .A1(n716), .A2(n433), .ZN(n432) );
  INV_X1 U459 ( .A(n713), .ZN(n433) );
  XNOR2_X1 U460 ( .A(n686), .B(KEYINPUT106), .ZN(n643) );
  XNOR2_X1 U461 ( .A(n416), .B(n415), .ZN(n709) );
  INV_X1 U462 ( .A(KEYINPUT100), .ZN(n415) );
  NOR2_X1 U463 ( .A1(n584), .A2(n585), .ZN(n416) );
  INV_X1 U464 ( .A(n619), .ZN(n620) );
  XNOR2_X1 U465 ( .A(n618), .B(n617), .ZN(n621) );
  NAND2_X1 U466 ( .A1(n614), .A2(KEYINPUT98), .ZN(n424) );
  INV_X1 U467 ( .A(KEYINPUT0), .ZN(n445) );
  XNOR2_X1 U468 ( .A(n543), .B(n544), .ZN(n657) );
  XNOR2_X1 U469 ( .A(n363), .B(n538), .ZN(n541) );
  XNOR2_X1 U470 ( .A(n540), .B(n364), .ZN(n363) );
  XNOR2_X1 U471 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U472 ( .A(n532), .B(n387), .ZN(n386) );
  XNOR2_X1 U473 ( .A(n530), .B(KEYINPUT93), .ZN(n384) );
  XNOR2_X1 U474 ( .A(n387), .B(n444), .ZN(n663) );
  XNOR2_X1 U475 ( .A(n522), .B(n417), .ZN(n494) );
  XNOR2_X1 U476 ( .A(n519), .B(n382), .ZN(n520) );
  XNOR2_X1 U477 ( .A(n362), .B(KEYINPUT43), .ZN(n397) );
  NOR2_X1 U478 ( .A1(n639), .A2(n641), .ZN(n611) );
  INV_X1 U479 ( .A(n631), .ZN(n390) );
  INV_X1 U480 ( .A(n686), .ZN(n438) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n567) );
  INV_X1 U482 ( .A(KEYINPUT85), .ZN(n419) );
  INV_X1 U483 ( .A(n683), .ZN(n437) );
  AND2_X2 U484 ( .A1(n556), .A2(n555), .ZN(n686) );
  XNOR2_X1 U485 ( .A(n485), .B(n484), .ZN(n603) );
  NAND2_X1 U486 ( .A1(n490), .A2(n697), .ZN(n352) );
  XOR2_X1 U487 ( .A(KEYINPUT13), .B(G475), .Z(n353) );
  XNOR2_X1 U488 ( .A(G478), .B(n512), .ZN(n574) );
  AND2_X1 U489 ( .A1(n397), .A2(n641), .ZN(n354) );
  AND2_X1 U490 ( .A1(n452), .A2(n456), .ZN(n355) );
  AND2_X1 U491 ( .A1(n377), .A2(n375), .ZN(n356) );
  INV_X1 U492 ( .A(n387), .ZN(n768) );
  AND2_X1 U493 ( .A1(n585), .A2(n424), .ZN(n357) );
  INV_X1 U494 ( .A(G140), .ZN(n382) );
  NOR2_X1 U495 ( .A1(n439), .A2(G900), .ZN(n358) );
  XNOR2_X1 U496 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n359) );
  INV_X1 U497 ( .A(KEYINPUT98), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n386), .B(n383), .ZN(n747) );
  OR2_X1 U499 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n361) );
  NAND2_X1 U500 ( .A1(n657), .A2(n545), .ZN(n546) );
  NAND2_X1 U501 ( .A1(n398), .A2(n640), .ZN(n362) );
  NAND2_X1 U502 ( .A1(n365), .A2(n578), .ZN(n580) );
  INV_X1 U503 ( .A(n779), .ZN(n365) );
  NAND2_X1 U504 ( .A1(n378), .A2(n377), .ZN(n376) );
  NAND2_X1 U505 ( .A1(n366), .A2(n356), .ZN(n370) );
  AND2_X1 U506 ( .A1(n367), .A2(n378), .ZN(n366) );
  NOR2_X1 U507 ( .A1(n780), .A2(n380), .ZN(n367) );
  NAND2_X1 U508 ( .A1(n368), .A2(n375), .ZN(n374) );
  OR2_X1 U509 ( .A1(n429), .A2(n379), .ZN(n375) );
  INV_X1 U510 ( .A(n780), .ZN(n368) );
  NAND2_X1 U511 ( .A1(n369), .A2(n430), .ZN(n378) );
  AND2_X1 U512 ( .A1(n429), .A2(n379), .ZN(n369) );
  NAND2_X1 U513 ( .A1(n371), .A2(n370), .ZN(n645) );
  NAND2_X1 U514 ( .A1(n376), .A2(n380), .ZN(n372) );
  NAND2_X1 U515 ( .A1(n374), .A2(n380), .ZN(n373) );
  NAND2_X1 U516 ( .A1(n388), .A2(KEYINPUT47), .ZN(n638) );
  INV_X1 U517 ( .A(n585), .ZN(n705) );
  NAND2_X1 U518 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U519 ( .A1(n405), .A2(n408), .ZN(n402) );
  NAND2_X1 U520 ( .A1(n403), .A2(KEYINPUT107), .ZN(n405) );
  NAND2_X1 U521 ( .A1(n410), .A2(n404), .ZN(n403) );
  INV_X1 U522 ( .A(n590), .ZN(n404) );
  NAND2_X1 U523 ( .A1(n435), .A2(n361), .ZN(n406) );
  NAND2_X1 U524 ( .A1(n583), .A2(n582), .ZN(n407) );
  NAND2_X1 U525 ( .A1(n410), .A2(n409), .ZN(n408) );
  NOR2_X1 U526 ( .A1(n590), .A2(KEYINPUT107), .ZN(n409) );
  INV_X1 U527 ( .A(n591), .ZN(n410) );
  NAND2_X1 U528 ( .A1(n412), .A2(n552), .ZN(n553) );
  NAND2_X1 U529 ( .A1(n412), .A2(n606), .ZN(n420) );
  NAND2_X1 U530 ( .A1(n412), .A2(n548), .ZN(n568) );
  NOR2_X2 U531 ( .A1(n598), .A2(n701), .ZN(n699) );
  NOR2_X2 U532 ( .A1(n423), .A2(n422), .ZN(n428) );
  INV_X1 U533 ( .A(n559), .ZN(n575) );
  XNOR2_X1 U534 ( .A(n593), .B(n413), .ZN(n441) );
  XNOR2_X1 U535 ( .A(n494), .B(n499), .ZN(n444) );
  NAND2_X1 U536 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U537 ( .A1(n581), .A2(n579), .ZN(n436) );
  XNOR2_X2 U538 ( .A(n577), .B(KEYINPUT35), .ZN(n779) );
  XNOR2_X2 U539 ( .A(n628), .B(n627), .ZN(n782) );
  BUF_X2 U540 ( .A(n624), .Z(n610) );
  NAND2_X1 U541 ( .A1(n436), .A2(n418), .ZN(n435) );
  NAND2_X1 U542 ( .A1(n440), .A2(n421), .ZN(n431) );
  NAND2_X1 U543 ( .A1(n645), .A2(n690), .ZN(n691) );
  AND2_X1 U544 ( .A1(n586), .A2(KEYINPUT98), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n425), .A2(n357), .ZN(n423) );
  XNOR2_X2 U546 ( .A(n446), .B(n445), .ZN(n586) );
  NOR2_X1 U547 ( .A1(n455), .A2(KEYINPUT102), .ZN(n450) );
  XNOR2_X2 U548 ( .A(n428), .B(KEYINPUT99), .ZN(n455) );
  NOR2_X2 U549 ( .A1(n431), .A2(n613), .ZN(n430) );
  NOR2_X1 U550 ( .A1(n717), .A2(n434), .ZN(n718) );
  OR2_X1 U551 ( .A1(n455), .A2(n437), .ZN(n558) );
  OR2_X1 U552 ( .A1(n455), .A2(n438), .ZN(n564) );
  NAND2_X1 U553 ( .A1(n439), .A2(G224), .ZN(n466) );
  NAND2_X1 U554 ( .A1(n439), .A2(G234), .ZN(n506) );
  NAND2_X1 U555 ( .A1(n439), .A2(G227), .ZN(n519) );
  OR2_X1 U556 ( .A1(n439), .A2(G952), .ZN(n666) );
  NAND2_X1 U557 ( .A1(n772), .A2(n439), .ZN(n778) );
  XNOR2_X2 U558 ( .A(n465), .B(G953), .ZN(n439) );
  NOR2_X2 U559 ( .A1(n567), .A2(n566), .ZN(n590) );
  NAND2_X1 U560 ( .A1(n685), .A2(n457), .ZN(n452) );
  NOR2_X2 U561 ( .A1(n782), .A2(n781), .ZN(n633) );
  INV_X1 U562 ( .A(n615), .ZN(n585) );
  NOR2_X2 U563 ( .A1(n726), .A2(n631), .ZN(n632) );
  NAND2_X1 U564 ( .A1(n441), .A2(n360), .ZN(n440) );
  NAND2_X1 U565 ( .A1(n442), .A2(G221), .ZN(n532) );
  NAND2_X1 U566 ( .A1(n442), .A2(G217), .ZN(n507) );
  XNOR2_X2 U567 ( .A(n506), .B(n443), .ZN(n442) );
  INV_X1 U568 ( .A(n714), .ZN(n629) );
  XNOR2_X2 U569 ( .A(n610), .B(n359), .ZN(n714) );
  NOR2_X2 U570 ( .A1(n603), .A2(n352), .ZN(n446) );
  XNOR2_X2 U571 ( .A(n448), .B(n447), .ZN(n542) );
  NOR2_X1 U572 ( .A1(n451), .A2(n450), .ZN(n591) );
  NAND2_X1 U573 ( .A1(n453), .A2(n355), .ZN(n451) );
  NAND2_X1 U574 ( .A1(n455), .A2(n454), .ZN(n453) );
  INV_X1 U575 ( .A(n592), .ZN(n456) );
  INV_X1 U576 ( .A(KEYINPUT102), .ZN(n457) );
  XNOR2_X2 U577 ( .A(KEYINPUT42), .B(n632), .ZN(n781) );
  BUF_X1 U578 ( .A(n669), .Z(n673) );
  INV_X1 U579 ( .A(n689), .ZN(n613) );
  INV_X1 U580 ( .A(KEYINPUT87), .ZN(n570) );
  XNOR2_X1 U581 ( .A(n570), .B(KEYINPUT33), .ZN(n571) );
  XNOR2_X1 U582 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U583 ( .A(n498), .B(n497), .ZN(n499) );
  NOR2_X1 U584 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n524) );
  BUF_X1 U586 ( .A(n691), .Z(n771) );
  INV_X1 U587 ( .A(KEYINPUT1), .ZN(n526) );
  INV_X1 U588 ( .A(n698), .ZN(n640) );
  INV_X1 U589 ( .A(KEYINPUT40), .ZN(n627) );
  XNOR2_X1 U590 ( .A(n459), .B(KEYINPUT72), .ZN(n460) );
  XNOR2_X2 U591 ( .A(n542), .B(n460), .ZN(n762) );
  INV_X1 U592 ( .A(G107), .ZN(n461) );
  XNOR2_X1 U593 ( .A(n462), .B(n461), .ZN(n760) );
  INV_X1 U594 ( .A(KEYINPUT68), .ZN(n463) );
  XNOR2_X1 U595 ( .A(n463), .B(G101), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n760), .B(n538), .ZN(n521) );
  XNOR2_X1 U597 ( .A(n762), .B(n521), .ZN(n474) );
  INV_X2 U598 ( .A(G146), .ZN(n464) );
  XNOR2_X2 U599 ( .A(n464), .B(G125), .ZN(n491) );
  XNOR2_X1 U600 ( .A(n491), .B(KEYINPUT4), .ZN(n468) );
  XNOR2_X1 U601 ( .A(n466), .B(n509), .ZN(n467) );
  XNOR2_X1 U602 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT80), .Z(n470) );
  XOR2_X1 U604 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n469) );
  XNOR2_X1 U605 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U606 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U607 ( .A(n474), .B(n473), .ZN(n669) );
  XNOR2_X1 U608 ( .A(n475), .B(G902), .ZN(n649) );
  OR2_X2 U609 ( .A1(n669), .A2(n649), .ZN(n481) );
  XNOR2_X1 U610 ( .A(n476), .B(KEYINPUT76), .ZN(n483) );
  INV_X1 U611 ( .A(G210), .ZN(n477) );
  OR2_X1 U612 ( .A1(n483), .A2(n477), .ZN(n479) );
  INV_X1 U613 ( .A(KEYINPUT90), .ZN(n478) );
  XNOR2_X1 U614 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X2 U615 ( .A(n481), .B(n480), .ZN(n624) );
  INV_X1 U616 ( .A(G214), .ZN(n482) );
  NAND2_X1 U617 ( .A1(n624), .A2(n713), .ZN(n485) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n484) );
  XNOR2_X1 U619 ( .A(G898), .B(KEYINPUT92), .ZN(n754) );
  NOR2_X1 U620 ( .A1(n755), .A2(n754), .ZN(n765) );
  NAND2_X1 U621 ( .A1(n765), .A2(G902), .ZN(n486) );
  NAND2_X1 U622 ( .A1(n755), .A2(G952), .ZN(n595) );
  NAND2_X1 U623 ( .A1(n486), .A2(n595), .ZN(n490) );
  XOR2_X1 U624 ( .A(KEYINPUT91), .B(KEYINPUT14), .Z(n489) );
  NAND2_X1 U625 ( .A1(G234), .A2(G237), .ZN(n487) );
  XNOR2_X1 U626 ( .A(n487), .B(KEYINPUT74), .ZN(n488) );
  XNOR2_X1 U627 ( .A(n489), .B(n488), .ZN(n697) );
  XNOR2_X1 U628 ( .A(G113), .B(KEYINPUT11), .ZN(n495) );
  XNOR2_X1 U629 ( .A(n496), .B(n495), .ZN(n498) );
  NOR2_X1 U630 ( .A1(G953), .A2(G237), .ZN(n539) );
  NAND2_X1 U631 ( .A1(G214), .A2(n539), .ZN(n497) );
  NAND2_X1 U632 ( .A1(n663), .A2(n545), .ZN(n500) );
  XNOR2_X1 U633 ( .A(G116), .B(G107), .ZN(n501) );
  XNOR2_X1 U634 ( .A(n501), .B(KEYINPUT9), .ZN(n505) );
  XNOR2_X1 U635 ( .A(G122), .B(KEYINPUT104), .ZN(n502) );
  XNOR2_X1 U636 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U637 ( .A(n505), .B(n504), .Z(n508) );
  XNOR2_X1 U638 ( .A(n508), .B(n507), .ZN(n511) );
  INV_X1 U639 ( .A(n523), .ZN(n510) );
  XNOR2_X1 U640 ( .A(n511), .B(n510), .ZN(n743) );
  NOR2_X1 U641 ( .A1(G902), .A2(n743), .ZN(n512) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n716) );
  XOR2_X1 U643 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n514) );
  INV_X1 U644 ( .A(n649), .ZN(n653) );
  NAND2_X1 U645 ( .A1(G234), .A2(n653), .ZN(n513) );
  XNOR2_X1 U646 ( .A(n514), .B(n513), .ZN(n533) );
  NAND2_X1 U647 ( .A1(n533), .A2(G221), .ZN(n517) );
  INV_X1 U648 ( .A(KEYINPUT97), .ZN(n515) );
  XNOR2_X1 U649 ( .A(n515), .B(KEYINPUT21), .ZN(n516) );
  XNOR2_X1 U650 ( .A(n517), .B(n516), .ZN(n701) );
  OR2_X1 U651 ( .A1(n716), .A2(n701), .ZN(n518) );
  XNOR2_X1 U652 ( .A(n544), .B(n524), .ZN(n739) );
  XOR2_X1 U653 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n528) );
  XNOR2_X1 U654 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U655 ( .A(KEYINPUT23), .B(KEYINPUT79), .Z(n531) );
  NAND2_X1 U656 ( .A1(G217), .A2(n533), .ZN(n534) );
  XNOR2_X2 U657 ( .A(n537), .B(n536), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n640), .A2(n598), .ZN(n547) );
  NAND2_X1 U659 ( .A1(n539), .A2(G210), .ZN(n540) );
  NOR2_X1 U660 ( .A1(n547), .A2(n705), .ZN(n548) );
  XNOR2_X1 U661 ( .A(n568), .B(G110), .ZN(G12) );
  INV_X1 U662 ( .A(KEYINPUT81), .ZN(n549) );
  XNOR2_X1 U663 ( .A(n606), .B(n549), .ZN(n551) );
  INV_X1 U664 ( .A(n598), .ZN(n565) );
  NOR2_X1 U665 ( .A1(n640), .A2(n565), .ZN(n550) );
  AND2_X1 U666 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X2 U667 ( .A(n553), .B(KEYINPUT32), .ZN(n569) );
  XNOR2_X1 U668 ( .A(n569), .B(G119), .ZN(G21) );
  INV_X1 U669 ( .A(n554), .ZN(n601) );
  NAND2_X1 U670 ( .A1(n601), .A2(n699), .ZN(n614) );
  XNOR2_X1 U671 ( .A(n559), .B(KEYINPUT103), .ZN(n556) );
  INV_X1 U672 ( .A(n574), .ZN(n555) );
  XOR2_X1 U673 ( .A(G104), .B(KEYINPUT113), .Z(n557) );
  XNOR2_X1 U674 ( .A(n558), .B(n557), .ZN(G6) );
  XOR2_X1 U675 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n561) );
  XNOR2_X1 U676 ( .A(G107), .B(KEYINPUT26), .ZN(n560) );
  XNOR2_X1 U677 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U678 ( .A(KEYINPUT114), .B(n562), .Z(n563) );
  XNOR2_X1 U679 ( .A(n564), .B(n563), .ZN(G9) );
  NAND2_X1 U680 ( .A1(n640), .A2(n565), .ZN(n566) );
  XOR2_X1 U681 ( .A(n590), .B(G101), .Z(G3) );
  INV_X1 U682 ( .A(KEYINPUT65), .ZN(n579) );
  NAND2_X1 U683 ( .A1(n699), .A2(n698), .ZN(n584) );
  XNOR2_X1 U684 ( .A(n573), .B(KEYINPUT34), .ZN(n576) );
  NOR2_X1 U685 ( .A1(n575), .A2(n574), .ZN(n636) );
  NAND2_X1 U686 ( .A1(n576), .A2(n636), .ZN(n577) );
  INV_X1 U687 ( .A(KEYINPUT44), .ZN(n578) );
  NAND2_X1 U688 ( .A1(n580), .A2(n579), .ZN(n583) );
  INV_X1 U689 ( .A(n581), .ZN(n582) );
  NOR2_X1 U690 ( .A1(n709), .A2(n586), .ZN(n588) );
  XNOR2_X1 U691 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n587) );
  INV_X1 U692 ( .A(KEYINPUT83), .ZN(n589) );
  XNOR2_X1 U693 ( .A(n717), .B(n589), .ZN(n592) );
  INV_X1 U694 ( .A(KEYINPUT2), .ZN(n652) );
  NOR2_X1 U695 ( .A1(n692), .A2(n652), .ZN(n647) );
  NOR2_X1 U696 ( .A1(n592), .A2(KEYINPUT47), .ZN(n593) );
  NAND2_X1 U697 ( .A1(G902), .A2(n358), .ZN(n594) );
  NAND2_X1 U698 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U699 ( .A1(n697), .A2(n596), .ZN(n597) );
  XOR2_X1 U700 ( .A(KEYINPUT82), .B(n597), .Z(n619) );
  NAND2_X1 U701 ( .A1(n598), .A2(n619), .ZN(n599) );
  NOR2_X2 U702 ( .A1(n701), .A2(n599), .ZN(n605) );
  XNOR2_X1 U703 ( .A(KEYINPUT28), .B(n600), .ZN(n602) );
  NAND2_X1 U704 ( .A1(n602), .A2(n601), .ZN(n631) );
  INV_X1 U705 ( .A(n603), .ZN(n604) );
  NAND2_X1 U706 ( .A1(n605), .A2(n683), .ZN(n609) );
  INV_X1 U707 ( .A(n606), .ZN(n607) );
  NAND2_X1 U708 ( .A1(n607), .A2(n713), .ZN(n608) );
  INV_X1 U709 ( .A(n610), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n611), .B(KEYINPUT36), .ZN(n612) );
  NAND2_X1 U711 ( .A1(n612), .A2(n698), .ZN(n689) );
  INV_X1 U712 ( .A(n614), .ZN(n623) );
  NAND2_X1 U713 ( .A1(n615), .A2(n713), .ZN(n618) );
  XOR2_X1 U714 ( .A(KEYINPUT30), .B(KEYINPUT111), .Z(n616) );
  NAND2_X1 U715 ( .A1(n623), .A2(n622), .ZN(n634) );
  INV_X1 U716 ( .A(KEYINPUT39), .ZN(n625) );
  XNOR2_X1 U717 ( .A(n626), .B(n625), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n644), .A2(n683), .ZN(n628) );
  NOR2_X1 U719 ( .A1(n634), .A2(n641), .ZN(n635) );
  XNOR2_X1 U720 ( .A(n635), .B(KEYINPUT112), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n680) );
  INV_X1 U722 ( .A(KEYINPUT109), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n354), .B(n642), .ZN(n780) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n690) );
  INV_X1 U725 ( .A(n691), .ZN(n646) );
  XNOR2_X2 U726 ( .A(n648), .B(KEYINPUT78), .ZN(n696) );
  XNOR2_X1 U727 ( .A(n691), .B(KEYINPUT77), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n655) );
  OR2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n654) );
  AND2_X2 U730 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X4 U731 ( .A1(n696), .A2(n656), .ZN(n735) );
  NAND2_X1 U732 ( .A1(n735), .A2(G472), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT62), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n660), .A2(n666), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U737 ( .A1(n735), .A2(G475), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n662) );
  XNOR2_X1 U739 ( .A(n665), .B(n664), .ZN(n667) );
  INV_X1 U740 ( .A(n666), .ZN(n750) );
  NOR2_X2 U741 ( .A1(n667), .A2(n750), .ZN(n668) );
  XNOR2_X1 U742 ( .A(n668), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U743 ( .A1(n735), .A2(G210), .ZN(n675) );
  XOR2_X1 U744 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n671) );
  XNOR2_X1 U745 ( .A(KEYINPUT55), .B(KEYINPUT86), .ZN(n670) );
  XNOR2_X1 U746 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U747 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X2 U748 ( .A1(n676), .A2(n750), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U750 ( .A(G128), .B(KEYINPUT29), .Z(n679) );
  NAND2_X1 U751 ( .A1(n360), .A2(n686), .ZN(n678) );
  XNOR2_X1 U752 ( .A(n679), .B(n678), .ZN(G30) );
  XNOR2_X1 U753 ( .A(G143), .B(KEYINPUT116), .ZN(n681) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(G45) );
  NAND2_X1 U755 ( .A1(n360), .A2(n683), .ZN(n682) );
  XNOR2_X1 U756 ( .A(n682), .B(G146), .ZN(G48) );
  NAND2_X1 U757 ( .A1(n683), .A2(n685), .ZN(n684) );
  XNOR2_X1 U758 ( .A(n684), .B(G113), .ZN(G15) );
  NAND2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(G116), .ZN(G18) );
  XOR2_X1 U761 ( .A(G125), .B(KEYINPUT37), .Z(n688) );
  XNOR2_X1 U762 ( .A(n689), .B(n688), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G134), .B(n690), .ZN(G36) );
  BUF_X1 U764 ( .A(n692), .Z(n693) );
  NOR2_X1 U765 ( .A1(n771), .A2(n693), .ZN(n694) );
  NOR2_X1 U766 ( .A1(n694), .A2(KEYINPUT2), .ZN(n695) );
  OR2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n733) );
  NAND2_X1 U768 ( .A1(G952), .A2(n697), .ZN(n725) );
  NOR2_X1 U769 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U770 ( .A(KEYINPUT50), .B(n700), .Z(n707) );
  XOR2_X1 U771 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n703) );
  NAND2_X1 U772 ( .A1(n701), .A2(n598), .ZN(n702) );
  XNOR2_X1 U773 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U775 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n710), .ZN(n711) );
  NOR2_X1 U778 ( .A1(n726), .A2(n711), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n712), .B(KEYINPUT118), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n414), .A2(n713), .ZN(n715) );
  NOR2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n719) );
  NOR2_X1 U782 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n727), .A2(n720), .ZN(n721) );
  NOR2_X1 U784 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U785 ( .A(n723), .B(KEYINPUT52), .ZN(n724) );
  NOR2_X1 U786 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U788 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U789 ( .A(n730), .B(KEYINPUT119), .ZN(n731) );
  NOR2_X1 U790 ( .A1(G953), .A2(n731), .ZN(n732) );
  NAND2_X1 U791 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U792 ( .A(KEYINPUT53), .B(n734), .Z(G75) );
  NAND2_X1 U793 ( .A1(n746), .A2(G469), .ZN(n741) );
  XOR2_X1 U794 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n737) );
  XNOR2_X1 U795 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n736) );
  XNOR2_X1 U796 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U797 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U798 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U799 ( .A1(n750), .A2(n742), .ZN(G54) );
  NAND2_X1 U800 ( .A1(n746), .A2(G478), .ZN(n744) );
  XNOR2_X1 U801 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U802 ( .A1(n750), .A2(n745), .ZN(G63) );
  NAND2_X1 U803 ( .A1(n746), .A2(G217), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n748), .B(n747), .ZN(n749) );
  NOR2_X1 U805 ( .A1(n750), .A2(n749), .ZN(G66) );
  XOR2_X1 U806 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n752) );
  NAND2_X1 U807 ( .A1(G224), .A2(G953), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n752), .B(n751), .ZN(n753) );
  NAND2_X1 U809 ( .A1(n754), .A2(n753), .ZN(n759) );
  NAND2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(KEYINPUT124), .ZN(n758) );
  NAND2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n767) );
  XOR2_X1 U813 ( .A(KEYINPUT125), .B(n760), .Z(n761) );
  XNOR2_X1 U814 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(G101), .ZN(n764) );
  NOR2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n767), .B(n766), .ZN(G69) );
  XNOR2_X1 U818 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U819 ( .A(n770), .B(KEYINPUT126), .ZN(n773) );
  XNOR2_X1 U820 ( .A(n771), .B(n773), .ZN(n772) );
  XNOR2_X1 U821 ( .A(G227), .B(n773), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n775), .A2(G953), .ZN(n776) );
  XOR2_X1 U824 ( .A(KEYINPUT127), .B(n776), .Z(n777) );
  NAND2_X1 U825 ( .A1(n778), .A2(n777), .ZN(G72) );
  XOR2_X1 U826 ( .A(G122), .B(n779), .Z(G24) );
  XOR2_X1 U827 ( .A(n780), .B(G140), .Z(G42) );
  XOR2_X1 U828 ( .A(n781), .B(G137), .Z(G39) );
  XOR2_X1 U829 ( .A(n782), .B(G131), .Z(G33) );
endmodule

