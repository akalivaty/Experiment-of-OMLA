//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882;
  INV_X1    g000(.A(KEYINPUT107), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT95), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT36), .ZN(new_n204));
  OR2_X1    g003(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(KEYINPUT28), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(new_n206), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(new_n210), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  OR3_X1    g019(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(new_n220), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n228), .B(new_n232), .C1(new_n230), .C2(new_n231), .ZN(new_n233));
  OR3_X1    g032(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n234), .A2(new_n235), .B1(G169gat), .B2(G176gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n236), .B(new_n239), .C1(new_n229), .C2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n238), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n243));
  INV_X1    g042(.A(G120gat), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G113gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n245), .A2(G120gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n243), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(G134gat), .ZN(new_n254));
  NOR3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT1), .ZN(new_n255));
  INV_X1    g054(.A(new_n250), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT69), .B(G113gat), .ZN(new_n257));
  OAI211_X1 g056(.A(KEYINPUT70), .B(new_n256), .C1(new_n257), .C2(new_n244), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n252), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G113gat), .B(G120gat), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n262), .A2(new_n253), .B1(KEYINPUT1), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n242), .B(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G227gat), .A2(G233gat), .ZN(new_n267));
  OR2_X1    g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT72), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n267), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n274), .B2(KEYINPUT32), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n271), .B(new_n273), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n278), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n268), .A2(new_n269), .A3(new_n272), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n272), .B1(new_n268), .B2(new_n269), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n280), .B(new_n276), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT33), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n274), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n279), .A2(new_n283), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n279), .B2(new_n283), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n204), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n283), .ZN(new_n294));
  INV_X1    g093(.A(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT36), .A3(new_n290), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G57gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G85gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G1gat), .B(G29gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G141gat), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n309), .A2(new_n311), .B1(KEYINPUT2), .B2(new_n306), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n313), .A3(new_n307), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n259), .A2(new_n315), .A3(new_n316), .A4(new_n264), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT76), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n316), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n320), .A2(new_n314), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(KEYINPUT76), .A3(new_n264), .A4(new_n259), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n317), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n315), .A2(new_n316), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n330), .A3(new_n265), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n326), .B1(new_n331), .B2(KEYINPUT4), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT5), .ZN(new_n334));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n335), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT77), .B1(new_n338), .B2(new_n324), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n340), .B(KEYINPUT4), .C1(new_n319), .C2(new_n322), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n324), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n337), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n265), .A2(new_n329), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n319), .A2(new_n322), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n335), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(KEYINPUT78), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT78), .B1(new_n347), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT5), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n302), .B(new_n336), .C1(new_n345), .C2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n347), .A2(new_n348), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n334), .B1(new_n358), .B2(new_n349), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n339), .A2(new_n341), .A3(new_n343), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n361), .A2(KEYINPUT79), .A3(new_n302), .A4(new_n336), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT6), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n336), .B1(new_n345), .B2(new_n352), .ZN(new_n366));
  INV_X1    g165(.A(new_n302), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n355), .A2(new_n368), .A3(new_n365), .A4(new_n362), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n242), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(KEYINPUT73), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT22), .ZN(new_n382));
  XOR2_X1   g181(.A(G211gat), .B(G218gat), .Z(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  INV_X1    g184(.A(G218gat), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT22), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n386), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n381), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT74), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n242), .A2(new_n391), .A3(new_n378), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n242), .B2(new_n378), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n380), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n390), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n242), .A2(new_n378), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n378), .B1(new_n242), .B2(new_n375), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G64gat), .ZN(new_n401));
  INV_X1    g200(.A(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n374), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n399), .A2(new_n403), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n373), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n395), .B2(KEYINPUT81), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n384), .A2(KEYINPUT81), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT3), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n409), .B1(new_n412), .B2(new_n321), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n390), .B1(new_n328), .B2(new_n375), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT3), .B1(new_n390), .B2(new_n375), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n321), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n413), .A2(new_n414), .B1(new_n417), .B2(new_n409), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT31), .B(G50gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  XOR2_X1   g219(.A(G78gat), .B(G106gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G22gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n420), .B(new_n422), .Z(new_n423));
  AOI21_X1  g222(.A(new_n298), .B1(new_n408), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n302), .B(KEYINPUT82), .Z(new_n425));
  NAND2_X1  g224(.A1(new_n366), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n355), .A2(new_n426), .A3(new_n365), .A4(new_n362), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n396), .A2(new_n397), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n390), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n380), .B1(new_n392), .B2(new_n393), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n395), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n428), .A2(KEYINPUT84), .A3(new_n390), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT38), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n394), .A2(new_n438), .A3(new_n398), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n436), .A2(new_n437), .A3(new_n403), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n399), .A2(KEYINPUT37), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n441), .A2(new_n403), .A3(new_n439), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n405), .B1(new_n442), .B2(KEYINPUT38), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n440), .A3(new_n370), .A4(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n348), .B1(new_n325), .B2(new_n332), .ZN(new_n445));
  OR2_X1    g244(.A1(new_n445), .A2(KEYINPUT39), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n323), .A2(new_n335), .A3(new_n346), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n448), .B2(KEYINPUT83), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n449), .B(new_n445), .C1(KEYINPUT83), .C2(new_n448), .ZN(new_n450));
  INV_X1    g249(.A(new_n425), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n446), .A2(new_n450), .A3(KEYINPUT40), .A4(new_n451), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n406), .A2(new_n426), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n423), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n444), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n444), .A2(new_n456), .A3(KEYINPUT85), .A4(new_n457), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n423), .B1(new_n296), .B2(new_n290), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n373), .A2(new_n407), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT35), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n427), .A2(new_n370), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n466), .B1(new_n467), .B2(new_n406), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n406), .B1(new_n427), .B2(new_n370), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT35), .B1(new_n469), .B2(KEYINPUT86), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n463), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n424), .A2(new_n462), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(KEYINPUT91), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n475), .A2(G1gat), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n476), .B2(KEYINPUT92), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT16), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n478), .B2(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n477), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n485), .A2(new_n487), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n487), .B2(new_n485), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(KEYINPUT15), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT15), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n487), .A2(new_n482), .B1(G29gat), .B2(G36gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n498), .B(KEYINPUT93), .Z(new_n499));
  NAND2_X1  g298(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(KEYINPUT90), .A2(KEYINPUT17), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n481), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT18), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n499), .B1(new_n481), .B2(new_n497), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n507), .B(KEYINPUT94), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(KEYINPUT13), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(KEYINPUT18), .A3(new_n507), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n510), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT11), .B(G169gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G197gat), .ZN(new_n518));
  XOR2_X1   g317(.A(G113gat), .B(G141gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT12), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n516), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n203), .B1(new_n472), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n460), .A2(new_n461), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n457), .B1(new_n373), .B2(new_n407), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n526), .A2(new_n527), .A3(new_n298), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n468), .A2(new_n463), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n529), .A2(new_n470), .B1(new_n464), .B2(KEYINPUT35), .ZN(new_n530));
  OAI211_X1 g329(.A(KEYINPUT95), .B(new_n523), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g333(.A(G99gat), .ZN(new_n535));
  INV_X1    g334(.A(G106gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT8), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT99), .B(G85gat), .Z(new_n538));
  OAI211_X1 g337(.A(new_n534), .B(new_n537), .C1(G92gat), .C2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G99gat), .B(G106gat), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n539), .B(new_n540), .Z(new_n541));
  NAND2_X1  g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  OR2_X1    g341(.A1(G71gat), .A2(G78gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT96), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n542), .B(new_n543), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n544), .B(KEYINPUT97), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n543), .B2(new_n546), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT101), .B1(new_n541), .B2(new_n551), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT10), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n555), .B1(new_n554), .B2(new_n553), .ZN(new_n556));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n558), .B(KEYINPUT102), .Z(new_n559));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n224), .ZN(new_n561));
  INV_X1    g360(.A(G204gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n552), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n541), .A2(new_n551), .ZN(new_n566));
  OAI211_X1 g365(.A(G230gat), .B(G233gat), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT103), .Z(new_n568));
  NAND3_X1  g367(.A1(new_n559), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n558), .B(KEYINPUT104), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n568), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n563), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n572), .A2(KEYINPUT105), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n572), .A2(KEYINPUT105), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT106), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT106), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n569), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n504), .B1(new_n580), .B2(new_n551), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n227), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT98), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n551), .A2(new_n580), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(new_n385), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n588), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n587), .B(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n503), .A2(new_n541), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n541), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n497), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT100), .ZN(new_n597));
  XOR2_X1   g396(.A(G190gat), .B(G218gat), .Z(new_n598));
  OAI211_X1 g397(.A(new_n594), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n597), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NOR3_X1   g404(.A1(new_n579), .A2(new_n592), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n202), .B1(new_n532), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n605), .ZN(new_n608));
  INV_X1    g407(.A(new_n579), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI211_X1 g409(.A(KEYINPUT107), .B(new_n610), .C1(new_n525), .C2(new_n531), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n373), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G1gat), .ZN(G1324gat));
  INV_X1    g415(.A(KEYINPUT108), .ZN(new_n617));
  XOR2_X1   g416(.A(KEYINPUT16), .B(G8gat), .Z(new_n618));
  OAI211_X1 g417(.A(new_n406), .B(new_n618), .C1(new_n607), .C2(new_n611), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT42), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n408), .A2(new_n423), .ZN(new_n622));
  INV_X1    g421(.A(new_n298), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n460), .A4(new_n461), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n465), .A2(new_n471), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT95), .B1(new_n626), .B2(new_n523), .ZN(new_n627));
  AOI211_X1 g426(.A(new_n203), .B(new_n524), .C1(new_n624), .C2(new_n625), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n606), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT107), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n532), .A2(new_n202), .A3(new_n606), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n407), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n632), .A2(KEYINPUT108), .A3(KEYINPUT42), .A4(new_n618), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n621), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n632), .B2(new_n473), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n619), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT109), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(new_n636), .A3(KEYINPUT109), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(G1325gat));
  NAND3_X1  g440(.A1(new_n613), .A2(G15gat), .A3(new_n298), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n291), .A2(new_n292), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n612), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n642), .B1(new_n644), .B2(G15gat), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n612), .A2(new_n457), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT43), .B(G22gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT110), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n647), .B(new_n649), .ZN(G1327gat));
  INV_X1    g449(.A(new_n592), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n579), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n532), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n605), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(G29gat), .A3(new_n373), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT45), .Z(new_n656));
  INV_X1    g455(.A(new_n605), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n472), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n660), .A2(new_n523), .A3(new_n652), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n661), .A2(KEYINPUT111), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(KEYINPUT111), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n373), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n665), .ZN(G1328gat));
  OAI21_X1  g465(.A(G36gat), .B1(new_n664), .B2(new_n407), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n654), .A2(G36gat), .A3(new_n407), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT46), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n668), .A2(KEYINPUT46), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(G1329gat));
  NOR3_X1   g470(.A1(new_n654), .A2(G43gat), .A3(new_n643), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G43gat), .B1(new_n661), .B2(new_n623), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(KEYINPUT47), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n298), .B1(new_n662), .B2(new_n663), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n672), .B1(new_n676), .B2(G43gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g477(.A1(new_n654), .A2(G50gat), .A3(new_n457), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G50gat), .B1(new_n661), .B2(new_n457), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(KEYINPUT48), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n423), .B1(new_n662), .B2(new_n663), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n679), .B1(new_n683), .B2(G50gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g484(.A1(new_n626), .A2(new_n524), .A3(new_n608), .A4(new_n579), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n373), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n407), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n689), .B2(new_n690), .ZN(G1333gat));
  OAI21_X1  g492(.A(G71gat), .B1(new_n686), .B2(new_n623), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n686), .A2(G71gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n695), .B2(new_n643), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT112), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g497(.A1(new_n686), .A2(new_n457), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n699), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g499(.A1(new_n651), .A2(new_n523), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n660), .A2(new_n579), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n538), .B1(new_n706), .B2(new_n373), .ZN(new_n707));
  INV_X1    g506(.A(new_n538), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n658), .A2(new_n701), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT51), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT114), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n658), .A2(KEYINPUT51), .A3(new_n701), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n712), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(KEYINPUT115), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(KEYINPUT115), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n708), .B(new_n579), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n707), .B1(new_n719), .B2(new_n373), .ZN(G1336gat));
  OAI21_X1  g519(.A(G92gat), .B1(new_n702), .B2(new_n407), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n609), .A2(G92gat), .A3(new_n407), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n721), .B(new_n722), .C1(new_n716), .C2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n406), .B1(new_n704), .B2(new_n705), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n713), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n726), .A2(G92gat), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n722), .ZN(G1337gat));
  OAI21_X1  g528(.A(G99gat), .B1(new_n706), .B2(new_n623), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n579), .B1(new_n717), .B2(new_n718), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n535), .B1(new_n291), .B2(new_n292), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(G1338gat));
  NOR3_X1   g532(.A1(new_n609), .A2(G106gat), .A3(new_n457), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n423), .B1(new_n704), .B2(new_n705), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(G106gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  OAI21_X1  g539(.A(G106gat), .B1(new_n702), .B2(new_n457), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n714), .A2(new_n715), .A3(new_n734), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n740), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT117), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(KEYINPUT117), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n739), .A2(new_n740), .B1(new_n744), .B2(new_n745), .ZN(G1339gat));
  INV_X1    g545(.A(new_n569), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n570), .A2(KEYINPUT54), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n564), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n559), .B(KEYINPUT54), .C1(new_n557), .C2(new_n556), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(KEYINPUT55), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(KEYINPUT55), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n747), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n516), .A2(new_n522), .ZN(new_n755));
  OAI22_X1  g554(.A1(new_n506), .A2(new_n507), .B1(new_n511), .B2(new_n513), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n520), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n657), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n579), .A2(new_n757), .B1(new_n754), .B2(new_n523), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(new_n657), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n760), .A2(new_n592), .B1(new_n524), .B2(new_n606), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n761), .A2(new_n643), .A3(new_n423), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n373), .A2(new_n406), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n523), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G113gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n257), .B2(new_n764), .ZN(G1340gat));
  NAND2_X1  g565(.A1(new_n762), .A2(new_n763), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n609), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(new_n244), .ZN(G1341gat));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n592), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n252), .ZN(G1342gat));
  NOR2_X1   g570(.A1(new_n767), .A2(new_n657), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n260), .A2(new_n261), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(KEYINPUT118), .B1(new_n774), .B2(KEYINPUT56), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n772), .A2(new_n776), .A3(new_n777), .A4(new_n773), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(KEYINPUT56), .ZN(new_n779));
  OAI21_X1  g578(.A(G134gat), .B1(new_n767), .B2(new_n657), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n775), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(G1343gat));
  OR2_X1    g580(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n623), .A2(new_n763), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT119), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n759), .A2(new_n657), .ZN(new_n785));
  INV_X1    g584(.A(new_n758), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n592), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n606), .A2(new_n524), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT57), .B1(new_n789), .B2(new_n423), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n791), .B(new_n457), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n523), .B(new_n784), .C1(new_n790), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G141gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n423), .ZN(new_n796));
  NOR4_X1   g595(.A1(new_n796), .A2(G141gat), .A3(new_n524), .A4(new_n783), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AND4_X1   g597(.A1(new_n782), .A2(new_n794), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n797), .B1(new_n793), .B2(G141gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n782), .B1(new_n800), .B2(new_n795), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(G1344gat));
  AOI21_X1  g601(.A(new_n457), .B1(new_n787), .B2(new_n788), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT57), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n791), .B1(new_n761), .B2(new_n457), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n807), .A3(new_n579), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n807), .A2(new_n308), .A3(KEYINPUT121), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n784), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT122), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n804), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n790), .A2(KEYINPUT122), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n579), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n784), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT59), .B(G148gat), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n796), .A2(new_n783), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n807), .B1(new_n819), .B2(new_n579), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n811), .B(new_n818), .C1(G148gat), .C2(new_n820), .ZN(G1345gat));
  INV_X1    g620(.A(new_n783), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n651), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n803), .A2(KEYINPUT123), .A3(new_n651), .A4(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n303), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n806), .A2(G155gat), .A3(new_n651), .A4(new_n784), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(G1346gat));
  AOI21_X1  g630(.A(G162gat), .B1(new_n819), .B2(new_n605), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n806), .A2(new_n784), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n657), .A2(new_n304), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(G1347gat));
  INV_X1    g634(.A(KEYINPUT126), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n614), .A2(new_n407), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n762), .A2(new_n523), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n223), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n836), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n836), .A3(new_n840), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(KEYINPUT125), .A3(G169gat), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n843), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n845), .A2(new_n841), .B1(new_n839), .B2(new_n223), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1348gat));
  NAND2_X1  g646(.A1(new_n762), .A2(new_n837), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n609), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(new_n224), .ZN(G1349gat));
  INV_X1    g649(.A(KEYINPUT127), .ZN(new_n851));
  OAI21_X1  g650(.A(G183gat), .B1(new_n848), .B2(new_n592), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n762), .A2(new_n214), .A3(new_n651), .A4(new_n837), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n851), .B(KEYINPUT60), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n851), .A2(KEYINPUT60), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n851), .A2(KEYINPUT60), .ZN(new_n856));
  AND4_X1   g655(.A1(new_n855), .A2(new_n852), .A3(new_n856), .A4(new_n853), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(new_n857), .ZN(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n848), .B2(new_n657), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(KEYINPUT61), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT61), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n848), .A2(new_n657), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n213), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n859), .B2(new_n863), .ZN(G1351gat));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n623), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n796), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(G197gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n523), .ZN(new_n868));
  INV_X1    g667(.A(new_n865), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n523), .A2(new_n813), .A3(new_n814), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n870), .B2(new_n867), .ZN(G1352gat));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n562), .A3(new_n579), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT62), .Z(new_n873));
  OAI21_X1  g672(.A(G204gat), .B1(new_n815), .B2(new_n865), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1353gat));
  NAND3_X1  g674(.A1(new_n866), .A2(new_n385), .A3(new_n651), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n813), .A2(new_n814), .A3(new_n651), .A4(new_n869), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT63), .B1(new_n877), .B2(G211gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(G1354gat));
  NAND3_X1  g679(.A1(new_n866), .A2(new_n386), .A3(new_n605), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n605), .A2(new_n813), .A3(new_n814), .A4(new_n869), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n882), .B2(new_n386), .ZN(G1355gat));
endmodule


