//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT31), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(G211gat), .B(G218gat), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT70), .ZN(new_n207));
  AND2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G197gat), .B(G204gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n211), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(KEYINPUT70), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n214), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(new_n205), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT71), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n210), .A2(new_n207), .A3(new_n211), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT70), .B1(new_n213), .B2(new_n214), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n205), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT71), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  INV_X1    g024(.A(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G141gat), .ZN(new_n227));
  INV_X1    g026(.A(G141gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G155gat), .B(G162gat), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(new_n228), .B2(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n228), .A2(G148gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n226), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G155gat), .ZN(new_n238));
  INV_X1    g037(.A(G162gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n225), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n232), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n219), .A2(new_n224), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n243), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n206), .A2(new_n213), .A3(new_n214), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n205), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT29), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n249), .B1(new_n252), .B2(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT78), .ZN(new_n255));
  INV_X1    g054(.A(G228gat), .ZN(new_n256));
  INV_X1    g055(.A(G233gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n249), .A2(KEYINPUT75), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT75), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n232), .B2(new_n243), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n223), .B1(new_n222), .B2(new_n250), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n216), .A2(KEYINPUT71), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n246), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n262), .B1(new_n265), .B2(new_n244), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n219), .A2(new_n224), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n245), .A2(KEYINPUT79), .A3(new_n246), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT79), .B1(new_n245), .B2(new_n246), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n255), .B(new_n258), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT80), .ZN(new_n272));
  INV_X1    g071(.A(new_n254), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n273), .A2(KEYINPUT78), .B1(new_n256), .B2(new_n257), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n271), .A2(new_n272), .A3(new_n274), .A4(G22gat), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n271), .A2(G22gat), .A3(new_n274), .ZN(new_n276));
  AOI21_X1  g075(.A(G22gat), .B1(new_n271), .B2(new_n274), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n204), .B(new_n275), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(G22gat), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n204), .A2(KEYINPUT80), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT81), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT81), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n278), .A2(new_n282), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT65), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n296), .A2(KEYINPUT65), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n292), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n296), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n294), .B2(new_n293), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT25), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n291), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT67), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT26), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT67), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n311), .A3(new_n291), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G183gat), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT27), .B1(new_n314), .B2(KEYINPUT66), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT27), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT27), .B(G183gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n321), .A2(G190gat), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n313), .B(new_n294), .C1(new_n322), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n330), .ZN(new_n333));
  INV_X1    g132(.A(G127gat), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n334), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n328), .B2(KEYINPUT68), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n305), .A2(new_n326), .A3(new_n337), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT34), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345));
  XNOR2_X1  g144(.A(G15gat), .B(G43gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G71gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G99gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n348), .B2(KEYINPUT69), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n349), .B1(KEYINPUT69), .B2(new_n348), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n342), .B(KEYINPUT64), .Z(new_n351));
  OAI211_X1 g150(.A(KEYINPUT32), .B(new_n350), .C1(new_n341), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n348), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n339), .B2(new_n340), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n345), .A2(KEYINPUT32), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT34), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n357), .A3(new_n351), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n344), .A2(new_n352), .A3(new_n356), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n344), .A2(new_n358), .B1(new_n352), .B2(new_n356), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n284), .A2(KEYINPUT35), .A3(new_n286), .A4(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n361), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(KEYINPUT36), .A3(new_n359), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT36), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n360), .B2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n278), .A2(new_n282), .A3(new_n285), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n285), .B1(new_n278), .B2(new_n282), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT3), .B1(new_n259), .B2(new_n261), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n338), .A3(new_n245), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n375), .B(KEYINPUT76), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n232), .A2(new_n243), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n337), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT4), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n337), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n374), .A2(new_n377), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n385), .A2(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n379), .B1(new_n262), .B2(new_n337), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n388), .B2(new_n376), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(new_n260), .ZN(new_n391));
  INV_X1    g190(.A(new_n261), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n337), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n379), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n376), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n384), .A3(new_n386), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G57gat), .ZN(new_n401));
  INV_X1    g200(.A(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT6), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n403), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n390), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n404), .B(new_n406), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n320), .A2(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n409));
  INV_X1    g208(.A(new_n294), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n300), .A2(new_n304), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT72), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n305), .A2(new_n326), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n327), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n267), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n327), .A2(new_n416), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n413), .A2(new_n415), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n421), .B1(new_n424), .B2(new_n267), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  INV_X1    g225(.A(G64gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  OR2_X1    g233(.A1(new_n425), .A2(new_n431), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n425), .A2(new_n431), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT73), .B1(new_n436), .B2(KEYINPUT30), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT73), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n432), .A2(new_n438), .A3(new_n433), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n434), .B(new_n435), .C1(new_n437), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n372), .A2(new_n407), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n406), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n390), .A2(KEYINPUT82), .A3(new_n397), .A4(new_n405), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n374), .A2(new_n383), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n376), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(KEYINPUT39), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(new_n405), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n448), .B(KEYINPUT39), .C1(new_n376), .C2(new_n388), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT40), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT40), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n446), .A3(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(KEYINPUT37), .B(new_n421), .C1(new_n424), .C2(new_n267), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n430), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(KEYINPUT85), .A3(new_n430), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT83), .B1(new_n425), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n425), .A2(KEYINPUT83), .A3(new_n463), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n461), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT38), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n432), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n446), .A2(new_n404), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n397), .A4(new_n405), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n463), .B1(new_n424), .B2(new_n267), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n418), .A2(new_n420), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n219), .A3(new_n224), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n431), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n472), .B(new_n476), .C1(new_n465), .C2(new_n464), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n469), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n457), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n369), .A2(new_n370), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n480), .A3(new_n368), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n469), .A2(new_n471), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n483), .A2(new_n284), .A3(new_n286), .A4(new_n362), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n482), .B1(new_n484), .B2(new_n440), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n442), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G1gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT16), .ZN(new_n488));
  INV_X1    g287(.A(G15gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(G22gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G15gat), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(G1gat), .B1(new_n490), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g293(.A(G8gat), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n491), .A2(G15gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n489), .A2(G22gat), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n488), .A2(new_n490), .A3(new_n492), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G71gat), .A2(G78gat), .ZN(new_n503));
  INV_X1    g302(.A(G71gat), .ZN(new_n504));
  INV_X1    g303(.A(G78gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n503), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G57gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G64gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n427), .A2(G57gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n503), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n503), .A2(new_n508), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n502), .B1(new_n517), .B2(KEYINPUT21), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT93), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT19), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(G127gat), .B(G155gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT20), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n524), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n517), .A2(KEYINPUT21), .ZN(new_n527));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n527), .B(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n525), .B2(new_n526), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G162gat), .B(G218gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G50gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G43gat), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G50gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT15), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT14), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT14), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT86), .ZN(new_n548));
  NAND2_X1  g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT86), .B1(new_n545), .B2(new_n547), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n542), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n538), .A2(new_n540), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n545), .A2(new_n547), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n541), .A4(new_n549), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n552), .A2(KEYINPUT17), .A3(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT7), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(G85gat), .A3(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n402), .B2(new_n429), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(G99gat), .ZN(new_n570));
  INV_X1    g369(.A(G106gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n567), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n576), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n573), .B1(new_n566), .B2(new_n568), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n558), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(G134gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(G134gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G190gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n585), .B2(new_n586), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n536), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n535), .A3(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n534), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n552), .A2(new_n495), .A3(new_n501), .A4(new_n557), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT89), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n558), .A2(new_n502), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n493), .A2(new_n494), .A3(G8gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n499), .B1(new_n498), .B2(new_n500), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT89), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n552), .A4(new_n557), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G229gat), .A2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT13), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT90), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n609), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(G197gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT11), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G169gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(G169gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n623), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT12), .A3(new_n621), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n560), .A2(new_n606), .A3(new_n561), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n603), .A2(KEYINPUT88), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n560), .A2(KEYINPUT88), .A3(new_n606), .A4(new_n561), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(KEYINPUT18), .A3(new_n610), .A4(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n610), .A3(new_n631), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT18), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n627), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT91), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n609), .A2(new_n614), .A3(new_n611), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n614), .B1(new_n609), .B2(new_n611), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n632), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n640), .B1(new_n616), .B2(new_n632), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT92), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT92), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n648), .B(new_n639), .C1(new_n644), .C2(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n638), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n600), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G176gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G204gat), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n509), .A2(new_n516), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n577), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n572), .A2(KEYINPUT96), .A3(new_n567), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n566), .A2(new_n658), .A3(new_n568), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n568), .B2(new_n566), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT95), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n582), .B2(new_n517), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n656), .B(KEYINPUT95), .C1(new_n581), .C2(new_n580), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n657), .B1(new_n665), .B2(new_n655), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT97), .Z(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n665), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n654), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n661), .ZN(new_n672));
  INV_X1    g471(.A(new_n664), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT95), .B1(new_n577), .B2(new_n656), .ZN(new_n674));
  OAI211_X1 g473(.A(new_n655), .B(new_n672), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n657), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n675), .A2(new_n676), .B1(G230gat), .B2(G233gat), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n677), .A2(new_n670), .A3(new_n654), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n486), .A2(new_n651), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n407), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n487), .ZN(G1324gat));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n441), .ZN(new_n684));
  OR2_X1    g483(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n684), .A2(KEYINPUT42), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(KEYINPUT98), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n684), .B2(new_n499), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n688), .B1(new_n692), .B2(new_n687), .ZN(G1325gat));
  INV_X1    g492(.A(new_n362), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n489), .B1(new_n681), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT99), .Z(new_n696));
  NOR3_X1   g495(.A1(new_n681), .A2(new_n489), .A3(new_n368), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n480), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND2_X1  g500(.A1(new_n486), .A2(new_n598), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n486), .A2(new_n704), .A3(new_n598), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n534), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(new_n650), .A3(new_n679), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G29gat), .B1(new_n709), .B2(new_n407), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n486), .A2(new_n543), .A3(new_n598), .A4(new_n708), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n711), .A2(KEYINPUT100), .A3(new_n407), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT100), .B1(new_n711), .B2(new_n407), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1328gat));
  AND2_X1   g518(.A1(new_n486), .A2(new_n598), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n708), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(G36gat), .A3(new_n441), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT46), .ZN(new_n723));
  OAI21_X1  g522(.A(G36gat), .B1(new_n709), .B2(new_n441), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1329gat));
  OAI21_X1  g524(.A(new_n539), .B1(new_n721), .B2(new_n694), .ZN(new_n726));
  INV_X1    g525(.A(new_n368), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G43gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n709), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g529(.A(new_n480), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n706), .A2(new_n731), .A3(new_n708), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT102), .B1(new_n732), .B2(G50gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n721), .A2(G50gat), .A3(new_n480), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n732), .B2(G50gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n735), .B(new_n737), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n599), .A2(new_n650), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n486), .A2(new_n679), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n407), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT103), .B(G57gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1332gat));
  AOI211_X1 g543(.A(new_n441), .B(new_n741), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(new_n504), .B1(new_n741), .B2(new_n694), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n727), .A2(G71gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g550(.A1(new_n741), .A2(new_n480), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n505), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n650), .A2(new_n534), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT104), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n486), .A2(new_n755), .A3(new_n598), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n759));
  INV_X1    g558(.A(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n756), .A2(new_n762), .A3(new_n757), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n407), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n766), .A2(new_n402), .A3(new_n767), .A4(new_n679), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n486), .A2(new_n704), .A3(new_n598), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n704), .B1(new_n486), .B2(new_n598), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n679), .B(new_n755), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n407), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1336gat));
  OAI21_X1  g572(.A(G92gat), .B1(new_n771), .B2(new_n441), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n441), .A2(G92gat), .A3(new_n680), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n760), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n756), .B1(new_n779), .B2(new_n757), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g580(.A(KEYINPUT107), .B(G92gat), .C1(new_n771), .C2(new_n441), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n771), .B2(new_n441), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n680), .B1(new_n703), .B2(new_n705), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(KEYINPUT109), .A3(new_n440), .A4(new_n755), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n788), .A3(G92gat), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n764), .B2(new_n777), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n784), .B1(new_n792), .B2(new_n793), .ZN(G1337gat));
  NAND4_X1  g593(.A1(new_n766), .A2(new_n570), .A3(new_n679), .A4(new_n362), .ZN(new_n795));
  OAI21_X1  g594(.A(G99gat), .B1(new_n771), .B2(new_n368), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(new_n771), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n571), .B1(new_n799), .B2(new_n731), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n778), .A2(new_n780), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n731), .A2(new_n571), .A3(new_n679), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT111), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n764), .A2(new_n804), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n798), .A2(new_n805), .B1(new_n806), .B2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n675), .A2(new_n668), .A3(new_n676), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n812), .B2(new_n677), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n675), .A2(new_n676), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n667), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n815), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n811), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n666), .A2(KEYINPUT54), .A3(new_n668), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n813), .A2(new_n816), .A3(new_n654), .A4(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(KEYINPUT113), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n678), .B1(new_n818), .B2(new_n819), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n650), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n610), .B1(new_n630), .B2(new_n631), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n609), .A2(new_n611), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n621), .B(new_n625), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n633), .B2(new_n637), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n679), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n597), .B1(new_n826), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(KEYINPUT114), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n837), .B(new_n829), .C1(new_n633), .C2(new_n637), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n822), .A3(new_n823), .ZN(new_n840));
  INV_X1    g639(.A(new_n825), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n598), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n835), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n822), .A2(new_n823), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n597), .A2(new_n825), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT115), .A4(new_n839), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n707), .B1(new_n834), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n739), .A2(new_n679), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n809), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n849), .ZN(new_n851));
  INV_X1    g650(.A(new_n638), .ZN(new_n852));
  INV_X1    g651(.A(new_n649), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n632), .B1(new_n641), .B2(new_n642), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT91), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n636), .A3(new_n643), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n648), .B1(new_n856), .B2(new_n639), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n852), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n844), .A3(new_n841), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n832), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n860), .A2(new_n597), .B1(new_n843), .B2(new_n846), .ZN(new_n861));
  OAI211_X1 g660(.A(KEYINPUT116), .B(new_n851), .C1(new_n861), .C2(new_n707), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n731), .A2(new_n694), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n407), .A2(new_n440), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n850), .A2(new_n862), .A3(new_n863), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n650), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g666(.A1(new_n865), .A2(new_n680), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(G120gat), .Z(G1341gat));
  NOR2_X1   g668(.A1(new_n865), .A2(new_n534), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G127gat), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n870), .A2(G127gat), .ZN(new_n874));
  OAI22_X1  g673(.A1(new_n872), .A2(new_n873), .B1(KEYINPUT117), .B2(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(G1342gat));
  NOR3_X1   g679(.A1(new_n865), .A2(G134gat), .A3(new_n597), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n882));
  OR3_X1    g681(.A1(new_n881), .A2(KEYINPUT119), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n865), .B2(new_n597), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n882), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n886), .ZN(G1343gat));
  INV_X1    g686(.A(new_n371), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n850), .A2(new_n862), .A3(new_n888), .A4(new_n864), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(G141gat), .A3(new_n650), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n864), .A2(new_n368), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n858), .A2(new_n820), .A3(new_n841), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n598), .B1(new_n892), .B2(new_n832), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n707), .B1(new_n894), .B2(new_n847), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n731), .B1(new_n895), .B2(new_n849), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n891), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n850), .A2(new_n862), .A3(new_n898), .A4(new_n731), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n899), .A3(new_n858), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n890), .B1(G141gat), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g700(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n902));
  NAND2_X1  g701(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1344gat));
  INV_X1    g705(.A(new_n889), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n226), .A3(new_n679), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n850), .A2(new_n731), .A3(new_n862), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n891), .A2(new_n680), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT121), .B1(new_n739), .B2(new_n679), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n599), .A2(new_n914), .A3(new_n650), .A4(new_n680), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n840), .A2(new_n842), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n534), .B1(new_n893), .B2(new_n917), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT57), .B(new_n480), .C1(new_n916), .C2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n911), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n226), .B1(new_n921), .B2(KEYINPUT122), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n919), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n912), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n909), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n897), .A2(new_n899), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n909), .B1(new_n927), .B2(new_n680), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n226), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n908), .B1(new_n926), .B2(new_n929), .ZN(G1345gat));
  NOR3_X1   g729(.A1(new_n927), .A2(new_n238), .A3(new_n534), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n889), .A2(new_n534), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n931), .B1(new_n934), .B2(new_n238), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n927), .B2(new_n597), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n907), .A2(new_n239), .A3(new_n598), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1347gat));
  NAND4_X1  g737(.A1(new_n850), .A2(new_n862), .A3(new_n407), .A4(new_n863), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n441), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n858), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n679), .ZN(new_n943));
  XOR2_X1   g742(.A(KEYINPUT124), .B(G176gat), .Z(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(G1349gat));
  NAND2_X1  g744(.A1(new_n940), .A2(new_n707), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n314), .ZN(new_n947));
  NAND2_X1  g746(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n939), .A2(new_n534), .A3(new_n323), .A4(new_n441), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OR2_X1    g749(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G183gat), .B1(new_n940), .B2(new_n707), .ZN(new_n953));
  OAI211_X1 g752(.A(KEYINPUT125), .B(KEYINPUT60), .C1(new_n953), .C2(new_n949), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n952), .A2(new_n954), .ZN(G1350gat));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n598), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(G190gat), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n956), .A2(G190gat), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n959), .B(new_n962), .C1(G190gat), .C2(new_n956), .ZN(G1351gat));
  AOI211_X1 g762(.A(new_n441), .B(new_n919), .C1(new_n910), .C2(KEYINPUT57), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n767), .A2(new_n727), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(new_n858), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G197gat), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n850), .A2(new_n862), .A3(new_n407), .A4(new_n888), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(new_n441), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OR2_X1    g769(.A1(new_n650), .A2(G197gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1352gat));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n964), .A2(new_n973), .A3(new_n679), .A4(new_n965), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n923), .A2(new_n679), .A3(new_n440), .A4(new_n965), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n974), .A2(new_n976), .A3(G204gat), .ZN(new_n977));
  INV_X1    g776(.A(G204gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n978), .A3(new_n679), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(G1353gat));
  OR3_X1    g781(.A1(new_n970), .A2(G211gat), .A3(new_n534), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n923), .A2(new_n707), .A3(new_n440), .A4(new_n965), .ZN(new_n984));
  AND3_X1   g783(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n985));
  AOI21_X1  g784(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n985), .B2(new_n986), .ZN(G1354gat));
  AND4_X1   g786(.A1(G218gat), .A2(new_n964), .A3(new_n598), .A4(new_n965), .ZN(new_n988));
  AOI21_X1  g787(.A(G218gat), .B1(new_n969), .B2(new_n598), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n988), .A2(new_n989), .ZN(G1355gat));
endmodule


