//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(G104), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  AOI21_X1  g004(.A(G107), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n191), .A2(new_n192), .B1(G104), .B2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n191), .A2(new_n192), .ZN(new_n195));
  OAI21_X1  g009(.A(G101), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n187), .A2(KEYINPUT3), .A3(G107), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n191), .B2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n188), .A2(new_n190), .A3(G107), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n206));
  INV_X1    g020(.A(G113), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n208), .A2(new_n209), .B1(new_n206), .B2(new_n207), .ZN(new_n210));
  XNOR2_X1  g024(.A(G116), .B(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G119), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT5), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n207), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n196), .A2(new_n204), .A3(new_n212), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G119), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(G116), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT69), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n210), .B(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n201), .B(new_n198), .C1(new_n191), .C2(new_n199), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT4), .B1(new_n200), .B2(new_n203), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n224), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n224), .B2(new_n229), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n219), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G110), .B(G122), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n219), .B(new_n234), .C1(new_n227), .C2(new_n232), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(KEYINPUT6), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(G143), .B2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n239), .B1(new_n242), .B2(KEYINPUT67), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(KEYINPUT67), .B2(new_n242), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n241), .B2(G143), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT64), .A3(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n241), .A2(G143), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n241), .B2(G143), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n247), .A2(KEYINPUT65), .A3(G146), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n253), .A2(new_n254), .B1(G143), .B2(new_n241), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n244), .A2(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n255), .A2(new_n263), .A3(new_n260), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n262), .A2(new_n264), .B1(new_n251), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n267), .B2(new_n258), .ZN(new_n268));
  INV_X1    g082(.A(G224), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G953), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT82), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n268), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n233), .A2(new_n273), .A3(new_n235), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n238), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT83), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n238), .A2(new_n272), .A3(new_n277), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G902), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n196), .A2(new_n204), .ZN(new_n281));
  XOR2_X1   g095(.A(new_n217), .B(KEYINPUT85), .Z(new_n282));
  XNOR2_X1  g096(.A(new_n213), .B(KEYINPUT84), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n212), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n234), .B(KEYINPUT8), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n212), .A2(new_n218), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(new_n286), .C1(new_n281), .C2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT7), .B1(new_n269), .B2(G953), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n259), .B(new_n290), .C1(new_n258), .C2(new_n267), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n268), .A2(new_n289), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n237), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n280), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n279), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT86), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n295), .B1(new_n276), .B2(new_n278), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G214), .B1(G237), .B2(G902), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n302), .A2(new_n301), .A3(new_n298), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n304), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT87), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n310), .A3(new_n307), .A4(new_n305), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT9), .B(G234), .ZN(new_n313));
  OAI21_X1  g127(.A(G221), .B1(new_n313), .B2(G902), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G469), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(new_n280), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n255), .A2(new_n256), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT80), .ZN(new_n320));
  OAI21_X1  g134(.A(G128), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n320), .B2(new_n319), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(new_n255), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n204), .A3(new_n196), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT10), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n257), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n324), .A2(new_n325), .B1(new_n281), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  INV_X1    g144(.A(G137), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(KEYINPUT11), .A3(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(G131), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI221_X1 g150(.A(new_n267), .B1(new_n225), .B2(new_n226), .C1(new_n230), .C2(new_n231), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n327), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G140), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G227), .ZN(new_n342));
  XOR2_X1   g156(.A(new_n340), .B(new_n342), .Z(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n327), .A2(new_n337), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT81), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n327), .A2(new_n347), .A3(new_n337), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n335), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT67), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n319), .A2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n243), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n251), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n318), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n324), .B1(new_n354), .B2(new_n281), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n355), .A2(KEYINPUT12), .A3(new_n335), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT12), .B1(new_n355), .B2(new_n335), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n338), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n344), .A2(new_n349), .B1(new_n358), .B2(new_n343), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n317), .B1(new_n359), .B2(G469), .ZN(new_n360));
  INV_X1    g174(.A(new_n343), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n349), .B2(new_n338), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(new_n339), .A3(new_n343), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n316), .B(new_n280), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n315), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n367), .A2(G143), .A3(G214), .ZN(new_n368));
  AOI21_X1  g182(.A(G143), .B1(new_n367), .B2(G214), .ZN(new_n369));
  OR2_X1    g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  INV_X1    g186(.A(G131), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT17), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G125), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n258), .A2(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(KEYINPUT16), .B2(new_n378), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n241), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n382), .B(G146), .C1(KEYINPUT16), .C2(new_n378), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n372), .A2(new_n373), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n376), .A2(new_n384), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n187), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n390), .B(KEYINPUT89), .Z(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT18), .A2(G131), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n372), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n381), .B2(new_n241), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n380), .A2(KEYINPUT74), .A3(G146), .ZN(new_n397));
  OAI22_X1  g211(.A1(new_n396), .A2(new_n397), .B1(new_n241), .B2(new_n381), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n381), .A2(KEYINPUT19), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT19), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n241), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n374), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n403), .B(new_n385), .C1(new_n404), .C2(new_n386), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n390), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT88), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n409), .B(new_n390), .C1(new_n399), .C2(new_n405), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n400), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT90), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n414), .B(new_n400), .C1(new_n408), .C2(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n418), .A3(new_n413), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n388), .A2(new_n399), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n407), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n422), .B2(new_n400), .ZN(new_n423));
  INV_X1    g237(.A(G475), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(G128), .A3(new_n247), .ZN(new_n430));
  XNOR2_X1  g244(.A(G128), .B(G143), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n430), .B(G134), .C1(new_n432), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n329), .ZN(new_n434));
  XNOR2_X1  g248(.A(G116), .B(G122), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(new_n193), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n431), .B(new_n329), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n214), .A2(KEYINPUT14), .A3(G122), .ZN(new_n439));
  INV_X1    g253(.A(new_n435), .ZN(new_n440));
  OAI211_X1 g254(.A(G107), .B(new_n439), .C1(new_n440), .C2(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n435), .A2(new_n193), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G217), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n313), .A2(new_n445), .A3(G953), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n444), .B(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n448), .A2(new_n280), .ZN(new_n449));
  INV_X1    g263(.A(G478), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(KEYINPUT15), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(KEYINPUT15), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n449), .A2(KEYINPUT93), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(KEYINPUT93), .A3(new_n280), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n455), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n457), .A2(KEYINPUT94), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT94), .B1(new_n457), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G952), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  INV_X1    g278(.A(G234), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n280), .B(new_n341), .C1(G234), .C2(G237), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT21), .B(G898), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n462), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n366), .A2(new_n428), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n312), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n384), .A2(new_n385), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT23), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n220), .B2(G128), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n480), .B(new_n481), .C1(G119), .C2(new_n239), .ZN(new_n482));
  XNOR2_X1  g296(.A(G119), .B(G128), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT24), .B(G110), .Z(new_n484));
  AOI22_X1  g298(.A1(new_n482), .A2(G110), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  OAI22_X1  g300(.A1(new_n482), .A2(G110), .B1(new_n483), .B2(new_n484), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n385), .B(new_n487), .C1(new_n397), .C2(new_n396), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT75), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT22), .B(G137), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n490), .B(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n486), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n486), .B2(new_n488), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n280), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT76), .A2(KEYINPUT25), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n495), .B2(new_n496), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n445), .B1(G234), .B2(new_n280), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(G902), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n493), .B2(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT73), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n334), .A2(G131), .ZN(new_n512));
  INV_X1    g326(.A(new_n333), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n329), .A2(G137), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n511), .B1(new_n257), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n354), .A2(new_n518), .A3(KEYINPUT70), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n223), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n262), .A2(new_n264), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n251), .A2(new_n266), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n335), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT72), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT26), .B(G101), .Z(new_n527));
  NAND2_X1  g341(.A1(new_n367), .A2(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n354), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n524), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT30), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n520), .A2(new_n524), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(KEYINPUT30), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n538), .B2(new_n521), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n517), .A2(new_n519), .B1(new_n335), .B2(new_n267), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n531), .B1(new_n540), .B2(new_n521), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n541), .A2(new_n526), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n510), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n534), .A2(new_n524), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n545), .B2(new_n540), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n547), .A2(new_n223), .B1(new_n541), .B2(new_n526), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n525), .A2(new_n532), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(KEYINPUT31), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n543), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT28), .B1(new_n544), .B2(new_n521), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n535), .A2(new_n223), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n525), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n531), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n509), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n507), .B1(new_n559), .B2(KEYINPUT32), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n543), .A2(new_n551), .B1(new_n531), .B2(new_n557), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT32), .ZN(new_n562));
  NOR4_X1   g376(.A1(new_n561), .A2(KEYINPUT73), .A3(new_n562), .A4(new_n509), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n540), .A2(new_n545), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n223), .B1(new_n565), .B2(new_n536), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n566), .A2(new_n525), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n532), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT29), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n557), .B2(new_n531), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n537), .A2(new_n223), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n572), .A2(new_n525), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n554), .B1(new_n573), .B2(new_n556), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n532), .A2(KEYINPUT29), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n280), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G472), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n562), .B1(new_n561), .B2(new_n509), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n506), .B1(new_n564), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n312), .A2(KEYINPUT95), .A3(new_n474), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n477), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(G101), .ZN(G3));
  OAI21_X1  g398(.A(G472), .B1(new_n561), .B2(G902), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n561), .B2(new_n509), .ZN(new_n586));
  INV_X1    g400(.A(new_n506), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n366), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n298), .B1(new_n279), .B2(new_n296), .ZN(new_n591));
  AOI211_X1 g405(.A(new_n299), .B(new_n295), .C1(new_n276), .C2(new_n278), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n305), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n447), .A2(KEYINPUT97), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n444), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n444), .B2(new_n596), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n448), .A2(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(G478), .A3(new_n280), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(G478), .B2(new_n449), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n427), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n471), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n594), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n590), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT34), .B(G104), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NAND4_X1  g422(.A1(new_n412), .A2(new_n418), .A3(new_n413), .A4(new_n415), .ZN(new_n609));
  OR2_X1    g423(.A1(new_n425), .A2(KEYINPUT98), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n425), .A2(KEYINPUT98), .ZN(new_n611));
  AOI22_X1  g425(.A1(new_n417), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n594), .A2(new_n462), .A3(new_n604), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n590), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT99), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G107), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n486), .A2(new_n488), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n492), .A2(KEYINPUT36), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n504), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n503), .A2(new_n618), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n502), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n497), .B2(new_n500), .ZN(new_n625));
  INV_X1    g439(.A(new_n622), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n586), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n477), .A2(new_n582), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT37), .B(G110), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT101), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(G12));
  INV_X1    g447(.A(new_n366), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n634), .A2(new_n628), .A3(new_n593), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n417), .A2(new_n609), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n610), .A2(new_n611), .ZN(new_n637));
  INV_X1    g451(.A(new_n469), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT102), .B(G900), .Z(new_n639));
  OAI21_X1  g453(.A(new_n467), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n636), .A2(new_n462), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n612), .A2(new_n643), .A3(new_n462), .A4(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT31), .B1(new_n548), .B2(new_n550), .ZN(new_n647));
  AND4_X1   g461(.A1(KEYINPUT31), .A2(new_n566), .A3(new_n550), .A4(new_n533), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n558), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(KEYINPUT32), .A3(new_n508), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT73), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n559), .A2(new_n507), .A3(KEYINPUT32), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(new_n652), .A3(new_n578), .A4(new_n577), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n635), .A2(new_n646), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NAND2_X1  g469(.A1(new_n548), .A2(new_n550), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n573), .A2(new_n532), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n280), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G472), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n651), .A2(new_n652), .A3(new_n578), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n591), .A2(new_n592), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n306), .B1(new_n664), .B2(new_n301), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n458), .B(new_n456), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT94), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n457), .A2(new_n459), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT94), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n426), .B2(new_n420), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n623), .A2(new_n627), .ZN(new_n674));
  INV_X1    g488(.A(new_n305), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n640), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n366), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n673), .B(new_n676), .C1(new_n678), .C2(KEYINPUT40), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n679), .B1(KEYINPUT40), .B2(new_n678), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n663), .A2(new_n666), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT105), .B(G143), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G45));
  NAND3_X1  g497(.A1(new_n427), .A2(new_n602), .A3(new_n640), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n635), .A2(new_n653), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NOR2_X1   g501(.A1(new_n362), .A2(new_n364), .ZN(new_n688));
  OAI21_X1  g502(.A(G469), .B1(new_n688), .B2(G902), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n314), .A3(new_n365), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(KEYINPUT106), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n691), .A2(new_n653), .A3(new_n587), .A4(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n605), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n693), .A2(new_n613), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n214), .ZN(G18));
  NOR2_X1   g512(.A1(new_n690), .A2(new_n593), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n428), .A2(new_n674), .A3(new_n472), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n653), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n574), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n556), .B1(new_n572), .B2(new_n525), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n705), .B2(new_n553), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n531), .ZN(new_n707));
  OAI22_X1  g521(.A1(new_n704), .A2(new_n707), .B1(new_n647), .B2(new_n648), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n508), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n585), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n710), .A2(new_n506), .A3(new_n471), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n673), .B(new_n305), .C1(new_n591), .C2(new_n592), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n691), .A3(new_n692), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NOR3_X1   g529(.A1(new_n710), .A2(new_n628), .A3(new_n684), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n699), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  NOR2_X1   g532(.A1(new_n665), .A2(new_n675), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n366), .ZN(new_n720));
  INV_X1    g534(.A(new_n650), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n685), .B(new_n587), .C1(new_n579), .C2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT42), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n581), .A2(new_n366), .A3(new_n719), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n373), .ZN(G33));
  NAND4_X1  g541(.A1(new_n581), .A2(new_n366), .A3(new_n646), .A4(new_n719), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  NAND2_X1  g543(.A1(new_n428), .A2(new_n602), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n586), .A3(new_n674), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  INV_X1    g550(.A(new_n719), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n359), .A2(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n359), .A2(KEYINPUT45), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(G469), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n317), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(KEYINPUT46), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n365), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n744), .B1(KEYINPUT108), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n747), .B1(KEYINPUT108), .B2(new_n746), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n748), .A2(new_n314), .A3(new_n677), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n738), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  NOR3_X1   g565(.A1(new_n579), .A2(new_n560), .A3(new_n563), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n719), .A3(new_n506), .A4(new_n685), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT109), .Z(new_n754));
  AND3_X1   g568(.A1(new_n748), .A2(KEYINPUT47), .A3(new_n314), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT47), .B1(new_n748), .B2(new_n314), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n732), .A2(new_n468), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n732), .A2(KEYINPUT114), .A3(new_n468), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n690), .B(new_n737), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n585), .A3(new_n674), .A4(new_n709), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n737), .A2(new_n690), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n662), .A2(new_n587), .A3(new_n468), .A4(new_n766), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n767), .A2(new_n427), .A3(new_n602), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n710), .A2(new_n506), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n762), .B2(new_n763), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n666), .A2(new_n305), .A3(new_n690), .ZN(new_n772));
  AND3_X1   g586(.A1(new_n771), .A2(KEYINPUT50), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT50), .B1(new_n771), .B2(new_n772), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n765), .B(new_n768), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n719), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n755), .A2(new_n756), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n689), .A2(new_n315), .A3(new_n365), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n759), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n771), .A2(new_n699), .ZN(new_n781));
  INV_X1    g595(.A(new_n603), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n781), .B(new_n464), .C1(new_n782), .C2(new_n767), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n506), .B1(new_n580), .B2(new_n650), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n764), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(KEYINPUT48), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(KEYINPUT48), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n775), .A2(new_n779), .A3(new_n759), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n645), .B1(new_n564), .B2(new_n580), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n792), .A2(new_n635), .B1(new_n699), .B2(new_n716), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n503), .A2(new_n622), .A3(new_n640), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n634), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n713), .A2(new_n661), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(KEYINPUT52), .A3(new_n686), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n654), .A2(new_n686), .A3(new_n717), .A4(new_n796), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n674), .A2(new_n667), .A3(new_n612), .A4(new_n640), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n564), .B2(new_n580), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n366), .B(new_n719), .C1(new_n803), .C2(new_n716), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n723), .A2(new_n804), .A3(new_n725), .A4(new_n728), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n714), .B(new_n701), .C1(new_n693), .C2(new_n605), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n697), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n312), .A2(new_n604), .A3(new_n589), .A4(new_n603), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n427), .A2(new_n667), .A3(new_n471), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n310), .B1(new_n665), .B2(new_n305), .ZN(new_n812));
  INV_X1    g626(.A(new_n311), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT112), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n312), .A2(new_n816), .A3(new_n811), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n589), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n583), .A2(new_n630), .A3(new_n810), .A4(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT95), .B1(new_n312), .B2(new_n474), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n476), .B(new_n473), .C1(new_n309), .C2(new_n311), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n590), .B1(new_n814), .B2(KEYINPUT112), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n824), .A2(new_n629), .B1(new_n825), .B2(new_n817), .ZN(new_n826));
  INV_X1    g640(.A(new_n810), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n824), .B2(new_n581), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n821), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n809), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n793), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n833), .B2(KEYINPUT52), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT54), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n819), .A2(KEYINPUT113), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n826), .A2(new_n828), .A3(new_n821), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n808), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n832), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n791), .A2(new_n836), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT115), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n791), .A2(new_n836), .A3(new_n848), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n463), .A2(new_n341), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n506), .A2(new_n675), .A3(new_n315), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT110), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n689), .A2(new_n365), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(KEYINPUT49), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n853), .A2(new_n730), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(KEYINPUT49), .B2(new_n854), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n663), .A3(new_n666), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT111), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n851), .A2(new_n859), .ZN(G75));
  NOR2_X1   g674(.A1(new_n341), .A2(G952), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n832), .A2(new_n844), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(G210), .A3(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n238), .A2(new_n274), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(new_n272), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT55), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n862), .B1(new_n866), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n863), .A2(new_n872), .A3(G210), .A4(G902), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n869), .A2(new_n865), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n871), .A2(KEYINPUT117), .A3(new_n873), .A4(new_n874), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(G51));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n741), .B(KEYINPUT120), .Z(new_n881));
  AOI211_X1 g695(.A(new_n280), .B(new_n881), .C1(new_n832), .C2(new_n844), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n317), .B(KEYINPUT118), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT57), .Z(new_n884));
  NOR2_X1   g698(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n842), .B(new_n808), .C1(new_n838), .C2(new_n839), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n837), .B1(new_n832), .B2(new_n844), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n688), .B(KEYINPUT119), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n882), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n880), .B1(new_n891), .B2(new_n861), .ZN(new_n892));
  INV_X1    g706(.A(new_n890), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT54), .B1(new_n885), .B2(new_n886), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n845), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n893), .B1(new_n895), .B2(new_n884), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT121), .B(new_n862), .C1(new_n896), .C2(new_n882), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n892), .A2(new_n897), .ZN(G54));
  NAND2_X1  g712(.A1(new_n412), .A2(new_n415), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n863), .A2(G902), .ZN(new_n900));
  AND3_X1   g714(.A1(KEYINPUT122), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(KEYINPUT58), .B2(G475), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n899), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n862), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n900), .A2(new_n899), .A3(new_n903), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G60));
  NAND2_X1  g721(.A1(new_n836), .A2(new_n845), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n600), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n895), .A2(new_n600), .A3(new_n910), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n861), .A3(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n863), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n493), .A2(new_n494), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n863), .A2(new_n621), .A3(new_n915), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n862), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G66));
  OAI21_X1  g736(.A(G953), .B1(new_n470), .B2(new_n269), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n697), .B(new_n806), .C1(new_n838), .C2(new_n839), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n867), .B1(G898), .B2(new_n341), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  NOR2_X1   g741(.A1(new_n401), .A2(new_n402), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n547), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n793), .A2(new_n686), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n681), .A2(KEYINPUT62), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n603), .B1(new_n428), .B2(new_n669), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n678), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n737), .A2(new_n752), .A3(new_n506), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n931), .A2(new_n750), .A3(new_n757), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n681), .B2(new_n930), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n929), .B1(new_n941), .B2(G953), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n929), .B1(G900), .B2(G953), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n784), .A2(new_n713), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n749), .B1(new_n738), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n728), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n930), .A2(new_n726), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n757), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n948), .B2(G953), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n942), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n341), .B1(G227), .B2(G900), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n949), .B2(KEYINPUT125), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n950), .B(new_n952), .Z(G72));
  XNOR2_X1  g767(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n835), .B(new_n957), .C1(new_n657), .C2(new_n568), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT127), .ZN(new_n959));
  AND4_X1   g773(.A1(new_n757), .A2(new_n924), .A3(new_n947), .A4(new_n945), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n531), .B(new_n567), .C1(new_n960), .C2(new_n956), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n941), .B2(new_n924), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n567), .A2(new_n531), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n961), .B(new_n862), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n959), .A2(new_n964), .ZN(G57));
endmodule


