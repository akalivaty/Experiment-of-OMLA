//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n206), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n209), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT0), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n219), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n222), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G50), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n252), .A2(new_n254), .B1(G50), .B2(new_n251), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n223), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n256), .B1(new_n257), .B2(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(new_n211), .C2(new_n268), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G1), .A3(G13), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT65), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G226), .ZN(new_n282));
  INV_X1    g0082(.A(new_n277), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(new_n274), .A3(G274), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n276), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT66), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G169), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  AOI211_X1 g0088(.A(new_n263), .B(new_n287), .C1(new_n288), .C2(new_n286), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n263), .B1(KEYINPUT71), .B2(KEYINPUT9), .ZN(new_n290));
  OR2_X1    g0090(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n293));
  INV_X1    g0093(.A(new_n286), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(KEYINPUT10), .B1(new_n294), .B2(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(KEYINPUT72), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n293), .A2(new_n297), .A3(new_n298), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n292), .B1(new_n301), .B2(new_n286), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT10), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n289), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  OAI211_X1 g0107(.A(G232), .B(new_n269), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G107), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n275), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n274), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n313));
  OAI21_X1  g0113(.A(G244), .B1(new_n313), .B2(new_n278), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n312), .A2(G190), .A3(new_n284), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT67), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n314), .A2(new_n284), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n318), .A2(KEYINPUT67), .A3(G190), .A4(new_n312), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G13), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n321), .A2(G1), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n322), .A2(new_n323), .A3(G20), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n251), .A2(KEYINPUT68), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n248), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(G77), .A3(new_n253), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n260), .A2(new_n259), .B1(new_n223), .B2(new_n211), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(new_n261), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n248), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n251), .B(new_n323), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT69), .B1(new_n332), .B2(new_n211), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n324), .A2(new_n325), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT69), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n334), .A2(new_n335), .A3(G77), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n327), .B(new_n331), .C1(new_n333), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n318), .A2(new_n312), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n320), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n318), .A2(new_n288), .A3(new_n312), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n337), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT70), .ZN(new_n346));
  OAI211_X1 g0146(.A(G232), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(new_n269), .C1(new_n306), .C2(new_n307), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n275), .ZN(new_n351));
  OAI21_X1  g0151(.A(G238), .B1(new_n313), .B2(new_n278), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n352), .A3(new_n284), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT13), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n351), .A2(new_n352), .A3(new_n355), .A4(new_n284), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(G190), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n326), .A2(G68), .A3(new_n253), .ZN(new_n358));
  INV_X1    g0158(.A(G68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G20), .ZN(new_n360));
  OAI221_X1 g0160(.A(new_n360), .B1(new_n261), .B2(new_n211), .C1(new_n259), .C2(new_n202), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  AND3_X1   g0162(.A1(new_n361), .A2(new_n362), .A3(new_n248), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n361), .B2(new_n248), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n322), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n366), .A2(new_n360), .A3(KEYINPUT12), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n332), .A2(new_n359), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(KEYINPUT12), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n357), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n301), .B1(new_n354), .B2(new_n356), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT73), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n354), .A2(new_n356), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G200), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n370), .A4(new_n357), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n346), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  INV_X1    g0179(.A(G58), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(new_n359), .ZN(new_n381));
  OAI21_X1  g0181(.A(G20), .B1(new_n381), .B2(new_n201), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n258), .A2(G159), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT74), .B(G33), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n223), .B(new_n266), .C1(new_n386), .C2(new_n264), .ZN(new_n387));
  OAI21_X1  g0187(.A(G68), .B1(new_n387), .B2(KEYINPUT7), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n265), .A2(KEYINPUT74), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT74), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G33), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n307), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n389), .B1(new_n394), .B2(new_n223), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT16), .B(new_n385), .C1(new_n388), .C2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n267), .A2(new_n223), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(new_n389), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(KEYINPUT3), .B2(new_n393), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n389), .B1(new_n398), .B2(new_n307), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n359), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(new_n384), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(new_n403), .A3(new_n248), .ZN(new_n404));
  INV_X1    g0204(.A(new_n260), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n253), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n406), .A2(new_n252), .B1(new_n251), .B2(new_n405), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT75), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n274), .A2(new_n277), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n284), .B1(new_n232), .B2(new_n410), .ZN(new_n411));
  MUX2_X1   g0211(.A(G223), .B(G226), .S(G1698), .Z(new_n412));
  AOI21_X1  g0212(.A(new_n264), .B1(new_n390), .B2(new_n392), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n307), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n411), .B1(new_n416), .B2(new_n275), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G179), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n341), .B2(new_n417), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n379), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n404), .A2(new_n408), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n274), .B1(new_n414), .B2(new_n415), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT76), .B(G190), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n423), .A2(KEYINPUT77), .A3(new_n411), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n411), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n266), .B1(new_n386), .B2(new_n264), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(new_n412), .B1(G33), .B2(G87), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n274), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT77), .B1(new_n430), .B2(new_n301), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n424), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n422), .A2(new_n433), .A3(KEYINPUT17), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n301), .B1(new_n423), .B2(new_n411), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT77), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n424), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n417), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n425), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n435), .B1(new_n441), .B2(new_n409), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n409), .A2(new_n379), .A3(new_n419), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n421), .A2(new_n434), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n370), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n374), .A2(new_n447), .A3(G169), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n354), .A2(G179), .A3(new_n356), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n447), .B1(new_n374), .B2(G169), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n446), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n304), .A2(new_n378), .A3(new_n445), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT80), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G238), .A2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n212), .B2(G1698), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n413), .B2(new_n307), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n458), .B1(new_n390), .B2(new_n392), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n274), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n250), .A2(G45), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(G250), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n274), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n274), .A2(G274), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n465), .B2(new_n462), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n454), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n465), .ZN(new_n468));
  INV_X1    g0268(.A(new_n462), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n468), .A2(new_n469), .B1(new_n274), .B2(new_n463), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n459), .B1(new_n428), .B2(new_n456), .ZN(new_n471));
  OAI211_X1 g0271(.A(KEYINPUT80), .B(new_n470), .C1(new_n471), .C2(new_n274), .ZN(new_n472));
  AOI21_X1  g0272(.A(G169), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n288), .A3(new_n472), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n249), .B(new_n251), .C1(G1), .C2(new_n265), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n329), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n334), .A2(new_n477), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n428), .A2(new_n223), .A3(G68), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT19), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n223), .B1(new_n349), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(new_n205), .A3(new_n206), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n261), .B2(new_n205), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n478), .B(new_n480), .C1(new_n489), .C2(new_n249), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n474), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n467), .A2(G190), .A3(new_n472), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n249), .B1(new_n481), .B2(new_n488), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n475), .A2(new_n484), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(new_n479), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n301), .B1(new_n467), .B2(new_n472), .ZN(new_n497));
  OAI22_X1  g0297(.A1(new_n473), .A2(new_n491), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n212), .A2(G1698), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G238), .B2(G1698), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n391), .A2(G33), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n265), .A2(KEYINPUT74), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT3), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(new_n266), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n275), .B1(new_n506), .B2(new_n459), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT80), .B1(new_n507), .B2(new_n470), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n461), .A2(new_n454), .A3(new_n466), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n341), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(new_n474), .A3(new_n490), .ZN(new_n511));
  OAI21_X1  g0311(.A(G200), .B1(new_n508), .B2(new_n509), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(new_n492), .A3(new_n495), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT81), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n500), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n458), .B1(new_n250), .B2(G33), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n334), .A2(new_n249), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n516), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT83), .B1(new_n334), .B2(G116), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT83), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n332), .A2(new_n522), .A3(new_n458), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G283), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(new_n223), .C1(G33), .C2(new_n205), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n458), .A2(G20), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n248), .A2(KEYINPUT84), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT84), .B1(new_n248), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT20), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT5), .B(G41), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n469), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n537), .A2(G270), .A3(new_n274), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n213), .A2(G1698), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(G257), .B2(G1698), .ZN(new_n540));
  INV_X1    g0340(.A(G303), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n394), .A2(new_n540), .B1(new_n541), .B2(new_n268), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n542), .B2(new_n275), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n536), .A2(new_n469), .A3(G274), .A4(new_n274), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n341), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n535), .A2(new_n545), .A3(KEYINPUT21), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n505), .B2(new_n266), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n268), .A2(new_n541), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n275), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n538), .ZN(new_n550));
  AND4_X1   g0350(.A1(G179), .A2(new_n549), .A3(new_n544), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n535), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT21), .B1(new_n535), .B2(new_n545), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(new_n424), .A3(new_n550), .A4(new_n544), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n524), .A3(new_n534), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n301), .B1(new_n543), .B2(new_n544), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g0358(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  MUX2_X1   g0359(.A(G250), .B(G257), .S(G1698), .Z(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n413), .B2(new_n307), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n393), .A2(G294), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n274), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n537), .A2(G264), .A3(new_n274), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n544), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n566), .A2(new_n341), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n563), .A2(new_n565), .A3(new_n288), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT85), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n223), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n459), .A2(new_n223), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n223), .A2(G87), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n309), .B2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n576), .A2(new_n484), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n428), .A2(new_n223), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n571), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n581), .A2(new_n571), .A3(new_n578), .A4(new_n575), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT24), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n578), .A3(new_n575), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT85), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT24), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n249), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n251), .A2(G107), .ZN(new_n591));
  XOR2_X1   g0391(.A(new_n591), .B(KEYINPUT25), .Z(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(G107), .B2(new_n476), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n570), .B1(new_n590), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n587), .A2(new_n588), .A3(new_n583), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n588), .B1(new_n587), .B2(new_n583), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n248), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n566), .A2(new_n301), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(G190), .B2(new_n566), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n212), .A2(G1698), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n602), .B1(new_n394), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n602), .A2(new_n212), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n606), .B(new_n269), .C1(new_n307), .C2(new_n306), .ZN(new_n607));
  OAI211_X1 g0407(.A(G250), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(new_n525), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n274), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n275), .B1(new_n469), .B2(new_n536), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G257), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n544), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT79), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT4), .B1(new_n428), .B2(new_n603), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n525), .A3(new_n608), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n275), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT79), .ZN(new_n618));
  INV_X1    g0418(.A(new_n544), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n611), .B2(G257), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n341), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n610), .A2(new_n613), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n258), .A2(G77), .ZN(new_n625));
  XNOR2_X1  g0425(.A(new_n625), .B(KEYINPUT78), .ZN(new_n626));
  NAND2_X1  g0426(.A1(G97), .A2(G107), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT6), .B1(new_n207), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n626), .B1(new_n223), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n206), .B1(new_n400), .B2(new_n401), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n248), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n251), .A2(G97), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n476), .B2(G97), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n624), .A2(new_n288), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n614), .A2(G190), .A3(new_n621), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n635), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n301), .B1(new_n617), .B2(new_n620), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n623), .A2(new_n636), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n559), .A2(new_n595), .A3(new_n601), .A4(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n453), .A2(new_n515), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n443), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(new_n420), .ZN(new_n645));
  INV_X1    g0445(.A(new_n452), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n375), .A2(new_n370), .A3(new_n357), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n342), .A2(new_n337), .A3(new_n343), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n434), .A2(new_n442), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n300), .A2(new_n303), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n289), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n507), .A2(new_n470), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n341), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n474), .A2(new_n656), .A3(new_n490), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(G200), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n492), .A2(new_n495), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n641), .A2(new_n601), .A3(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n553), .A2(new_n554), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n595), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n657), .A2(new_n665), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n623), .A2(new_n657), .A3(new_n659), .A4(new_n636), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(KEYINPUT26), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n623), .A2(new_n636), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n500), .A2(new_n514), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n669), .B1(new_n672), .B2(KEYINPUT26), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT87), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n664), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI211_X1 g0475(.A(KEYINPUT87), .B(new_n669), .C1(KEYINPUT26), .C2(new_n672), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n654), .B1(new_n677), .B2(new_n453), .ZN(G369));
  OR3_X1    g0478(.A1(new_n366), .A2(KEYINPUT27), .A3(G20), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT27), .B1(new_n366), .B2(G20), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n535), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n662), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n559), .A2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n683), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT88), .B1(new_n595), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n569), .B1(new_n598), .B2(new_n593), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT88), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(new_n683), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n683), .B1(new_n590), .B2(new_n594), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(new_n595), .A3(new_n601), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n689), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n595), .A2(new_n683), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n662), .A2(new_n683), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n226), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n485), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n221), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n511), .A2(new_n513), .A3(KEYINPUT81), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT81), .B1(new_n511), .B2(new_n513), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n713), .A3(new_n670), .ZN(new_n714));
  OAI21_X1  g0514(.A(KEYINPUT90), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n671), .A2(KEYINPUT26), .A3(new_n660), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT90), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT26), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n672), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n667), .A2(new_n666), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n661), .B2(new_n663), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n683), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n690), .B1(new_n675), .B2(new_n676), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n725), .A2(KEYINPUT89), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT89), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n568), .A2(new_n467), .A3(new_n472), .A4(new_n543), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n730), .B1(new_n622), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n624), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n543), .A2(new_n544), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n566), .A2(G179), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n733), .A2(new_n655), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n622), .A2(new_n731), .A3(new_n730), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n683), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR3_X1    g0541(.A1(new_n622), .A2(new_n731), .A3(new_n730), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(new_n736), .A3(new_n732), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT31), .B1(new_n743), .B2(new_n683), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n595), .A2(new_n641), .A3(new_n601), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n712), .A2(new_n713), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n746), .A2(new_n747), .A3(new_n559), .A4(new_n690), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G330), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n729), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n711), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n321), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n250), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n705), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n687), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n341), .A2(KEYINPUT93), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n223), .B1(KEYINPUT93), .B2(new_n341), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n222), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n765), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n245), .A2(G45), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT92), .Z(new_n774));
  NOR2_X1   g0574(.A1(new_n428), .A2(new_n704), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(G45), .C2(new_n709), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n268), .A2(new_n226), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT91), .Z(new_n778));
  AOI22_X1  g0578(.A1(new_n778), .A2(G355), .B1(new_n458), .B2(new_n704), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n772), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(G20), .A2(G179), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n301), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G190), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n783), .A2(new_n439), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n223), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n309), .B1(new_n792), .B2(new_n541), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n789), .A2(new_n790), .B1(new_n793), .B2(KEYINPUT99), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n782), .A2(new_n295), .A3(G200), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n787), .B(new_n794), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(new_n295), .A3(new_n301), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G329), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n791), .A2(new_n295), .A3(G200), .ZN(new_n803));
  INV_X1    g0603(.A(G294), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n805), .A2(new_n223), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n801), .B1(new_n802), .B2(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(KEYINPUT99), .B2(new_n793), .ZN(new_n808));
  INV_X1    g0608(.A(G326), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n782), .A2(G200), .A3(new_n424), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n798), .B(new_n808), .C1(new_n809), .C2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n806), .B(KEYINPUT97), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n205), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G68), .B2(new_n796), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT98), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n800), .A2(G159), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT32), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n785), .A2(new_n211), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(G58), .C2(new_n788), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n803), .A2(new_n206), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n792), .A2(new_n484), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n825), .A2(new_n826), .A3(new_n309), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n824), .B(new_n828), .C1(new_n202), .C2(new_n814), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n815), .B1(new_n820), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n780), .B1(new_n830), .B2(new_n770), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n761), .B1(new_n766), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n762), .A2(new_n751), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n760), .B1(new_n833), .B2(new_n688), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT100), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  INV_X1    g0637(.A(new_n770), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G159), .A2(new_n784), .B1(new_n796), .B2(G150), .ZN(new_n839));
  INV_X1    g0639(.A(G143), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n789), .C1(new_n814), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n806), .A2(new_n380), .B1(new_n803), .B2(new_n359), .ZN(new_n844));
  INV_X1    g0644(.A(G132), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n428), .B1(new_n845), .B2(new_n799), .ZN(new_n846));
  INV_X1    g0646(.A(new_n792), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n844), .B(new_n846), .C1(G50), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n309), .B1(new_n799), .B2(new_n786), .C1(new_n484), .C2(new_n803), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n850), .B(new_n818), .C1(G107), .C2(new_n847), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n789), .A2(new_n804), .B1(new_n802), .B2(new_n795), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G116), .B2(new_n784), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(new_n541), .C2(new_n814), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n838), .B1(new_n849), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n770), .A2(new_n763), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n761), .B(new_n855), .C1(new_n211), .C2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n337), .A2(KEYINPUT101), .A3(new_n683), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT101), .B1(new_n337), .B2(new_n683), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n648), .B1(new_n861), .B2(new_n340), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n344), .A2(new_n683), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT102), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n320), .A2(new_n339), .ZN(new_n865));
  INV_X1    g0665(.A(new_n860), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n858), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n344), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  INV_X1    g0669(.A(new_n863), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n857), .B1(new_n764), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n872), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n725), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n690), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n675), .B2(new_n676), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n760), .B1(new_n879), .B2(new_n753), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n879), .A2(new_n753), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(G384));
  INV_X1    g0683(.A(new_n630), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n224), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT36), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n709), .A2(new_n211), .A3(new_n381), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT103), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(G50), .B2(new_n359), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n889), .A2(KEYINPUT103), .ZN(new_n892));
  OAI211_X1 g0692(.A(G1), .B(new_n321), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT104), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n453), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n727), .B2(new_n728), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n654), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n396), .A2(new_n248), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n394), .A2(new_n389), .A3(new_n223), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n387), .A2(KEYINPUT7), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n902), .A3(G68), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT16), .B1(new_n903), .B2(new_n385), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n408), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n681), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n422), .A2(new_n433), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n419), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n436), .A2(new_n437), .B1(new_n417), .B2(new_n439), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n404), .B(new_n408), .C1(new_n910), .C2(new_n425), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n409), .A2(new_n419), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n409), .A2(new_n906), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .A4(new_n899), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT105), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n905), .A2(new_n906), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n908), .A2(new_n917), .A3(new_n911), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT105), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n914), .ZN(new_n921));
  INV_X1    g0721(.A(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n444), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT38), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n921), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n446), .A2(new_n683), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n373), .A2(new_n377), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n450), .A2(new_n451), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n647), .A2(new_n929), .ZN(new_n933));
  INV_X1    g0733(.A(new_n451), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n449), .A3(new_n448), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n446), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n661), .A2(new_n663), .ZN(new_n939));
  INV_X1    g0739(.A(new_n669), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n714), .B2(new_n718), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n939), .B1(new_n941), .B2(KEYINPUT87), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n673), .A2(new_n674), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n876), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n928), .B(new_n938), .C1(new_n944), .C2(new_n863), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n899), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n913), .B1(new_n650), .B2(new_n645), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n925), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n927), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT39), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n927), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n646), .A2(new_n690), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n645), .A2(new_n906), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n945), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n898), .B(new_n959), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n862), .A2(KEYINPUT102), .A3(new_n863), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n869), .B1(new_n868), .B2(new_n870), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n932), .B2(new_n936), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n748), .B2(new_n745), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n919), .A2(new_n914), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n965), .A2(KEYINPUT105), .B1(new_n444), .B2(new_n922), .ZN(new_n966));
  AOI21_X1  g0766(.A(KEYINPUT38), .B1(new_n966), .B2(new_n921), .ZN(new_n967));
  INV_X1    g0767(.A(new_n927), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT40), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n453), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n964), .A2(new_n950), .A3(KEYINPUT40), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n971), .A2(new_n972), .A3(new_n749), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(KEYINPUT40), .B1(new_n928), .B2(new_n964), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n927), .A2(new_n949), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n930), .A2(new_n931), .ZN(new_n977));
  INV_X1    g0777(.A(new_n929), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n452), .A2(new_n647), .A3(new_n929), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n979), .A2(new_n980), .B1(new_n864), .B2(new_n871), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n642), .A2(new_n515), .A3(new_n683), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n739), .A2(new_n740), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n981), .B(KEYINPUT40), .C1(new_n982), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n975), .A2(new_n987), .B1(new_n453), .B2(new_n750), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n974), .A2(new_n988), .A3(G330), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n960), .A2(KEYINPUT106), .A3(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n250), .B2(new_n757), .C1(new_n960), .C2(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT106), .B1(new_n960), .B2(new_n989), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n895), .B1(new_n991), .B2(new_n992), .ZN(G367));
  NOR2_X1   g0793(.A1(new_n495), .A2(new_n690), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n721), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n660), .B1(new_n495), .B2(new_n690), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n640), .A2(new_n637), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n692), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n683), .B1(new_n1003), .B2(new_n670), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n638), .A2(new_n683), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n641), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n670), .B2(new_n690), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n698), .A2(new_n701), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1004), .B1(new_n1008), .B2(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1008), .A2(KEYINPUT42), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1000), .B(new_n1001), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1014), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1011), .B1(new_n1009), .B2(KEYINPUT107), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1016), .A2(new_n1017), .A3(new_n999), .A4(new_n998), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1007), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n699), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1015), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n705), .B(KEYINPUT41), .Z(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n698), .A2(new_n701), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n701), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n695), .B2(new_n697), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n688), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT108), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1007), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1030), .B2(new_n700), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1036), .B1(new_n1034), .B2(new_n1035), .C1(new_n1030), .C2(new_n700), .ZN(new_n1040));
  AOI21_X1  g0840(.A(KEYINPUT45), .B1(new_n702), .B2(new_n1007), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT45), .ZN(new_n1042));
  NOR4_X1   g0842(.A1(new_n1030), .A2(new_n1042), .A3(new_n700), .A4(new_n1020), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1039), .B(new_n1040), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n699), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n699), .A3(KEYINPUT109), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1033), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1027), .B1(new_n1049), .B2(new_n754), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1025), .B1(new_n1050), .B2(new_n758), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n775), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1052), .A2(new_n238), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n771), .B1(new_n226), .B2(new_n329), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n760), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n309), .B1(new_n800), .B2(G137), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n380), .B2(new_n792), .C1(new_n211), .C2(new_n803), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n816), .A2(G68), .ZN(new_n1058));
  INV_X1    g0858(.A(G159), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n795), .C1(new_n257), .C2(new_n789), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(G50), .C2(new_n784), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n840), .B2(new_n814), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n785), .A2(new_n802), .B1(new_n804), .B2(new_n795), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G303), .B2(new_n788), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n792), .A2(new_n458), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT46), .ZN(new_n1066));
  INV_X1    g0866(.A(G317), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n394), .B1(new_n1067), .B2(new_n799), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n803), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(G97), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n206), .B2(new_n806), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1066), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1064), .B(new_n1072), .C1(new_n786), .C2(new_n814), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1062), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT47), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1055), .B1(new_n1075), .B2(new_n770), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n765), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n997), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1051), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(G387));
  NAND3_X1  g0881(.A1(new_n695), .A2(new_n697), .A3(new_n765), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n778), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n1083), .A2(new_n707), .B1(G107), .B2(new_n226), .ZN(new_n1084));
  INV_X1    g0884(.A(G45), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n235), .A2(new_n1085), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n707), .B(new_n1085), .C1(new_n359), .C2(new_n211), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1088));
  NOR3_X1   g0888(.A1(new_n1088), .A2(G50), .A3(new_n260), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(G50), .B2(new_n260), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1052), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1084), .B1(new_n1086), .B2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n760), .B1(new_n1093), .B2(new_n772), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n792), .A2(new_n211), .B1(new_n799), .B2(new_n257), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n784), .A2(G68), .B1(new_n1095), .B2(KEYINPUT111), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT111), .B2(new_n1095), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n789), .A2(new_n202), .B1(new_n260), .B2(new_n795), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n817), .A2(new_n329), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1070), .A2(new_n428), .ZN(new_n1100));
  NOR4_X1   g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n814), .ZN(new_n1102));
  AOI21_X1  g0902(.A(KEYINPUT112), .B1(new_n1102), .B2(G159), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1102), .A2(KEYINPUT112), .A3(G159), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n806), .A2(new_n802), .B1(new_n792), .B2(new_n804), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G317), .A2(new_n788), .B1(new_n796), .B2(G311), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n541), .B2(new_n785), .C1(new_n814), .C2(new_n790), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT48), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT49), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n394), .B1(new_n809), .B2(new_n799), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G116), .B2(new_n1069), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1105), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1094), .B1(new_n1117), .B2(new_n770), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1032), .A2(new_n759), .B1(new_n1082), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n755), .A2(new_n1032), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n705), .B1(new_n754), .B2(new_n1033), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(G393));
  NOR2_X1   g0922(.A1(new_n754), .A2(new_n1033), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1123), .A2(new_n705), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n771), .B1(new_n205), .B2(new_n226), .C1(new_n1052), .C2(new_n242), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT113), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(new_n761), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n814), .A2(new_n257), .B1(new_n1059), .B2(new_n789), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT115), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n817), .A2(new_n211), .B1(new_n202), .B2(new_n795), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n394), .B1(G143), .B2(new_n800), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n847), .A2(G68), .B1(new_n1069), .B2(G87), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n785), .C2(new_n260), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n814), .A2(new_n1067), .B1(new_n786), .B2(new_n789), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT52), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n268), .B(new_n825), .C1(G322), .C2(new_n800), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n806), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(G116), .B1(new_n847), .B2(G283), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n541), .C2(new_n795), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G294), .B2(new_n784), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1131), .A2(new_n1136), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1127), .B1(new_n1077), .B2(new_n1007), .C1(new_n1144), .C2(new_n838), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1121), .A2(new_n758), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1044), .B(new_n699), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1124), .B(new_n1145), .C1(new_n1146), .C2(new_n1148), .ZN(G390));
  XOR2_X1   g0949(.A(new_n954), .B(KEYINPUT116), .Z(new_n1150));
  NAND2_X1  g0950(.A1(new_n950), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n863), .B1(new_n723), .B2(new_n872), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n937), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n952), .A2(new_n953), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n937), .B1(new_n878), .B2(new_n870), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n955), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n749), .A2(G330), .A3(new_n872), .A4(new_n938), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1154), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g0961(.A(G330), .B(new_n872), .C1(new_n982), .C2(new_n985), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n937), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1158), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n878), .A2(new_n870), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n719), .A2(new_n716), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n717), .B1(new_n672), .B2(new_n718), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n722), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n690), .A3(new_n872), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1170), .A2(new_n870), .A3(new_n1158), .A4(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n752), .A2(new_n972), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n897), .A2(new_n1172), .A3(new_n654), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n706), .B1(new_n1161), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT117), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1158), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n952), .A2(new_n953), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1165), .A2(new_n938), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1180), .B2(new_n954), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1170), .A2(new_n870), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1151), .B1(new_n1182), .B2(new_n938), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1178), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1154), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1177), .B1(new_n1186), .B2(new_n1174), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1177), .B(new_n1174), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1176), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1179), .A2(new_n764), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1102), .A2(G128), .B1(G132), .B2(new_n788), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT118), .Z(new_n1193));
  NOR3_X1   g0993(.A1(new_n792), .A2(KEYINPUT53), .A3(new_n257), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n309), .B1(new_n800), .B2(G125), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT53), .B1(new_n792), .B2(new_n257), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n202), .C2(new_n803), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT54), .B(G143), .Z(new_n1198));
  NAND2_X1  g0998(.A1(new_n784), .A2(new_n1198), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n841), .B2(new_n795), .C1(new_n817), .C2(new_n1059), .ZN(new_n1200));
  NOR4_X1   g1000(.A1(new_n1193), .A2(new_n1194), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G116), .A2(new_n788), .B1(new_n796), .B2(G107), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n205), .B2(new_n785), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n268), .B(new_n826), .C1(G294), .C2(new_n800), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n359), .B2(new_n803), .C1(new_n211), .C2(new_n817), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G283), .C2(new_n1102), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n770), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n856), .A2(new_n260), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(new_n760), .A3(new_n1208), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1186), .A2(new_n758), .B1(new_n1191), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1190), .A2(new_n1211), .ZN(G378));
  INV_X1    g1012(.A(KEYINPUT57), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n897), .A2(new_n654), .A3(new_n1173), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1161), .B2(new_n1175), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT120), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n975), .A2(new_n987), .A3(new_n1216), .A4(new_n751), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n959), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n971), .A2(KEYINPUT120), .A3(G330), .A4(new_n973), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n957), .B1(new_n1156), .B2(new_n928), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n956), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n971), .A2(G330), .A3(new_n973), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n263), .A2(new_n681), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n304), .B(new_n1224), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1223), .A2(new_n1216), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1222), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1218), .A2(new_n1229), .A3(new_n1221), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1213), .B1(new_n1215), .B2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1218), .A2(new_n1229), .A3(new_n1221), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1229), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1214), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1186), .B2(new_n1174), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1239), .A3(KEYINPUT57), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1234), .A2(new_n705), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1228), .A2(new_n763), .A3(new_n1227), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n428), .A2(G41), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G33), .A2(G41), .ZN(new_n1244));
  OR3_X1    g1044(.A1(new_n1243), .A2(G50), .A3(new_n1244), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G77), .A2(new_n847), .B1(new_n800), .B2(G283), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1246), .B(new_n1243), .C1(new_n380), .C2(new_n803), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n784), .A2(new_n477), .B1(new_n788), .B2(G107), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n1058), .C1(new_n205), .C2(new_n795), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1247), .B(new_n1249), .C1(G116), .C2(new_n1102), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1245), .B1(new_n1250), .B2(KEYINPUT58), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT119), .Z(new_n1252));
  OAI22_X1  g1052(.A1(new_n817), .A2(new_n257), .B1(new_n785), .B2(new_n841), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(G128), .B2(new_n788), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1102), .A2(G125), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n796), .A2(G132), .B1(new_n847), .B2(new_n1198), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(KEYINPUT59), .ZN(new_n1258));
  INV_X1    g1058(.A(G124), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1244), .B1(new_n799), .B2(new_n1259), .C1(new_n1059), .C2(new_n803), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1257), .B2(KEYINPUT59), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1258), .A2(new_n1261), .B1(new_n1250), .B2(KEYINPUT58), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n838), .B1(new_n1252), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n761), .B(new_n1263), .C1(new_n202), .C2(new_n856), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1237), .A2(new_n759), .B1(new_n1242), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1241), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT121), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(G375));
  INV_X1    g1068(.A(new_n1172), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1214), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n1027), .A3(new_n1174), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n785), .A2(new_n206), .B1(new_n458), .B2(new_n795), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1102), .B2(G294), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT122), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n789), .A2(new_n802), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n268), .B1(new_n800), .B2(G303), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1276), .B1(new_n211), .B2(new_n803), .C1(new_n205), .C2(new_n792), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(new_n1274), .A2(new_n1099), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n394), .B1(G128), .B2(new_n800), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n847), .A2(G159), .B1(new_n1069), .B2(G58), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1279), .B(new_n1280), .C1(new_n785), .C2(new_n257), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G50), .B2(new_n816), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G137), .A2(new_n788), .B1(new_n796), .B2(new_n1198), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n814), .B2(new_n845), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1282), .B1(new_n1284), .B2(KEYINPUT123), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(KEYINPUT123), .B2(new_n1284), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n770), .B1(new_n1278), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n761), .B1(new_n856), .B2(new_n359), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1287), .B(new_n1288), .C1(new_n938), .C2(new_n764), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1172), .B2(new_n759), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1271), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(G381));
  NOR2_X1   g1093(.A1(G375), .A2(G378), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  OAI211_X1 g1095(.A(new_n836), .B(new_n1119), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(G381), .A2(G390), .A3(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1294), .A2(new_n1295), .A3(new_n1080), .A4(new_n1297), .ZN(G407));
  NAND2_X1  g1098(.A1(new_n682), .A2(G213), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1294), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(G407), .A2(G213), .A3(new_n1301), .ZN(G409));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1051), .B2(new_n1079), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1296), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1305), .B(new_n1296), .C1(new_n1051), .C2(new_n1079), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1307), .A2(G390), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1241), .A2(G378), .A3(new_n1265), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1237), .A2(new_n1239), .A3(new_n1027), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1265), .A2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(KEYINPUT117), .B1(new_n1161), .B2(new_n1175), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1188), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1210), .B1(new_n1316), .B2(new_n1176), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1300), .B1(new_n1312), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1174), .A2(KEYINPUT60), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1320), .A2(new_n1270), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1214), .A2(new_n1269), .A3(KEYINPUT60), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n705), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1291), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1295), .ZN(new_n1325));
  OAI211_X1 g1125(.A(G384), .B(new_n1291), .C1(new_n1321), .C2(new_n1323), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1319), .A2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1311), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1327), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1319), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1300), .A2(KEYINPUT124), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1325), .A2(new_n1326), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1300), .A2(G2897), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1325), .A2(new_n1326), .A3(new_n1335), .A4(new_n1333), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1332), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1330), .A2(new_n1331), .A3(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1319), .A2(new_n1327), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1319), .B2(new_n1339), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT126), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(KEYINPUT62), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1319), .B2(new_n1327), .ZN(new_n1349));
  NOR3_X1   g1149(.A1(new_n1344), .A2(new_n1346), .A3(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1310), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1307), .A2(G390), .A3(new_n1308), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1342), .B1(new_n1350), .B2(new_n1353), .ZN(G405));
  NOR2_X1   g1154(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1355), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1351), .B(new_n1352), .C1(KEYINPUT127), .C2(new_n1327), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1317), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1360));
  AND2_X1   g1160(.A1(new_n1360), .A2(new_n1312), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1358), .A2(new_n1362), .ZN(new_n1363));
  NAND4_X1  g1163(.A1(new_n1356), .A2(new_n1359), .A3(new_n1361), .A4(new_n1357), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(G402));
endmodule


