

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  NOR2_X1 U323 ( .A1(n439), .A2(n438), .ZN(n440) );
  NOR2_X2 U324 ( .A1(n443), .A2(n529), .ZN(n567) );
  XOR2_X1 U325 ( .A(n414), .B(n413), .Z(n575) );
  XNOR2_X1 U326 ( .A(G1GAT), .B(G57GAT), .ZN(n335) );
  NOR2_X2 U327 ( .A1(n446), .A2(n455), .ZN(n563) );
  XNOR2_X1 U328 ( .A(n440), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U329 ( .A(n309), .B(n341), .Z(n531) );
  XNOR2_X1 U330 ( .A(n349), .B(n348), .ZN(n529) );
  XNOR2_X1 U331 ( .A(n402), .B(KEYINPUT72), .ZN(n403) );
  XNOR2_X1 U332 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U333 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U334 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  XOR2_X1 U335 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n292) );
  XNOR2_X1 U336 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U338 ( .A(KEYINPUT19), .B(n293), .Z(n362) );
  XOR2_X1 U339 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U342 ( .A(G176GAT), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U343 ( .A(G15GAT), .B(KEYINPUT64), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U345 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n410) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G134GAT), .Z(n375) );
  XOR2_X1 U348 ( .A(n410), .B(n375), .Z(n301) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(n302), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n362), .B(n305), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT81), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT82), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(n308), .ZN(n341) );
  INV_X1 U358 ( .A(n531), .ZN(n455) );
  XOR2_X1 U359 ( .A(G141GAT), .B(G22GAT), .Z(n418) );
  XOR2_X1 U360 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n311) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(KEYINPUT86), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(n418), .B(n312), .Z(n314) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n330) );
  XOR2_X1 U366 ( .A(G204GAT), .B(KEYINPUT22), .Z(n316) );
  XNOR2_X1 U367 ( .A(KEYINPUT87), .B(KEYINPUT23), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n319) );
  XOR2_X1 U369 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n404) );
  XOR2_X1 U372 ( .A(n319), .B(n404), .Z(n328) );
  XOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT3), .Z(n321) );
  XNOR2_X1 U374 ( .A(KEYINPUT89), .B(KEYINPUT2), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U376 ( .A(n322), .B(KEYINPUT88), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT90), .B(G162GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n342) );
  XOR2_X1 U379 ( .A(G211GAT), .B(KEYINPUT21), .Z(n326) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(G218GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n356) );
  XNOR2_X1 U382 ( .A(n342), .B(n356), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n459) );
  XOR2_X1 U385 ( .A(G148GAT), .B(G120GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(G134GAT), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U388 ( .A(G29GAT), .B(G85GAT), .Z(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n347) );
  XOR2_X1 U390 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n336) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U392 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n338) );
  XNOR2_X1 U393 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n340), .B(n339), .Z(n345) );
  INV_X1 U396 ( .A(n341), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n349) );
  NAND2_X1 U400 ( .A1(G225GAT), .A2(G233GAT), .ZN(n348) );
  INV_X1 U401 ( .A(KEYINPUT54), .ZN(n442) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G64GAT), .Z(n351) );
  XNOR2_X1 U403 ( .A(G176GAT), .B(KEYINPUT74), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U405 ( .A(G204GAT), .B(n352), .Z(n414) );
  XOR2_X1 U406 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n354) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n414), .B(n355), .ZN(n360) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XOR2_X1 U411 ( .A(n356), .B(n421), .Z(n358) );
  NAND2_X1 U412 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U414 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n476) );
  XOR2_X1 U416 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n364) );
  XNOR2_X1 U417 ( .A(G218GAT), .B(KEYINPUT66), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n380) );
  XOR2_X1 U419 ( .A(G99GAT), .B(G85GAT), .Z(n399) );
  XOR2_X1 U420 ( .A(n399), .B(G92GAT), .Z(n366) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n368) );
  XNOR2_X1 U424 ( .A(G162GAT), .B(G106GAT), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U426 ( .A(n370), .B(n369), .Z(n378) );
  XOR2_X1 U427 ( .A(G29GAT), .B(KEYINPUT7), .Z(n372) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G36GAT), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U430 ( .A(G50GAT), .B(KEYINPUT8), .Z(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n427) );
  INV_X1 U432 ( .A(n427), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(n380), .B(n379), .Z(n468) );
  XOR2_X1 U436 ( .A(G78GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G155GAT), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U439 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n384) );
  XNOR2_X1 U440 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n383) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n397) );
  XOR2_X1 U443 ( .A(G57GAT), .B(KEYINPUT13), .Z(n398) );
  XOR2_X1 U444 ( .A(G71GAT), .B(G127GAT), .Z(n388) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G183GAT), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U447 ( .A(n398), .B(n389), .Z(n391) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U450 ( .A(n392), .B(KEYINPUT79), .Z(n395) );
  XNOR2_X1 U451 ( .A(G15GAT), .B(G1GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n393), .B(KEYINPUT70), .ZN(n417) );
  XNOR2_X1 U453 ( .A(n417), .B(KEYINPUT78), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n578) );
  XOR2_X1 U456 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n430) );
  XOR2_X1 U457 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n401) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U459 ( .A(n401), .B(n400), .Z(n406) );
  AND2_X1 U460 ( .A1(G230GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n412) );
  XOR2_X1 U462 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n407) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U467 ( .A(KEYINPUT41), .B(n575), .Z(n552) );
  XOR2_X1 U468 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n416) );
  XNOR2_X1 U469 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n426) );
  XOR2_X1 U471 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U472 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U474 ( .A(n422), .B(n421), .Z(n424) );
  XNOR2_X1 U475 ( .A(G113GAT), .B(G197GAT), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U478 ( .A(n428), .B(n427), .Z(n570) );
  AND2_X1 U479 ( .A1(n552), .A2(n570), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n430), .B(n429), .ZN(n431) );
  NOR2_X1 U481 ( .A1(n578), .A2(n431), .ZN(n432) );
  NAND2_X1 U482 ( .A1(n468), .A2(n432), .ZN(n433) );
  XNOR2_X1 U483 ( .A(KEYINPUT47), .B(n433), .ZN(n439) );
  XOR2_X1 U484 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n435) );
  INV_X1 U485 ( .A(n468), .ZN(n564) );
  XNOR2_X1 U486 ( .A(KEYINPUT36), .B(n564), .ZN(n581) );
  NAND2_X1 U487 ( .A1(n578), .A2(n581), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U489 ( .A(n570), .ZN(n498) );
  XOR2_X1 U490 ( .A(KEYINPUT71), .B(n498), .Z(n534) );
  NAND2_X1 U491 ( .A1(n436), .A2(n534), .ZN(n437) );
  NOR2_X1 U492 ( .A1(n575), .A2(n437), .ZN(n438) );
  NOR2_X1 U493 ( .A1(n476), .A2(n527), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U495 ( .A1(n459), .A2(n567), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n444), .B(KEYINPUT123), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U498 ( .A1(n563), .A2(n552), .ZN(n450) );
  XOR2_X1 U499 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n448) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n447) );
  XOR2_X1 U501 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n474) );
  XNOR2_X1 U502 ( .A(KEYINPUT27), .B(KEYINPUT96), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(n476), .ZN(n526) );
  XNOR2_X1 U504 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(n459), .ZN(n530) );
  NOR2_X1 U506 ( .A1(n526), .A2(n530), .ZN(n453) );
  NAND2_X1 U507 ( .A1(n455), .A2(n453), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n454), .A2(n529), .ZN(n466) );
  INV_X1 U509 ( .A(n459), .ZN(n457) );
  NOR2_X1 U510 ( .A1(n455), .A2(n476), .ZN(n456) );
  NOR2_X1 U511 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(KEYINPUT25), .B(n458), .ZN(n464) );
  NOR2_X1 U513 ( .A1(n531), .A2(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(n568) );
  NOR2_X1 U516 ( .A1(n568), .A2(n526), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n529), .A2(n462), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U520 ( .A(KEYINPUT98), .B(n467), .ZN(n483) );
  NAND2_X1 U521 ( .A1(n578), .A2(n468), .ZN(n469) );
  XNOR2_X1 U522 ( .A(n469), .B(KEYINPUT80), .ZN(n470) );
  XNOR2_X1 U523 ( .A(n470), .B(KEYINPUT16), .ZN(n471) );
  NOR2_X1 U524 ( .A1(n483), .A2(n471), .ZN(n499) );
  NOR2_X1 U525 ( .A1(n575), .A2(n534), .ZN(n487) );
  NAND2_X1 U526 ( .A1(n499), .A2(n487), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT99), .ZN(n480) );
  NAND2_X1 U528 ( .A1(n480), .A2(n529), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n475), .Z(G1324GAT) );
  INV_X1 U531 ( .A(n476), .ZN(n516) );
  NAND2_X1 U532 ( .A1(n480), .A2(n516), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U535 ( .A1(n480), .A2(n531), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT101), .Z(n482) );
  NAND2_X1 U538 ( .A1(n480), .A2(n530), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  NOR2_X1 U540 ( .A1(n578), .A2(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT102), .B(n484), .ZN(n485) );
  NAND2_X1 U542 ( .A1(n485), .A2(n581), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(KEYINPUT37), .ZN(n511) );
  NAND2_X1 U544 ( .A1(n511), .A2(n487), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT38), .B(n488), .Z(n495) );
  NAND2_X1 U546 ( .A1(n529), .A2(n495), .ZN(n490) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  XOR2_X1 U549 ( .A(G36GAT), .B(KEYINPUT103), .Z(n492) );
  NAND2_X1 U550 ( .A1(n516), .A2(n495), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1329GAT) );
  NAND2_X1 U552 ( .A1(n495), .A2(n531), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT40), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NAND2_X1 U555 ( .A1(n495), .A2(n530), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(KEYINPUT104), .ZN(n497) );
  XNOR2_X1 U557 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT42), .B(KEYINPUT105), .Z(n502) );
  NAND2_X1 U559 ( .A1(n552), .A2(n498), .ZN(n512) );
  INV_X1 U560 ( .A(n499), .ZN(n500) );
  NOR2_X1 U561 ( .A1(n512), .A2(n500), .ZN(n508) );
  NAND2_X1 U562 ( .A1(n508), .A2(n529), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n508), .A2(n516), .ZN(n504) );
  XNOR2_X1 U566 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U568 ( .A1(n508), .A2(n531), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U572 ( .A1(n508), .A2(n530), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(KEYINPUT108), .ZN(n515) );
  INV_X1 U575 ( .A(n511), .ZN(n513) );
  NOR2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n529), .A2(n521), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  XOR2_X1 U579 ( .A(G92GAT), .B(KEYINPUT109), .Z(n518) );
  NAND2_X1 U580 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n531), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n525) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n530), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n536) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  NAND2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n546) );
  NOR2_X1 U593 ( .A1(n530), .A2(n546), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(KEYINPUT115), .ZN(n543) );
  INV_X1 U596 ( .A(n534), .ZN(n559) );
  NAND2_X1 U597 ( .A1(n543), .A2(n559), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U601 ( .A1(n543), .A2(n552), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n541) );
  NAND2_X1 U604 ( .A1(n543), .A2(n578), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n564), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT119), .Z(n548) );
  NOR2_X1 U611 ( .A1(n568), .A2(n546), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n557), .A2(n570), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT53), .B(n551), .Z(n554) );
  NAND2_X1 U618 ( .A1(n557), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n557), .A2(n578), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT122), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n578), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  INV_X1 U633 ( .A(n567), .ZN(n569) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n582) );
  AND2_X1 U635 ( .A1(n570), .A2(n582), .ZN(n574) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT126), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  AND2_X1 U640 ( .A1(n575), .A2(n582), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  AND2_X1 U643 ( .A1(n578), .A2(n582), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

