

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U550 ( .A(KEYINPUT13), .B(n594), .Z(n517) );
  NOR2_X2 U551 ( .A1(n703), .A2(n702), .ZN(n719) );
  XNOR2_X2 U552 ( .A(KEYINPUT27), .B(n701), .ZN(n702) );
  NAND2_X2 U553 ( .A1(n697), .A2(n787), .ZN(n710) );
  NAND2_X2 U554 ( .A1(n597), .A2(n596), .ZN(n971) );
  NOR2_X2 U555 ( .A1(n595), .A2(n517), .ZN(n597) );
  OR2_X1 U556 ( .A1(n707), .A2(n971), .ZN(n708) );
  XNOR2_X1 U557 ( .A(n520), .B(n519), .ZN(n1002) );
  NOR2_X1 U558 ( .A1(G1966), .A2(n782), .ZN(n741) );
  NAND2_X1 U559 ( .A1(n1002), .A2(G137), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n770), .A2(n769), .ZN(n518) );
  NOR2_X1 U561 ( .A1(n710), .A2(n913), .ZN(n706) );
  NOR2_X1 U562 ( .A1(n709), .A2(n708), .ZN(n716) );
  OR2_X1 U563 ( .A1(n972), .A2(n716), .ZN(n717) );
  BUF_X1 U564 ( .A(n710), .Z(n748) );
  INV_X1 U565 ( .A(n935), .ZN(n769) );
  INV_X1 U566 ( .A(KEYINPUT105), .ZN(n759) );
  INV_X1 U567 ( .A(KEYINPUT106), .ZN(n772) );
  NAND2_X1 U568 ( .A1(G8), .A2(n710), .ZN(n782) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n519) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n656) );
  INV_X1 U571 ( .A(KEYINPUT65), .ZN(n529) );
  XNOR2_X1 U572 ( .A(n530), .B(n529), .ZN(n531) );
  NOR2_X1 U573 ( .A1(n532), .A2(n531), .ZN(n696) );
  BUF_X1 U574 ( .A(n696), .Z(G160) );
  NOR2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n998) );
  NAND2_X1 U577 ( .A1(G113), .A2(n998), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(n523), .ZN(n532) );
  INV_X1 U580 ( .A(G2104), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n526), .A2(G2105), .ZN(n524) );
  XNOR2_X1 U582 ( .A(n524), .B(KEYINPUT64), .ZN(n569) );
  NAND2_X1 U583 ( .A1(n569), .A2(G101), .ZN(n525) );
  XOR2_X1 U584 ( .A(n525), .B(KEYINPUT23), .Z(n528) );
  AND2_X1 U585 ( .A1(n526), .A2(G2105), .ZN(n999) );
  NAND2_X1 U586 ( .A1(n999), .A2(G125), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n530) );
  NAND2_X1 U588 ( .A1(G85), .A2(n656), .ZN(n534) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  INV_X1 U590 ( .A(G651), .ZN(n535) );
  NOR2_X2 U591 ( .A1(n650), .A2(n535), .ZN(n653) );
  NAND2_X1 U592 ( .A1(G72), .A2(n653), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U594 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X2 U595 ( .A(KEYINPUT1), .B(n536), .Z(n655) );
  NAND2_X1 U596 ( .A1(G60), .A2(n655), .ZN(n538) );
  NOR2_X2 U597 ( .A1(G651), .A2(n650), .ZN(n659) );
  NAND2_X1 U598 ( .A1(G47), .A2(n659), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U600 ( .A1(n540), .A2(n539), .ZN(G290) );
  XOR2_X1 U601 ( .A(G2443), .B(G2435), .Z(n542) );
  XNOR2_X1 U602 ( .A(G2451), .B(G2446), .ZN(n541) );
  XNOR2_X1 U603 ( .A(n542), .B(n541), .ZN(n549) );
  XOR2_X1 U604 ( .A(G2427), .B(G2438), .Z(n544) );
  XNOR2_X1 U605 ( .A(G1341), .B(G2430), .ZN(n543) );
  XNOR2_X1 U606 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U607 ( .A(n545), .B(KEYINPUT107), .Z(n547) );
  XNOR2_X1 U608 ( .A(G1348), .B(G2454), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n549), .B(n548), .ZN(n550) );
  AND2_X1 U611 ( .A1(n550), .A2(G14), .ZN(G401) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G120), .ZN(G236) );
  INV_X1 U614 ( .A(G69), .ZN(G235) );
  INV_X1 U615 ( .A(G108), .ZN(G238) );
  NAND2_X1 U616 ( .A1(G64), .A2(n655), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G52), .A2(n659), .ZN(n551) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G90), .A2(n656), .ZN(n554) );
  NAND2_X1 U620 ( .A1(G77), .A2(n653), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U624 ( .A1(n659), .A2(G50), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT79), .B(n558), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n655), .A2(G62), .ZN(n559) );
  XOR2_X1 U627 ( .A(KEYINPUT78), .B(n559), .Z(n560) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT80), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G88), .A2(n656), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G75), .A2(n653), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT81), .B(n565), .ZN(n566) );
  NOR2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT82), .B(n568), .Z(G303) );
  NAND2_X1 U636 ( .A1(n1002), .A2(G138), .ZN(n572) );
  INV_X1 U637 ( .A(n569), .ZN(n570) );
  INV_X1 U638 ( .A(n570), .ZN(n1004) );
  NAND2_X1 U639 ( .A1(G102), .A2(n1004), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G114), .A2(n998), .ZN(n574) );
  NAND2_X1 U642 ( .A1(G126), .A2(n999), .ZN(n573) );
  NAND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U644 ( .A1(n576), .A2(n575), .ZN(G164) );
  NAND2_X1 U645 ( .A1(n656), .A2(G89), .ZN(n577) );
  XNOR2_X1 U646 ( .A(n577), .B(KEYINPUT4), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G76), .A2(n653), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT5), .ZN(n585) );
  NAND2_X1 U650 ( .A1(G63), .A2(n655), .ZN(n582) );
  NAND2_X1 U651 ( .A1(G51), .A2(n659), .ZN(n581) );
  NAND2_X1 U652 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U653 ( .A(KEYINPUT6), .B(n583), .Z(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U656 ( .A(G168), .B(KEYINPUT8), .Z(n587) );
  XNOR2_X1 U657 ( .A(KEYINPUT72), .B(n587), .ZN(G286) );
  NAND2_X1 U658 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U659 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U660 ( .A(G223), .ZN(n838) );
  NAND2_X1 U661 ( .A1(n838), .A2(G567), .ZN(n589) );
  XOR2_X1 U662 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U663 ( .A1(G56), .A2(n655), .ZN(n590) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(n590), .Z(n595) );
  NAND2_X1 U665 ( .A1(n656), .A2(G81), .ZN(n591) );
  XNOR2_X1 U666 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U667 ( .A1(G68), .A2(n653), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n659), .A2(G43), .ZN(n596) );
  INV_X1 U670 ( .A(G860), .ZN(n622) );
  OR2_X1 U671 ( .A1(n971), .A2(n622), .ZN(G153) );
  INV_X1 U672 ( .A(G171), .ZN(G301) );
  NAND2_X1 U673 ( .A1(G868), .A2(G301), .ZN(n611) );
  NAND2_X1 U674 ( .A1(n656), .A2(G92), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT68), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G66), .A2(n655), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U678 ( .A(KEYINPUT69), .B(n601), .Z(n608) );
  NAND2_X1 U679 ( .A1(n653), .A2(G79), .ZN(n602) );
  XNOR2_X1 U680 ( .A(n602), .B(KEYINPUT70), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G54), .A2(n659), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n605), .ZN(n606) );
  INV_X1 U684 ( .A(n606), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X2 U686 ( .A(KEYINPUT15), .B(n609), .Z(n972) );
  OR2_X1 U687 ( .A1(n972), .A2(G868), .ZN(n610) );
  NAND2_X1 U688 ( .A1(n611), .A2(n610), .ZN(G284) );
  NAND2_X1 U689 ( .A1(G65), .A2(n655), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G53), .A2(n659), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U692 ( .A1(G91), .A2(n656), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G78), .A2(n653), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n938) );
  XNOR2_X1 U696 ( .A(n938), .B(KEYINPUT67), .ZN(G299) );
  XNOR2_X1 U697 ( .A(KEYINPUT73), .B(G868), .ZN(n618) );
  NOR2_X1 U698 ( .A1(G286), .A2(n618), .ZN(n619) );
  XNOR2_X1 U699 ( .A(n619), .B(KEYINPUT74), .ZN(n621) );
  NOR2_X1 U700 ( .A1(G299), .A2(G868), .ZN(n620) );
  NOR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(G297) );
  NAND2_X1 U702 ( .A1(n622), .A2(G559), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(n972), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U705 ( .A1(G868), .A2(n971), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n972), .A2(G868), .ZN(n625) );
  NOR2_X1 U707 ( .A1(G559), .A2(n625), .ZN(n626) );
  NOR2_X1 U708 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U709 ( .A1(n998), .A2(G111), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G99), .A2(n1004), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n999), .A2(G123), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n630), .B(KEYINPUT18), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G135), .A2(n1002), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT75), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n994) );
  XNOR2_X1 U718 ( .A(n994), .B(G2096), .ZN(n637) );
  INV_X1 U719 ( .A(G2100), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(G156) );
  NAND2_X1 U721 ( .A1(G67), .A2(n655), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G80), .A2(n653), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n656), .A2(G93), .ZN(n640) );
  XOR2_X1 U725 ( .A(KEYINPUT76), .B(n640), .Z(n641) );
  NOR2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n659), .A2(G55), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n675) );
  NAND2_X1 U729 ( .A1(G559), .A2(n972), .ZN(n645) );
  XNOR2_X1 U730 ( .A(n645), .B(n971), .ZN(n671) );
  NOR2_X1 U731 ( .A1(G860), .A2(n671), .ZN(n646) );
  XOR2_X1 U732 ( .A(n675), .B(n646), .Z(G145) );
  NAND2_X1 U733 ( .A1(G49), .A2(n659), .ZN(n648) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U736 ( .A1(n655), .A2(n649), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n650), .A2(G87), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U739 ( .A1(G73), .A2(n653), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n654), .B(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U741 ( .A1(G61), .A2(n655), .ZN(n658) );
  NAND2_X1 U742 ( .A1(G86), .A2(n656), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U744 ( .A1(G48), .A2(n659), .ZN(n660) );
  XNOR2_X1 U745 ( .A(KEYINPUT77), .B(n660), .ZN(n661) );
  NOR2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n664), .A2(n663), .ZN(G305) );
  XNOR2_X1 U748 ( .A(G290), .B(G288), .ZN(n669) );
  XNOR2_X1 U749 ( .A(G305), .B(G299), .ZN(n667) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n665) );
  XNOR2_X1 U751 ( .A(n665), .B(n675), .ZN(n666) );
  XNOR2_X1 U752 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U753 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U754 ( .A(G303), .B(n670), .ZN(n970) );
  XNOR2_X1 U755 ( .A(KEYINPUT84), .B(n671), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n970), .B(n672), .ZN(n673) );
  NAND2_X1 U757 ( .A1(n673), .A2(G868), .ZN(n677) );
  INV_X1 U758 ( .A(G868), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U764 ( .A(n680), .B(KEYINPUT86), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n681) );
  XNOR2_X1 U766 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U768 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U769 ( .A1(G235), .A2(G236), .ZN(n684) );
  XOR2_X1 U770 ( .A(KEYINPUT88), .B(n684), .Z(n685) );
  NOR2_X1 U771 ( .A1(G238), .A2(n685), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G57), .A2(n686), .ZN(n968) );
  NAND2_X1 U773 ( .A1(G567), .A2(n968), .ZN(n692) );
  XOR2_X1 U774 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n688) );
  NAND2_X1 U775 ( .A1(G132), .A2(G82), .ZN(n687) );
  XNOR2_X1 U776 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n689), .A2(G218), .ZN(n690) );
  NAND2_X1 U778 ( .A1(G96), .A2(n690), .ZN(n969) );
  NAND2_X1 U779 ( .A1(G2106), .A2(n969), .ZN(n691) );
  NAND2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U781 ( .A(KEYINPUT89), .B(n693), .ZN(G319) );
  INV_X1 U782 ( .A(G319), .ZN(n1023) );
  NAND2_X1 U783 ( .A1(G661), .A2(G483), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n1023), .A2(n694), .ZN(n842) );
  NAND2_X1 U785 ( .A1(G36), .A2(n842), .ZN(n695) );
  XNOR2_X1 U786 ( .A(n695), .B(KEYINPUT90), .ZN(G176) );
  NAND2_X1 U787 ( .A1(n696), .A2(G40), .ZN(n786) );
  INV_X1 U788 ( .A(n786), .ZN(n697) );
  NOR2_X1 U789 ( .A1(G164), .A2(G1384), .ZN(n787) );
  AND2_X1 U790 ( .A1(G1956), .A2(n710), .ZN(n699) );
  INV_X1 U791 ( .A(KEYINPUT101), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n699), .B(n698), .ZN(n703) );
  INV_X1 U793 ( .A(n710), .ZN(n700) );
  NAND2_X1 U794 ( .A1(n700), .A2(G2072), .ZN(n701) );
  NOR2_X1 U795 ( .A1(n938), .A2(n719), .ZN(n705) );
  INV_X1 U796 ( .A(KEYINPUT28), .ZN(n704) );
  XNOR2_X1 U797 ( .A(n705), .B(n704), .ZN(n723) );
  INV_X1 U798 ( .A(G1996), .ZN(n913) );
  XNOR2_X1 U799 ( .A(n706), .B(KEYINPUT26), .ZN(n709) );
  AND2_X1 U800 ( .A1(n710), .A2(G1341), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n972), .A2(n716), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n748), .A2(G1348), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(KEYINPUT102), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n700), .A2(G2067), .ZN(n712) );
  NAND2_X1 U805 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U808 ( .A1(n938), .A2(n719), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U811 ( .A(n724), .B(KEYINPUT29), .ZN(n729) );
  XOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .Z(n911) );
  NOR2_X1 U813 ( .A1(n911), .A2(n748), .ZN(n725) );
  XNOR2_X1 U814 ( .A(n725), .B(KEYINPUT100), .ZN(n727) );
  XOR2_X1 U815 ( .A(G1961), .B(KEYINPUT99), .Z(n904) );
  NOR2_X1 U816 ( .A1(n700), .A2(n904), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n733) );
  NOR2_X1 U818 ( .A1(G301), .A2(n733), .ZN(n728) );
  NOR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n738) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n748), .ZN(n743) );
  NOR2_X1 U821 ( .A1(n743), .A2(n741), .ZN(n730) );
  NAND2_X1 U822 ( .A1(G8), .A2(n730), .ZN(n731) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n731), .ZN(n732) );
  NOR2_X1 U824 ( .A1(n732), .A2(G168), .ZN(n735) );
  AND2_X1 U825 ( .A1(G301), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U827 ( .A(n736), .B(KEYINPUT31), .ZN(n737) );
  NOR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U829 ( .A(n739), .B(KEYINPUT103), .ZN(n747) );
  INV_X1 U830 ( .A(n747), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U832 ( .A(n742), .B(KEYINPUT104), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n743), .A2(G8), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n758) );
  AND2_X1 U835 ( .A1(G286), .A2(G8), .ZN(n746) );
  NAND2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n755) );
  INV_X1 U837 ( .A(G8), .ZN(n753) );
  NOR2_X1 U838 ( .A1(G1971), .A2(n782), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n751), .A2(G303), .ZN(n752) );
  OR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U846 ( .A(n760), .B(n759), .ZN(n779) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n939) );
  NOR2_X1 U848 ( .A1(G303), .A2(G1971), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n939), .A2(n761), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n779), .A2(n762), .ZN(n763) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n940) );
  NAND2_X1 U852 ( .A1(n763), .A2(n940), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n782), .A2(n764), .ZN(n765) );
  INV_X1 U854 ( .A(n765), .ZN(n767) );
  INV_X1 U855 ( .A(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n939), .A2(KEYINPUT33), .ZN(n768) );
  NOR2_X1 U858 ( .A1(n768), .A2(n782), .ZN(n770) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n935) );
  NAND2_X1 U860 ( .A1(n771), .A2(n518), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(n772), .ZN(n778) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U863 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  NOR2_X1 U864 ( .A1(n782), .A2(n775), .ZN(n776) );
  XNOR2_X1 U865 ( .A(n776), .B(KEYINPUT98), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n778), .A2(n777), .ZN(n785) );
  NOR2_X1 U867 ( .A1(G2090), .A2(G303), .ZN(n780) );
  NAND2_X1 U868 ( .A1(G8), .A2(n780), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n779), .A2(n781), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n823) );
  XNOR2_X1 U872 ( .A(G1986), .B(G290), .ZN(n944) );
  NOR2_X1 U873 ( .A1(n787), .A2(n786), .ZN(n833) );
  NAND2_X1 U874 ( .A1(n944), .A2(n833), .ZN(n821) );
  NAND2_X1 U875 ( .A1(n1002), .A2(G140), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G104), .A2(n1004), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U878 ( .A(n790), .B(KEYINPUT91), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n791), .B(KEYINPUT34), .ZN(n797) );
  XNOR2_X1 U880 ( .A(KEYINPUT35), .B(KEYINPUT92), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G116), .A2(n998), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G128), .A2(n999), .ZN(n792) );
  NAND2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U884 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U886 ( .A(KEYINPUT36), .B(n798), .Z(n1016) );
  XNOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NOR2_X1 U888 ( .A1(n1016), .A2(n831), .ZN(n851) );
  NAND2_X1 U889 ( .A1(n851), .A2(n833), .ZN(n799) );
  XOR2_X1 U890 ( .A(KEYINPUT93), .B(n799), .Z(n829) );
  NAND2_X1 U891 ( .A1(n999), .A2(G119), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G95), .A2(n1004), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n998), .A2(G107), .ZN(n802) );
  XOR2_X1 U895 ( .A(KEYINPUT94), .B(n802), .Z(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n1002), .A2(G131), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n1010) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n1010), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT95), .ZN(n817) );
  NAND2_X1 U901 ( .A1(n1004), .A2(G105), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT38), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G141), .A2(n1002), .ZN(n810) );
  NAND2_X1 U904 ( .A1(G117), .A2(n998), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n999), .A2(G129), .ZN(n811) );
  XOR2_X1 U907 ( .A(KEYINPUT96), .B(n811), .Z(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n995) );
  AND2_X1 U910 ( .A1(G1996), .A2(n995), .ZN(n816) );
  NOR2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n853) );
  XNOR2_X1 U912 ( .A(KEYINPUT97), .B(n833), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n853), .A2(n818), .ZN(n826) );
  INV_X1 U914 ( .A(n826), .ZN(n819) );
  AND2_X1 U915 ( .A1(n829), .A2(n819), .ZN(n820) );
  AND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n836) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n995), .ZN(n855) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n824) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n1010), .ZN(n870) );
  NOR2_X1 U921 ( .A1(n824), .A2(n870), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  NOR2_X1 U923 ( .A1(n855), .A2(n827), .ZN(n828) );
  XNOR2_X1 U924 ( .A(n828), .B(KEYINPUT39), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n1016), .A2(n831), .ZN(n868) );
  NAND2_X1 U927 ( .A1(n832), .A2(n868), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT108), .B(n839), .Z(n840) );
  NAND2_X1 U934 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(G188) );
  NAND2_X1 U938 ( .A1(G124), .A2(n999), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U940 ( .A1(n1004), .A2(G100), .ZN(n844) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(n844), .Z(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G136), .A2(n1002), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G112), .A2(n998), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G162) );
  INV_X1 U947 ( .A(n851), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(n879) );
  XOR2_X1 U949 ( .A(G2090), .B(G162), .Z(n854) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U951 ( .A(KEYINPUT51), .B(n856), .Z(n877) );
  NAND2_X1 U952 ( .A1(n1002), .A2(G139), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G103), .A2(n1004), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U955 ( .A1(G115), .A2(n998), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G127), .A2(n999), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT47), .B(n861), .ZN(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(n862), .ZN(n863) );
  NOR2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n1015) );
  XOR2_X1 U961 ( .A(G2072), .B(n1015), .Z(n866) );
  XOR2_X1 U962 ( .A(G164), .B(G2078), .Z(n865) );
  NOR2_X1 U963 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U964 ( .A(n867), .B(KEYINPUT50), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n875) );
  XNOR2_X1 U966 ( .A(G160), .B(G2084), .ZN(n872) );
  NOR2_X1 U967 ( .A1(n870), .A2(n994), .ZN(n871) );
  NAND2_X1 U968 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U969 ( .A(KEYINPUT115), .B(n873), .Z(n874) );
  NOR2_X1 U970 ( .A1(n875), .A2(n874), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT52), .B(n880), .ZN(n882) );
  INV_X1 U974 ( .A(KEYINPUT55), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n883), .A2(G29), .ZN(n966) );
  XNOR2_X1 U977 ( .A(G1971), .B(G22), .ZN(n885) );
  XNOR2_X1 U978 ( .A(G23), .B(G1976), .ZN(n884) );
  NOR2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n887) );
  XOR2_X1 U980 ( .A(G1986), .B(G24), .Z(n886) );
  NAND2_X1 U981 ( .A1(n887), .A2(n886), .ZN(n889) );
  XOR2_X1 U982 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n888) );
  XNOR2_X1 U983 ( .A(n889), .B(n888), .ZN(n903) );
  XOR2_X1 U984 ( .A(G4), .B(KEYINPUT125), .Z(n891) );
  XNOR2_X1 U985 ( .A(G1348), .B(KEYINPUT59), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n895) );
  XNOR2_X1 U987 ( .A(G1956), .B(G20), .ZN(n893) );
  XNOR2_X1 U988 ( .A(G19), .B(G1341), .ZN(n892) );
  NOR2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n898) );
  XNOR2_X1 U991 ( .A(KEYINPUT124), .B(G1981), .ZN(n896) );
  XNOR2_X1 U992 ( .A(G6), .B(n896), .ZN(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT60), .B(n899), .Z(n901) );
  XNOR2_X1 U995 ( .A(G1966), .B(G21), .ZN(n900) );
  NOR2_X1 U996 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n903), .A2(n902), .ZN(n906) );
  XNOR2_X1 U998 ( .A(G5), .B(n904), .ZN(n905) );
  NOR2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(KEYINPUT61), .B(n907), .ZN(n909) );
  INV_X1 U1001 ( .A(G16), .ZN(n908) );
  NAND2_X1 U1002 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(n910), .A2(G11), .ZN(n964) );
  XOR2_X1 U1004 ( .A(n911), .B(G27), .Z(n923) );
  XNOR2_X1 U1005 ( .A(KEYINPUT117), .B(G2072), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(G33), .ZN(n918) );
  XNOR2_X1 U1007 ( .A(G32), .B(n913), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n914), .A2(G28), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(G25), .B(G1991), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(n921) );
  XNOR2_X1 U1012 ( .A(KEYINPUT116), .B(G2067), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(G26), .B(n919), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1016 ( .A(KEYINPUT53), .B(n924), .ZN(n928) );
  XOR2_X1 U1017 ( .A(KEYINPUT118), .B(G34), .Z(n926) );
  XNOR2_X1 U1018 ( .A(G2084), .B(KEYINPUT54), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G35), .B(G2090), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1023 ( .A(KEYINPUT55), .B(n931), .Z(n932) );
  NOR2_X1 U1024 ( .A1(G29), .A2(n932), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(n933), .ZN(n962) );
  XOR2_X1 U1026 ( .A(G16), .B(KEYINPUT56), .Z(n959) );
  XNOR2_X1 U1027 ( .A(G1966), .B(G168), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(n934), .B(KEYINPUT120), .ZN(n936) );
  NAND2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(n937), .B(KEYINPUT57), .ZN(n954) );
  XNOR2_X1 U1031 ( .A(G171), .B(G1961), .ZN(n950) );
  XNOR2_X1 U1032 ( .A(n938), .B(G1956), .ZN(n946) );
  INV_X1 U1033 ( .A(n939), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1035 ( .A(KEYINPUT121), .B(n942), .Z(n943) );
  NOR2_X1 U1036 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1038 ( .A(G1341), .B(n971), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1040 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(G1971), .B(G303), .ZN(n951) );
  NOR2_X1 U1042 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1043 ( .A1(n954), .A2(n953), .ZN(n956) );
  XOR2_X1 U1044 ( .A(G1348), .B(n972), .Z(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1046 ( .A(KEYINPUT122), .B(n957), .ZN(n958) );
  NOR2_X1 U1047 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(KEYINPUT123), .B(n960), .ZN(n961) );
  NAND2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1050 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1051 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1052 ( .A(KEYINPUT62), .B(n967), .Z(G311) );
  XNOR2_X1 U1053 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1054 ( .A(G132), .ZN(G219) );
  INV_X1 U1055 ( .A(G96), .ZN(G221) );
  INV_X1 U1056 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1057 ( .A1(n969), .A2(n968), .ZN(G325) );
  INV_X1 U1058 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1059 ( .A(n971), .B(n970), .ZN(n974) );
  XNOR2_X1 U1060 ( .A(G171), .B(n972), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1062 ( .A(n975), .B(G286), .Z(n976) );
  NOR2_X1 U1063 ( .A1(G37), .A2(n976), .ZN(G397) );
  XOR2_X1 U1064 ( .A(G2100), .B(G2096), .Z(n978) );
  XNOR2_X1 U1065 ( .A(G2072), .B(G2090), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n978), .B(n977), .ZN(n982) );
  XOR2_X1 U1067 ( .A(G2678), .B(KEYINPUT42), .Z(n980) );
  XNOR2_X1 U1068 ( .A(G2067), .B(KEYINPUT43), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1070 ( .A(n982), .B(n981), .Z(n984) );
  XNOR2_X1 U1071 ( .A(G2084), .B(G2078), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n984), .B(n983), .ZN(G227) );
  XOR2_X1 U1073 ( .A(G1976), .B(G1971), .Z(n986) );
  XNOR2_X1 U1074 ( .A(G1986), .B(G1966), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n986), .B(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(n987), .B(G2474), .Z(n989) );
  XNOR2_X1 U1077 ( .A(G1996), .B(G1956), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(n989), .B(n988), .ZN(n993) );
  XOR2_X1 U1079 ( .A(KEYINPUT41), .B(G1981), .Z(n991) );
  XNOR2_X1 U1080 ( .A(G1991), .B(G1961), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n991), .B(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n993), .B(n992), .ZN(G229) );
  XOR2_X1 U1083 ( .A(n994), .B(G162), .Z(n997) );
  XOR2_X1 U1084 ( .A(G160), .B(n995), .Z(n996) );
  XNOR2_X1 U1085 ( .A(n997), .B(n996), .ZN(n1021) );
  NAND2_X1 U1086 ( .A1(G118), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(G130), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1009) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(G142), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(KEYINPUT110), .ZN(n1006) );
  NAND2_X1 U1091 ( .A1(G106), .A2(n1004), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(KEYINPUT45), .B(n1007), .Z(n1008) );
  NOR2_X1 U1094 ( .A1(n1009), .A2(n1008), .ZN(n1014) );
  XNOR2_X1 U1095 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1010), .B(KEYINPUT112), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1014), .B(n1013), .ZN(n1019) );
  XNOR2_X1 U1099 ( .A(G164), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1100 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(n1019), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1022), .ZN(G395) );
  NOR2_X1 U1104 ( .A1(G401), .A2(n1023), .ZN(n1028) );
  NOR2_X1 U1105 ( .A1(G227), .A2(G229), .ZN(n1024) );
  XOR2_X1 U1106 ( .A(KEYINPUT113), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1107 ( .A(n1025), .B(KEYINPUT49), .ZN(n1026) );
  NOR2_X1 U1108 ( .A1(G397), .A2(n1026), .ZN(n1027) );
  NAND2_X1 U1109 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1110 ( .A1(n1029), .A2(G395), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(n1030), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1112 ( .A(G308), .ZN(G225) );
  INV_X1 U1113 ( .A(G57), .ZN(G237) );
  INV_X1 U1114 ( .A(G303), .ZN(G166) );
endmodule

