//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XOR2_X1   g0006(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT66), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n208), .B(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  INV_X1    g0019(.A(new_n201), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n215), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT67), .B(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n223), .B1(KEYINPUT1), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n217), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G274), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n258), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n259), .B1(G226), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G222), .A2(G1698), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G223), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n256), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n270), .B(new_n271), .C1(G77), .C2(new_n266), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G190), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n202), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n211), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n218), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n209), .B2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n279), .B1(new_n283), .B2(new_n202), .ZN(new_n284));
  INV_X1    g0084(.A(new_n281), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT8), .A2(G58), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT71), .B(G58), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(KEYINPUT8), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n254), .A2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n285), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n276), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n297), .B1(new_n298), .B2(KEYINPUT10), .C1(new_n299), .C2(new_n273), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT10), .B1(new_n297), .B2(new_n298), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n299), .B2(new_n273), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n273), .A2(G169), .ZN(new_n304));
  INV_X1    g0104(.A(G179), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n273), .ZN(new_n306));
  INV_X1    g0106(.A(new_n294), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(G77), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n289), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT8), .B(G58), .Z(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n309), .B1(G77), .B2(new_n277), .C1(new_n315), .C2(new_n285), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n260), .A2(new_n224), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n266), .A2(G232), .A3(new_n268), .ZN(new_n318));
  INV_X1    g0118(.A(G107), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n266), .A2(G1698), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n318), .B1(new_n319), .B2(new_n266), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  AOI211_X1 g0122(.A(new_n259), .B(new_n317), .C1(new_n322), .C2(new_n271), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n316), .B1(G190), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n299), .B2(new_n323), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n305), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n316), .B(new_n326), .C1(G169), .C2(new_n323), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AND4_X1   g0128(.A1(new_n300), .A2(new_n303), .A3(new_n308), .A4(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(G226), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(G232), .B2(new_n268), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n264), .A2(new_n265), .ZN(new_n332));
  INV_X1    g0132(.A(G97), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n331), .A2(new_n332), .B1(new_n254), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n259), .B1(new_n334), .B2(new_n271), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n321), .B1(new_n260), .B2(KEYINPUT74), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(KEYINPUT74), .B2(new_n260), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT13), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT14), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(G179), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n344), .A3(G169), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n343), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G68), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n291), .A2(G50), .B1(G20), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n289), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n225), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n354), .A2(new_n281), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT12), .B1(new_n277), .B2(G68), .ZN(new_n357));
  OR3_X1    g0157(.A1(new_n277), .A2(KEYINPUT12), .A3(G68), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n282), .A2(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g0161(.A(new_n361), .B(KEYINPUT75), .Z(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT77), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n350), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n362), .B1(new_n275), .B2(new_n339), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n340), .A2(new_n299), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n329), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n288), .A2(new_n278), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n370), .B1(new_n283), .B2(new_n288), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT71), .A2(G58), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT71), .A2(G58), .ZN(new_n373));
  OAI21_X1  g0173(.A(G68), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n210), .B1(new_n374), .B2(new_n220), .ZN(new_n375));
  INV_X1    g0175(.A(new_n291), .ZN(new_n376));
  INV_X1    g0176(.A(G159), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT80), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT80), .ZN(new_n380));
  INV_X1    g0180(.A(new_n378), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n201), .B1(new_n287), .B2(G68), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n380), .B(new_n381), .C1(new_n382), .C2(new_n210), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  AND2_X1   g0186(.A1(KEYINPUT78), .A2(G33), .ZN(new_n387));
  NOR2_X1   g0187(.A1(KEYINPUT78), .A2(G33), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n387), .A2(new_n388), .A3(new_n263), .ZN(new_n389));
  INV_X1    g0189(.A(new_n264), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n386), .B(new_n210), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT79), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n254), .ZN(new_n395));
  NAND2_X1  g0195(.A1(KEYINPUT78), .A2(G33), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT3), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n264), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n386), .B1(new_n398), .B2(new_n210), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n392), .A2(new_n393), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(G20), .B1(new_n397), .B2(new_n264), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n351), .B1(new_n401), .B2(new_n386), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n387), .A2(new_n388), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n390), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT7), .B1(new_n404), .B2(G20), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT79), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n385), .C1(new_n400), .C2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n332), .B2(new_n210), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n263), .A2(KEYINPUT81), .A3(G33), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n265), .A2(KEYINPUT81), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n403), .C2(KEYINPUT3), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n386), .A2(G20), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n383), .B(new_n379), .C1(new_n413), .C2(new_n351), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT82), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n281), .B(new_n407), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT83), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n414), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT82), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT83), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n281), .A4(new_n407), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n371), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n259), .B1(G232), .B2(new_n261), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  XOR2_X1   g0229(.A(new_n429), .B(KEYINPUT84), .Z(new_n430));
  MUX2_X1   g0230(.A(G223), .B(G226), .S(G1698), .Z(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n404), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n428), .B1(new_n256), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(new_n305), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(G169), .B2(new_n433), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n427), .A2(KEYINPUT18), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n420), .A2(new_n426), .ZN(new_n437));
  INV_X1    g0237(.A(new_n371), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(G200), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n275), .B2(new_n433), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT18), .B1(new_n427), .B2(new_n435), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n427), .A2(KEYINPUT17), .A3(new_n441), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n436), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n369), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  INV_X1    g0251(.A(G250), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n320), .ZN(new_n453));
  INV_X1    g0253(.A(G244), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT4), .B1(new_n404), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n271), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g0257(.A(KEYINPUT5), .B(G41), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G257), .A3(new_n256), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n257), .A2(new_n461), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n305), .A3(new_n464), .ZN(new_n465));
  XOR2_X1   g0265(.A(G97), .B(G107), .Z(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(KEYINPUT6), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n319), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n469), .A2(new_n210), .B1(new_n225), .B2(new_n376), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n413), .A2(new_n319), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n281), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR3_X1    g0272(.A1(new_n254), .A2(KEYINPUT85), .A3(G1), .ZN(new_n473));
  OAI21_X1  g0273(.A(KEYINPUT85), .B1(new_n254), .B2(G1), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n277), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n281), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n472), .B(new_n477), .C1(G97), .C2(new_n277), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n457), .A2(new_n462), .A3(new_n464), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n341), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n465), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT86), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n299), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n483), .B2(new_n479), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n479), .A2(new_n275), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n487), .A3(KEYINPUT87), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n403), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(G238), .A2(G1698), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n454), .B2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n404), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n256), .ZN(new_n498));
  INV_X1    g0298(.A(new_n460), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n256), .A2(G250), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(new_n257), .B2(new_n499), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n299), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n503), .B1(G190), .B2(new_n502), .ZN(new_n504));
  NAND3_X1  g0304(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  INV_X1    g0306(.A(G87), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n210), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT88), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n404), .A2(new_n210), .A3(G68), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n353), .A2(new_n333), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(KEYINPUT19), .C2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n311), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n512), .A2(new_n281), .B1(new_n278), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n476), .A2(G87), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n504), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n502), .A2(G169), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n305), .B2(new_n502), .ZN(new_n518));
  XOR2_X1   g0318(.A(new_n311), .B(KEYINPUT89), .Z(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n476), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n404), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n210), .B2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n319), .A2(KEYINPUT23), .A3(G20), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n494), .A2(new_n210), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n332), .A2(G20), .A3(new_n507), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n525), .B(new_n529), .C1(KEYINPUT22), .C2(new_n530), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT24), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n281), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n277), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n278), .A2(KEYINPUT25), .A3(new_n319), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n476), .A2(G107), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G264), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n461), .A2(new_n256), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n464), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G294), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n403), .A2(new_n542), .ZN(new_n543));
  MUX2_X1   g0343(.A(G250), .B(G257), .S(G1698), .Z(new_n544));
  AOI21_X1  g0344(.A(new_n543), .B1(new_n404), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n256), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n299), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n524), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n492), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n538), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n305), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(G169), .B2(new_n547), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n277), .A2(G116), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n476), .B2(G116), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n451), .B(new_n210), .C1(G33), .C2(new_n333), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT90), .ZN(new_n561));
  XNOR2_X1  g0361(.A(new_n560), .B(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(new_n281), .C1(new_n210), .C2(G116), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  OR2_X1    g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT91), .ZN(new_n570));
  INV_X1    g0370(.A(G270), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G257), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n539), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n404), .A2(new_n573), .B1(G303), .B2(new_n332), .ZN(new_n574));
  OAI221_X1 g0374(.A(new_n464), .B1(new_n571), .B2(new_n540), .C1(new_n574), .C2(new_n256), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n568), .A2(G169), .A3(new_n570), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(G169), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT91), .B(new_n569), .C1(new_n567), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n305), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n568), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n576), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n575), .A2(new_n275), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n575), .A2(G200), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n567), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OR3_X1    g0384(.A1(new_n556), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n449), .A2(new_n552), .A3(new_n585), .ZN(G372));
  OAI21_X1  g0386(.A(new_n364), .B1(new_n367), .B2(new_n327), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(new_n444), .A3(new_n446), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n436), .A2(new_n445), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n303), .A2(new_n300), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n307), .B2(new_n306), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n556), .A2(new_n581), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n492), .A3(new_n551), .ZN(new_n594));
  INV_X1    g0394(.A(new_n523), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT26), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n524), .B2(new_n481), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n482), .A2(KEYINPUT26), .A3(new_n523), .A4(new_n516), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n592), .B1(new_n449), .B2(new_n600), .ZN(G369));
  NAND3_X1  g0401(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n602), .A2(KEYINPUT27), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(KEYINPUT27), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(G213), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G343), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n567), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n581), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n609), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n576), .A2(new_n611), .A3(new_n578), .A4(new_n580), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n584), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G330), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n538), .A2(new_n607), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n556), .A2(new_n608), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n618), .A2(new_n581), .A3(new_n608), .A4(new_n619), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n619), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n625), .ZN(G399));
  INV_X1    g0426(.A(new_n213), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(G41), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n506), .A2(new_n507), .A3(new_n493), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(G1), .A3(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n221), .B2(new_n629), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT28), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n607), .B1(new_n594), .B2(new_n599), .ZN(new_n635));
  XNOR2_X1  g0435(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT92), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT29), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  OR3_X1    g0441(.A1(new_n552), .A2(new_n585), .A3(new_n607), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n579), .A2(new_n463), .A3(new_n502), .A4(new_n547), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT30), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n547), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n502), .A2(G179), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n479), .A4(new_n575), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n607), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT31), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n642), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n637), .A2(new_n641), .B1(new_n653), .B2(G330), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n634), .B1(new_n654), .B2(G1), .ZN(G364));
  INV_X1    g0455(.A(G330), .ZN(new_n656));
  AOI211_X1 g0456(.A(new_n656), .B(new_n584), .C1(new_n610), .C2(new_n612), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n216), .A2(G20), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n209), .B1(new_n658), .B2(G45), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n628), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(G330), .B1(new_n613), .B2(new_n614), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n613), .A2(new_n614), .ZN(new_n665));
  NOR2_X1   g0465(.A1(G13), .A2(G33), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n213), .A2(new_n266), .ZN(new_n670));
  INV_X1    g0470(.A(G355), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n670), .A2(new_n671), .B1(G116), .B2(new_n213), .ZN(new_n672));
  AOI211_X1 g0472(.A(new_n404), .B(new_n627), .C1(new_n459), .C2(new_n222), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n252), .A2(G45), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n217), .B1(new_n210), .B2(G169), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT93), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT93), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n668), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n661), .B1(new_n675), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n210), .A2(G179), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(G190), .A3(G200), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n507), .ZN(new_n685));
  NOR2_X1   g0485(.A1(G190), .A2(G200), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n377), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(KEYINPUT32), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n275), .A2(G179), .A3(G200), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n210), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n685), .B(new_n690), .C1(G97), .C2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n210), .A2(new_n305), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n686), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n266), .B1(new_n696), .B2(new_n225), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(G190), .A3(new_n299), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n697), .B1(new_n287), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(G200), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G190), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n683), .A2(new_n275), .A3(G200), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n702), .A2(G68), .B1(new_n704), .B2(G107), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n701), .A2(new_n275), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n689), .A2(KEYINPUT32), .B1(new_n706), .B2(G50), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n694), .A2(new_n700), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n687), .A2(KEYINPUT94), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n687), .A2(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G329), .ZN(new_n713));
  INV_X1    g0513(.A(G283), .ZN(new_n714));
  INV_X1    g0514(.A(G303), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n714), .A2(new_n703), .B1(new_n684), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT33), .B(G317), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n716), .B1(new_n702), .B2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G311), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n332), .B1(new_n696), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(G322), .B2(new_n699), .ZN(new_n721));
  AOI22_X1  g0521(.A1(G294), .A2(new_n693), .B1(new_n706), .B2(G326), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n713), .A2(new_n718), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n708), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n682), .B1(new_n724), .B2(new_n679), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n662), .A2(new_n664), .B1(new_n669), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(G396));
  NOR2_X1   g0527(.A1(new_n327), .A2(new_n607), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n316), .A2(new_n607), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n325), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n730), .B2(new_n327), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n635), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n653), .A2(G330), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n661), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n679), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n667), .ZN(new_n738));
  INV_X1    g0538(.A(new_n702), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n739), .A2(new_n714), .B1(new_n703), .B2(new_n507), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n332), .B1(new_n696), .B2(new_n493), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(G294), .B2(new_n699), .ZN(new_n742));
  INV_X1    g0542(.A(new_n684), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n693), .A2(G97), .B1(new_n743), .B2(G107), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n742), .B(new_n744), .C1(new_n719), .C2(new_n711), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n740), .B(new_n745), .C1(G303), .C2(new_n706), .ZN(new_n746));
  XOR2_X1   g0546(.A(KEYINPUT95), .B(G143), .Z(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n696), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n699), .A2(new_n748), .B1(new_n749), .B2(G159), .ZN(new_n750));
  INV_X1    g0550(.A(G150), .ZN(new_n751));
  INV_X1    g0551(.A(G137), .ZN(new_n752));
  INV_X1    g0552(.A(new_n706), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n750), .B1(new_n739), .B2(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT34), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n693), .A2(new_n287), .B1(new_n743), .B2(G50), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n398), .B1(G68), .B2(new_n704), .ZN(new_n758));
  INV_X1    g0558(.A(G132), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n757), .B(new_n758), .C1(new_n711), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n754), .A2(new_n755), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n746), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n661), .B1(G77), .B2(new_n738), .C1(new_n763), .C2(new_n737), .ZN(new_n764));
  INV_X1    g0564(.A(new_n731), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n666), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n736), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(G384));
  AOI211_X1 g0569(.A(new_n371), .B(new_n440), .C1(new_n420), .C2(new_n426), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n385), .B1(new_n400), .B2(new_n406), .ZN(new_n771));
  AOI21_X1  g0571(.A(KEYINPUT16), .B1(new_n771), .B2(KEYINPUT97), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n393), .B1(new_n392), .B2(new_n399), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n402), .A2(KEYINPUT79), .A3(new_n405), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n384), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT97), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n285), .B1(new_n772), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT98), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n407), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n416), .B1(new_n775), .B2(new_n776), .ZN(new_n781));
  AOI211_X1 g0581(.A(KEYINPUT97), .B(new_n384), .C1(new_n773), .C2(new_n774), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n779), .B(new_n281), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n438), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n435), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n770), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT99), .ZN(new_n788));
  INV_X1    g0588(.A(new_n407), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n281), .B1(new_n781), .B2(new_n782), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(KEYINPUT98), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n371), .B1(new_n791), .B2(new_n783), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n788), .B1(new_n792), .B2(new_n605), .ZN(new_n793));
  INV_X1    g0593(.A(new_n605), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n785), .A2(KEYINPUT99), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n787), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(KEYINPUT37), .ZN(new_n797));
  INV_X1    g0597(.A(new_n427), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n786), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n794), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT37), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n442), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT38), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n793), .A2(new_n795), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n447), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n803), .A2(KEYINPUT100), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n805), .A2(new_n447), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(KEYINPUT38), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n442), .B1(new_n427), .B2(new_n435), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n427), .A2(new_n605), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n811), .A2(KEYINPUT37), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n796), .B2(KEYINPUT37), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n808), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n447), .A2(new_n812), .ZN(new_n816));
  OAI21_X1  g0616(.A(KEYINPUT37), .B1(new_n811), .B2(new_n812), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n802), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n804), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n807), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n363), .A2(new_n607), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n364), .A2(new_n368), .A3(new_n822), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n363), .B(new_n607), .C1(new_n350), .C2(new_n367), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND4_X1   g0625(.A1(KEYINPUT40), .A2(new_n825), .A3(new_n653), .A4(new_n731), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT102), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n821), .A2(KEYINPUT102), .A3(new_n826), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n803), .A2(new_n806), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n805), .A2(new_n447), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n804), .B1(new_n814), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n825), .A2(new_n653), .A3(new_n731), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT40), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT103), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n449), .B1(new_n642), .B2(new_n652), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n656), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n841), .B2(new_n842), .ZN(new_n844));
  INV_X1    g0644(.A(new_n364), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n608), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT38), .B1(new_n803), .B2(new_n809), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n810), .A2(new_n814), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT39), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT39), .B1(new_n819), .B2(new_n804), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n807), .A2(new_n815), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n846), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n823), .A2(new_n824), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n728), .B1(new_n635), .B2(new_n731), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n835), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n589), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n605), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n641), .B1(new_n635), .B2(new_n636), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n449), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT101), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n861), .A2(new_n449), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n592), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n860), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n844), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n844), .A2(new_n870), .ZN(new_n874));
  OAI21_X1  g0674(.A(G1), .B1(new_n216), .B2(G20), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n469), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n219), .A4(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n880), .B(KEYINPUT36), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n222), .A2(G77), .A3(new_n374), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(G50), .B2(new_n351), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(G1), .A3(new_n216), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n876), .A2(new_n881), .A3(new_n884), .ZN(G367));
  AOI21_X1  g0685(.A(new_n608), .B1(new_n514), .B2(new_n515), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n524), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n595), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT43), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n889), .A2(KEYINPUT43), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n478), .A2(new_n607), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n492), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n492), .A2(KEYINPUT105), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n482), .A2(new_n607), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT106), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n623), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n894), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n907), .A2(KEYINPUT42), .A3(new_n623), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n556), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n607), .B1(new_n910), .B2(new_n481), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n892), .B(new_n893), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n911), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n906), .A2(new_n908), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n891), .A4(new_n890), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n907), .A2(new_n622), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n912), .A2(new_n915), .A3(new_n917), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n628), .B(KEYINPUT41), .Z(new_n922));
  NAND2_X1  g0722(.A1(new_n907), .A2(new_n624), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT44), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n904), .A2(KEYINPUT45), .A3(new_n625), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT45), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n907), .B2(new_n624), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n622), .B1(new_n925), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT108), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n581), .A2(new_n608), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n620), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT107), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n934), .A2(new_n623), .B1(new_n657), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n657), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n615), .A2(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n934), .A2(new_n623), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n654), .A2(new_n932), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n941), .A2(new_n861), .A3(new_n733), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT108), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n925), .A2(new_n622), .A3(new_n929), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n931), .A2(new_n942), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n922), .B1(new_n946), .B2(new_n654), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n921), .B1(new_n947), .B2(new_n660), .ZN(new_n948));
  INV_X1    g0748(.A(new_n661), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n680), .B1(new_n213), .B2(new_n513), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n627), .A2(new_n404), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n242), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n704), .A2(G77), .ZN(new_n953));
  INV_X1    g0753(.A(new_n287), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n953), .B1(new_n954), .B2(new_n684), .C1(new_n739), .C2(new_n377), .ZN(new_n955));
  INV_X1    g0755(.A(new_n687), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n332), .B1(new_n956), .B2(G137), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n202), .B2(new_n696), .C1(new_n751), .C2(new_n698), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n753), .A2(new_n747), .B1(new_n351), .B2(new_n692), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n704), .A2(G97), .ZN(new_n961));
  INV_X1    g0761(.A(G317), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n961), .B(new_n398), .C1(new_n962), .C2(new_n687), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n963), .B(KEYINPUT109), .Z(new_n964));
  AOI22_X1  g0764(.A1(new_n699), .A2(G303), .B1(new_n749), .B2(G283), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n319), .B2(new_n692), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n739), .A2(new_n542), .B1(new_n753), .B2(new_n719), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n684), .A2(new_n493), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT46), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n960), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT47), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n737), .B1(new_n971), .B2(KEYINPUT47), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n949), .B(new_n952), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n668), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n889), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT110), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n948), .A2(new_n978), .ZN(G387));
  NAND2_X1  g0779(.A1(new_n313), .A2(new_n202), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT112), .Z(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT50), .ZN(new_n983));
  AOI211_X1 g0783(.A(G45), .B(new_n630), .C1(G68), .C2(G77), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT111), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n951), .C1(new_n459), .C2(new_n239), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(G107), .B2(new_n213), .C1(new_n631), .C2(new_n670), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n949), .B1(new_n988), .B2(new_n680), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n699), .A2(G50), .B1(new_n749), .B2(G68), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n751), .B2(new_n687), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n288), .B2(new_n702), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n706), .A2(G159), .B1(new_n743), .B2(G77), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n992), .A2(new_n404), .A3(new_n961), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n520), .A2(new_n692), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n699), .A2(G317), .B1(new_n749), .B2(G303), .ZN(new_n997));
  INV_X1    g0797(.A(G322), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n739), .B2(new_n719), .C1(new_n998), .C2(new_n753), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n693), .A2(G283), .B1(new_n743), .B2(G294), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT49), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n703), .A2(new_n493), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n404), .B(new_n1006), .C1(G326), .C2(new_n956), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n996), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n989), .B1(new_n737), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n620), .B2(new_n668), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n941), .B2(new_n660), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n944), .A2(new_n942), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(KEYINPUT113), .A3(new_n628), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n654), .B2(new_n941), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT113), .B1(new_n1012), .B2(new_n628), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(G393));
  INV_X1    g0816(.A(new_n945), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1012), .B1(new_n1017), .B2(new_n930), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n946), .A2(new_n1018), .A3(new_n628), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1017), .A2(new_n930), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n907), .A2(new_n668), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n313), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n404), .B1(new_n687), .B2(new_n747), .C1(new_n1022), .C2(new_n696), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n739), .A2(new_n202), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n351), .A2(new_n684), .B1(new_n703), .B2(new_n507), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n692), .A2(new_n225), .ZN(new_n1026));
  NOR4_X1   g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n753), .A2(new_n751), .B1(new_n377), .B2(new_n698), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n753), .A2(new_n962), .B1(new_n719), .B2(new_n698), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n739), .A2(new_n715), .B1(new_n493), .B2(new_n692), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n332), .B1(new_n687), .B2(new_n998), .C1(new_n542), .C2(new_n696), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n319), .A2(new_n703), .B1(new_n684), .B2(new_n714), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1027), .A2(new_n1029), .B1(new_n1031), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1036), .A2(new_n737), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n248), .A2(new_n951), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n681), .B1(G97), .B2(new_n627), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n949), .B(new_n1037), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1020), .A2(new_n660), .B1(new_n1021), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1019), .A2(new_n1041), .ZN(G390));
  OAI21_X1  g0842(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n849), .A2(new_n851), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1043), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n821), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n825), .A2(new_n653), .A3(G330), .A4(new_n731), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1044), .A2(new_n1048), .A3(new_n1046), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(new_n660), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n849), .A2(new_n666), .A3(new_n851), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n661), .B1(new_n738), .B2(new_n288), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n332), .B1(new_n698), .B2(new_n493), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(G97), .B2(new_n749), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n685), .B1(G68), .B2(new_n704), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n542), .C2(new_n711), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1026), .B1(G107), .B2(new_n702), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n714), .B2(new_n753), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT54), .B(G143), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n266), .B1(new_n696), .B2(new_n1063), .C1(new_n759), .C2(new_n698), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n712), .B2(G125), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n684), .A2(new_n751), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT53), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G128), .A2(new_n706), .B1(new_n702), .B2(G137), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n693), .A2(G159), .B1(new_n704), .B2(G50), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1062), .B1(KEYINPUT115), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT115), .B2(new_n1070), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1055), .B1(new_n1072), .B2(new_n679), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1054), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n863), .A2(G330), .A3(new_n653), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n592), .B(new_n1075), .C1(new_n864), .C2(new_n866), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n552), .A2(new_n585), .A3(new_n607), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n652), .ZN(new_n1078));
  OAI211_X1 g0878(.A(G330), .B(new_n731), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n853), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1048), .A2(new_n1080), .A3(new_n854), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n854), .B1(new_n1048), .B2(new_n1080), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1050), .A2(new_n1051), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT114), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n628), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1052), .B2(new_n1084), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1086), .B1(new_n1085), .B2(new_n628), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1053), .B(new_n1074), .C1(new_n1088), .C2(new_n1089), .ZN(G378));
  OAI21_X1  g0890(.A(new_n661), .B1(new_n738), .B2(G50), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n692), .A2(new_n351), .B1(new_n698), .B2(new_n319), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n702), .A2(G97), .B1(new_n704), .B2(new_n287), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n493), .B2(new_n753), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1092), .B(new_n1094), .C1(G283), .C2(new_n712), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n398), .A2(new_n255), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G77), .B2(new_n743), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT116), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1095), .B(new_n1098), .C1(new_n520), .C2(new_n696), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT58), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1096), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n706), .A2(G125), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n739), .B2(new_n759), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n699), .A2(G128), .B1(new_n749), .B2(G137), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n684), .B2(new_n1063), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1105), .B(new_n1107), .C1(G150), .C2(new_n693), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n704), .A2(G159), .ZN(new_n1112));
  AOI211_X1 g0912(.A(G33), .B(G41), .C1(new_n956), .C2(G124), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n1103), .B1(new_n1100), .B2(new_n1099), .C1(new_n1110), .C2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1091), .B1(new_n1115), .B2(new_n679), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n591), .A2(new_n308), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n294), .A2(new_n605), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT55), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1117), .B(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1121));
  XNOR2_X1  g0921(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1116), .B1(new_n1122), .B2(new_n667), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT118), .B1(new_n852), .B2(new_n859), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n846), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n807), .A2(new_n815), .A3(new_n850), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT39), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n832), .B2(new_n834), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1126), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n835), .A2(new_n855), .B1(new_n857), .B2(new_n605), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n656), .B1(new_n837), .B2(new_n838), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n821), .A2(KEYINPUT102), .A3(new_n826), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT102), .B1(new_n821), .B2(new_n826), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1122), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1122), .B1(new_n831), .B2(new_n1135), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1134), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1122), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n860), .A3(new_n1138), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1124), .B1(new_n1146), .B2(new_n660), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT57), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1076), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1085), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n1144), .A2(new_n860), .A3(new_n1138), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n860), .B1(new_n1144), .B2(new_n1138), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT119), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1150), .B(KEYINPUT119), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n1141), .A2(new_n1145), .B1(new_n1149), .B2(new_n1085), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n628), .B1(new_n1158), .B2(KEYINPUT57), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1147), .B1(new_n1157), .B2(new_n1159), .ZN(G375));
  NOR2_X1   g0960(.A1(new_n1083), .A2(new_n659), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n853), .A2(new_n666), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n661), .B1(new_n738), .B2(G68), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n711), .A2(new_n715), .B1(new_n333), .B2(new_n684), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT121), .Z(new_n1165));
  OAI221_X1 g0965(.A(new_n332), .B1(new_n696), .B2(new_n319), .C1(new_n714), .C2(new_n698), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n953), .B1(new_n739), .B2(new_n493), .C1(new_n542), .C2(new_n753), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n995), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n712), .A2(G128), .B1(G159), .B2(new_n743), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT122), .Z(new_n1170));
  OAI221_X1 g0970(.A(new_n404), .B1(new_n752), .B2(new_n698), .C1(new_n751), .C2(new_n696), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G50), .A2(new_n693), .B1(new_n706), .B2(G132), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n954), .B2(new_n703), .C1(new_n739), .C2(new_n1063), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1168), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1163), .B1(new_n1175), .B2(new_n679), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1161), .B1(new_n1162), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1084), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n922), .B(KEYINPUT120), .Z(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1076), .A2(new_n1083), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1177), .B1(new_n1180), .B2(new_n1181), .ZN(G381));
  OR4_X1    g0982(.A1(G384), .A2(G387), .A3(G390), .A4(G381), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n726), .B(new_n1011), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1184));
  OR4_X1    g0984(.A1(G378), .A2(G375), .A3(new_n1183), .A4(new_n1184), .ZN(G407));
  INV_X1    g0985(.A(G378), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n606), .A2(G213), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(G407), .B(G213), .C1(G375), .C2(new_n1189), .ZN(G409));
  INV_X1    g0990(.A(KEYINPUT63), .ZN(new_n1191));
  OAI211_X1 g0991(.A(G378), .B(new_n1147), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1158), .A2(new_n1179), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n660), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1123), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1186), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1187), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1181), .B1(new_n1178), .B2(KEYINPUT60), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1076), .A2(KEYINPUT60), .A3(new_n1083), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n628), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1177), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n768), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G384), .B(new_n1177), .C1(new_n1199), .C2(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1191), .B1(new_n1198), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1207), .A3(new_n1204), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1188), .A2(G2897), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1205), .A2(KEYINPUT123), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT61), .B1(new_n1198), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(G393), .A2(G396), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1184), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G390), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n919), .A2(new_n920), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n922), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1017), .A2(new_n1012), .A3(new_n930), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n654), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1221), .B1(new_n1225), .B2(new_n659), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1220), .B(KEYINPUT124), .C1(new_n1226), .C2(new_n977), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n948), .A2(new_n978), .A3(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT124), .B1(G387), .B2(new_n1220), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1219), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(KEYINPUT125), .B(new_n1219), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT126), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G387), .B2(new_n1220), .ZN(new_n1236));
  AOI211_X1 g1036(.A(KEYINPUT126), .B(G390), .C1(new_n948), .C2(new_n978), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1228), .A2(new_n1218), .ZN(new_n1238));
  OR3_X1    g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1233), .A2(new_n1234), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1188), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1205), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1206), .A2(new_n1216), .A3(new_n1240), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1241), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1241), .B2(new_n1214), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1246), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1244), .B1(new_n1250), .B2(new_n1240), .ZN(G405));
  NAND3_X1  g1051(.A1(new_n1240), .A2(KEYINPUT127), .A3(new_n1205), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1205), .A2(KEYINPUT127), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1233), .A2(new_n1234), .A3(new_n1239), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G375), .A2(new_n1186), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n1192), .C1(KEYINPUT127), .C2(new_n1205), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1255), .B(new_n1257), .ZN(G402));
endmodule


