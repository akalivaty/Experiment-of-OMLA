//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n208), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n202), .B2(new_n226), .C1(new_n203), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n210), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n218), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT64), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n237), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G274), .ZN(new_n252));
  AND2_X1   g0052(.A1(G1), .A2(G13), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n255), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT68), .B1(new_n255), .B2(new_n257), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n253), .A2(new_n254), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n260), .B1(G238), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n265), .A2(new_n266), .A3(KEYINPUT69), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT69), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G226), .A2(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n226), .B2(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n261), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT77), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT77), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n282), .B(new_n261), .C1(new_n277), .C2(new_n278), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n264), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT13), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(new_n264), .C1(new_n281), .C2(new_n283), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g0088(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G169), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT80), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n292), .B1(new_n285), .B2(new_n287), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT80), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n294), .A3(new_n289), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT14), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  OAI22_X1  g0098(.A1(new_n293), .A2(new_n297), .B1(new_n288), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT74), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n305), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n302), .B1(new_n307), .B2(G68), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT12), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(new_n311), .A3(G20), .A4(new_n203), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n216), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT71), .B1(new_n270), .B2(G20), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n208), .A3(G33), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n319), .A3(G77), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n316), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT11), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n313), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n315), .B1(new_n304), .B2(new_n306), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n207), .A2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G68), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n323), .B2(KEYINPUT11), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n301), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n288), .A2(G200), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n285), .A2(G190), .A3(new_n287), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n330), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n208), .B1(new_n267), .B2(new_n273), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n265), .A2(new_n266), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n203), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n202), .A2(new_n203), .ZN(new_n344));
  NOR2_X1   g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n321), .A2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(KEYINPUT81), .B(new_n337), .C1(new_n343), .C2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT69), .B1(new_n265), .B2(new_n266), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n271), .A2(new_n268), .A3(new_n272), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n342), .B1(new_n353), .B2(KEYINPUT7), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(G68), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n350), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  INV_X1    g0156(.A(new_n342), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n341), .B2(new_n208), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n348), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n361), .A2(new_n315), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n349), .A2(new_n356), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT8), .B(G58), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n327), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n316), .A2(new_n303), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n303), .B2(new_n365), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n363), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n271), .A2(new_n272), .ZN(new_n372));
  INV_X1    g0172(.A(G223), .ZN(new_n373));
  INV_X1    g0173(.A(G1698), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n372), .B(new_n375), .C1(G226), .C2(new_n374), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n270), .A2(new_n222), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n280), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n262), .A2(new_n226), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n255), .A2(new_n257), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT68), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n255), .A2(KEYINPUT68), .A3(new_n257), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT82), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n379), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n258), .A2(new_n259), .B1(new_n226), .B2(new_n262), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(KEYINPUT82), .ZN(new_n389));
  OAI21_X1  g0189(.A(G169), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n386), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(KEYINPUT82), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(G179), .A4(new_n379), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n370), .A2(new_n371), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n371), .B1(new_n370), .B2(new_n394), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G200), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n387), .B2(new_n389), .ZN(new_n399));
  INV_X1    g0199(.A(G190), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n391), .A2(new_n392), .A3(new_n400), .A4(new_n379), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n363), .A2(new_n402), .A3(new_n369), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n374), .A2(G222), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n274), .B(new_n406), .C1(new_n373), .C2(new_n374), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n280), .C1(G77), .C2(new_n274), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n260), .B1(G226), .B2(new_n263), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT70), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n321), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n317), .A2(new_n319), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n364), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n315), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n327), .A2(G50), .ZN(new_n421));
  OAI221_X1 g0221(.A(new_n420), .B1(G50), .B2(new_n303), .C1(new_n367), .C2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n414), .A2(new_n298), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n416), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n412), .A2(G200), .A3(new_n413), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n422), .B(KEYINPUT9), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n415), .C2(new_n400), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT10), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT76), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n430), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n321), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n434), .A2(KEYINPUT73), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(KEYINPUT73), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n365), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT15), .B(G87), .ZN(new_n438));
  OAI221_X1 g0238(.A(new_n437), .B1(new_n208), .B2(new_n220), .C1(new_n418), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n315), .ZN(new_n440));
  INV_X1    g0240(.A(new_n307), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n220), .B1(new_n207), .B2(G20), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n441), .A2(new_n220), .B1(new_n326), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n227), .A2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G232), .B2(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n274), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G107), .B2(new_n274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT72), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT72), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n448), .B(new_n451), .C1(G107), .C2(new_n274), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(new_n280), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n260), .B1(G244), .B2(new_n263), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n445), .B1(new_n455), .B2(new_n292), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT75), .B1(new_n455), .B2(G179), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n453), .A2(new_n458), .A3(new_n298), .A4(new_n454), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n444), .B1(new_n455), .B2(G200), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n400), .B2(new_n455), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n336), .A2(new_n405), .A3(new_n433), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G257), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n374), .ZN(new_n466));
  OAI221_X1 g0266(.A(new_n466), .B1(G264), .B2(new_n374), .C1(new_n265), .C2(new_n266), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G303), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n351), .B2(new_n352), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n280), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G41), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n207), .B(G45), .C1(new_n472), .C2(KEYINPUT5), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n255), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n261), .B(G270), .C1(new_n473), .C2(new_n474), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n471), .A2(G179), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G116), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n207), .B2(G33), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n307), .A2(new_n316), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n304), .A2(new_n480), .A3(new_n306), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n314), .A2(new_n216), .B1(G20), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n208), .C1(G33), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n482), .B(new_n483), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(KEYINPUT88), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT88), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n441), .A2(new_n480), .B1(new_n326), .B2(new_n481), .ZN(new_n494));
  INV_X1    g0294(.A(new_n490), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n488), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n479), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n491), .A2(KEYINPUT88), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n494), .A2(new_n496), .A3(new_n493), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT89), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n479), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n471), .A2(new_n478), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT87), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n502), .B1(new_n510), .B2(G190), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n398), .B2(new_n510), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT21), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n502), .A2(G169), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n510), .ZN(new_n515));
  INV_X1    g0315(.A(new_n510), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n292), .B1(new_n500), .B2(new_n501), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(KEYINPUT21), .A3(new_n517), .ZN(new_n518));
  AND4_X1   g0318(.A1(new_n505), .A2(new_n512), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n351), .A2(new_n352), .A3(G250), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n374), .B1(new_n520), .B2(KEYINPUT4), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT4), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n522), .A2(new_n221), .A3(G1698), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n351), .A2(new_n352), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n341), .B2(new_n221), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(new_n485), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n280), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n476), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n475), .A2(new_n280), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n292), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n303), .A2(G97), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n367), .B1(new_n207), .B2(G33), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G97), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT6), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n536), .A2(new_n486), .A3(G107), .ZN(new_n537));
  XNOR2_X1  g0337(.A(G97), .B(G107), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n539), .A2(new_n208), .B1(new_n220), .B2(new_n434), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n354), .B2(G107), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n535), .B1(new_n541), .B2(new_n316), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n527), .A2(new_n298), .A3(new_n530), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT84), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT84), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n532), .A2(new_n542), .A3(new_n546), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n527), .A2(new_n550), .A3(new_n530), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(G200), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n531), .A2(new_n400), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n542), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n548), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n418), .B2(new_n486), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n208), .B1(new_n278), .B2(new_n557), .ZN(new_n559));
  INV_X1    g0359(.A(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n222), .A2(new_n486), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT85), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n372), .A2(new_n208), .A3(G68), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT85), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n565), .A3(new_n561), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n558), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n315), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n441), .A2(new_n438), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n534), .A2(G87), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n227), .A2(new_n374), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n221), .A2(G1698), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n572), .B(new_n573), .C1(new_n265), .C2(new_n266), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G33), .A2(G116), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n261), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n207), .A2(new_n252), .A3(G45), .ZN(new_n577));
  INV_X1    g0377(.A(G45), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n223), .B1(new_n578), .B2(G1), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n261), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G190), .ZN(new_n583));
  OAI21_X1  g0383(.A(G200), .B1(new_n576), .B2(new_n581), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n571), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n574), .A2(new_n575), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n298), .B(new_n580), .C1(new_n587), .C2(new_n261), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n292), .B1(new_n576), .B2(new_n581), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n567), .A2(new_n315), .B1(new_n441), .B2(new_n438), .ZN(new_n591));
  INV_X1    g0391(.A(new_n438), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n534), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n556), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(new_n590), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n591), .A2(new_n570), .A3(new_n584), .A4(new_n583), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(KEYINPUT86), .A3(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n534), .A2(G107), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n303), .A2(G107), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT25), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT22), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n351), .A2(new_n352), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n208), .A2(G87), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n606), .A2(new_n222), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n208), .C1(new_n266), .C2(new_n265), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT23), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n208), .B2(G107), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n560), .A2(KEYINPUT23), .A3(G20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT24), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n609), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n605), .B1(new_n622), .B2(new_n315), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n261), .B(G264), .C1(new_n473), .C2(new_n474), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n223), .A2(new_n374), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n465), .A2(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n627), .C1(new_n265), .C2(new_n266), .ZN(new_n628));
  NAND2_X1  g0428(.A1(G33), .A2(G294), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n261), .B1(new_n630), .B2(KEYINPUT90), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT90), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n628), .A2(new_n632), .A3(new_n629), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n625), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n400), .A3(new_n476), .ZN(new_n635));
  AOI211_X1 g0435(.A(new_n625), .B(new_n528), .C1(new_n631), .C2(new_n633), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(G200), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n476), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n292), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n636), .A2(new_n298), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n316), .B1(new_n619), .B2(new_n621), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n605), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n601), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n464), .A2(new_n519), .A3(new_n555), .A4(new_n645), .ZN(G372));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n598), .A2(new_n599), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n544), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n601), .A2(new_n548), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n647), .ZN(new_n651));
  INV_X1    g0451(.A(new_n548), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n505), .A2(new_n518), .A3(new_n515), .A4(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n554), .A2(new_n552), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n586), .B1(new_n623), .B2(new_n637), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n651), .A2(new_n598), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n464), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n424), .ZN(new_n659));
  INV_X1    g0459(.A(new_n335), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(new_n460), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(new_n331), .B2(new_n301), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n363), .A2(new_n402), .A3(new_n369), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n397), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n431), .A2(new_n432), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n659), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n658), .A2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n310), .A2(new_n208), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n670), .B(KEYINPUT91), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT27), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(G213), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G343), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n644), .B1(new_n623), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n679));
  INV_X1    g0479(.A(new_n643), .ZN(new_n680));
  INV_X1    g0480(.A(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n681), .A2(new_n502), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n519), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n518), .A2(new_n515), .ZN(new_n687));
  INV_X1    g0487(.A(new_n505), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n689), .B2(new_n685), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT92), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n690), .A2(new_n691), .A3(G330), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n690), .B2(G330), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n684), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n679), .A2(new_n683), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n677), .B1(new_n687), .B2(new_n688), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n680), .A2(new_n677), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n694), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n211), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n207), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n561), .A2(G116), .ZN(new_n707));
  INV_X1    g0507(.A(new_n704), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n706), .A2(new_n707), .B1(new_n214), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT29), .B1(new_n657), .B2(new_n677), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n595), .A2(new_n600), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n545), .B2(new_n547), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT96), .B1(new_n713), .B2(KEYINPUT26), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n650), .A2(new_n715), .A3(new_n647), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n648), .A2(new_n544), .A3(new_n647), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n505), .A2(new_n518), .A3(new_n515), .A4(new_n643), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n654), .A2(new_n545), .A3(new_n655), .A4(new_n547), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n598), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n681), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n711), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT94), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n479), .A2(new_n582), .A3(new_n634), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n531), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n725), .B(new_n729), .C1(new_n726), .C2(new_n531), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n636), .A2(G179), .A3(new_n582), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n516), .A2(new_n731), .A3(new_n531), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n519), .A2(new_n555), .A3(new_n645), .A4(new_n677), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n734), .A2(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT31), .B1(new_n733), .B2(new_n681), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n735), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n724), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n710), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n692), .A2(new_n693), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n309), .A2(new_n578), .A3(G20), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT97), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n706), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n745), .B(new_n749), .C1(G330), .C2(new_n690), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n274), .A2(G355), .A3(new_n211), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G116), .B2(new_n211), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n247), .A2(new_n578), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n703), .A2(new_n372), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n578), .B2(new_n215), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n752), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n216), .B1(G20), .B2(new_n292), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n748), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n208), .A2(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(G179), .A3(G200), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n398), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n771), .A2(G329), .B1(G283), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT101), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n766), .A2(new_n298), .A3(new_n398), .ZN(new_n777));
  INV_X1    g0577(.A(G317), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n778), .A2(KEYINPUT33), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n208), .A2(new_n298), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(new_n400), .A3(new_n398), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n772), .A2(G20), .A3(G190), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G311), .A2(new_n784), .B1(new_n786), .B2(G303), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n782), .A2(G190), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n398), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G326), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n790), .A2(new_n791), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n298), .A2(new_n398), .A3(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G294), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n607), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n776), .A2(new_n781), .A3(new_n787), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n771), .A2(G159), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n803), .A2(KEYINPUT32), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n607), .B1(G87), .B2(new_n786), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(KEYINPUT32), .B1(KEYINPUT99), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n773), .A2(new_n560), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G77), .B2(new_n784), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n202), .B2(new_n790), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n807), .B(new_n810), .C1(G50), .C2(new_n792), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n777), .A2(G68), .B1(new_n797), .B2(G97), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT100), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n804), .A2(new_n806), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n802), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n764), .B1(new_n815), .B2(new_n761), .ZN(new_n816));
  INV_X1    g0616(.A(new_n760), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n690), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n750), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(G396));
  NOR2_X1   g0620(.A1(new_n677), .A2(new_n445), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n460), .A2(new_n462), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n456), .A2(new_n457), .A3(new_n459), .A4(new_n821), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n649), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n713), .B2(KEYINPUT26), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n677), .C1(new_n827), .C2(new_n721), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT103), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n657), .A2(new_n830), .A3(new_n677), .A4(new_n825), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n681), .B1(new_n722), .B2(new_n651), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n825), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n741), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n748), .B1(new_n834), .B2(new_n741), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n761), .A2(new_n758), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n748), .B1(G77), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G150), .A2(new_n777), .B1(new_n784), .B2(G159), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n789), .A2(G143), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n841), .B(new_n842), .C1(new_n843), .C2(new_n793), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT34), .ZN(new_n845));
  OR2_X1    g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n771), .A2(G132), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n785), .A2(new_n201), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n372), .B1(new_n773), .B2(new_n203), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(G58), .C2(new_n797), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n771), .A2(G311), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n274), .B1(G97), .B2(new_n797), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G294), .A2(new_n789), .B1(new_n792), .B2(G303), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n783), .A2(new_n480), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n785), .A2(new_n560), .B1(new_n773), .B2(new_n222), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(G283), .C2(new_n777), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n840), .B1(new_n860), .B2(new_n761), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n825), .B2(new_n759), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT102), .Z(new_n863));
  NOR2_X1   g0663(.A1(new_n838), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  INV_X1    g0665(.A(new_n539), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT35), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT35), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n867), .A2(G116), .A3(new_n217), .A4(new_n868), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI211_X1 g0670(.A(new_n215), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n201), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n207), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n301), .A2(new_n331), .A3(new_n677), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n361), .A2(new_n315), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT16), .B1(new_n359), .B2(new_n360), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n369), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n394), .B2(new_n676), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n877), .B1(new_n881), .B2(new_n403), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n370), .A2(new_n394), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n403), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n337), .B1(new_n343), .B2(new_n348), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n878), .B1(new_n885), .B2(new_n350), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n368), .B1(new_n886), .B2(new_n349), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n877), .B1(new_n887), .B2(new_n675), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT104), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n363), .A2(new_n369), .B1(new_n390), .B2(new_n393), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n663), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT104), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT37), .B1(new_n370), .B2(new_n676), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n882), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n880), .A2(new_n676), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n397), .B2(new_n404), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n876), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n900), .B(new_n876), .C1(new_n895), .C2(new_n897), .ZN(new_n901));
  INV_X1    g0701(.A(new_n897), .ZN(new_n902));
  NOR3_X1   g0702(.A1(new_n884), .A2(new_n888), .A3(KEYINPUT104), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n902), .B(KEYINPUT38), .C1(new_n905), .C2(new_n882), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n901), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT39), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n370), .A2(new_n676), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n891), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT37), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n903), .B2(new_n904), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n909), .B1(new_n397), .B2(new_n404), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n889), .A2(new_n894), .B1(new_n910), .B2(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n876), .B1(new_n917), .B2(new_n913), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n916), .A2(new_n920), .A3(new_n921), .A4(new_n906), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n875), .B1(new_n908), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n677), .A2(new_n330), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n299), .B1(new_n291), .B2(new_n295), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n335), .B(new_n925), .C1(new_n926), .C2(new_n330), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n301), .A2(new_n924), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n460), .A2(new_n681), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n832), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n907), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n675), .B1(new_n395), .B2(new_n396), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n464), .A2(new_n724), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n668), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G330), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n927), .A2(new_n928), .ZN(new_n941));
  INV_X1    g0741(.A(new_n825), .ZN(new_n942));
  INV_X1    g0742(.A(new_n734), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n738), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n942), .B1(new_n944), .B2(new_n736), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n907), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT40), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n916), .A2(new_n920), .A3(new_n906), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n941), .A2(new_n945), .A3(KEYINPUT40), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n948), .A2(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n944), .A2(new_n736), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n464), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n940), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n952), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n939), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(G1), .B1(new_n309), .B2(G20), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n939), .A2(new_n956), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n874), .B1(new_n959), .B2(new_n960), .ZN(G367));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  INV_X1    g0762(.A(new_n694), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n681), .A2(new_n542), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n555), .A2(new_n964), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n544), .A2(new_n677), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n962), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n681), .A2(new_n571), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n598), .A3(new_n599), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n598), .B2(new_n969), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(new_n967), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n694), .A2(KEYINPUT108), .A3(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n968), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n972), .B1(new_n968), .B2(new_n974), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n695), .A2(new_n697), .A3(new_n967), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT107), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n967), .A2(new_n680), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n681), .B1(new_n981), .B2(new_n652), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n979), .B2(KEYINPUT42), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n980), .A2(new_n983), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n977), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n704), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(KEYINPUT110), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n698), .B1(new_n684), .B2(new_n697), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n745), .B(new_n988), .Z(new_n989));
  AOI21_X1  g0789(.A(new_n987), .B1(new_n989), .B2(new_n743), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n987), .A3(new_n743), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n700), .B2(new_n973), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n997));
  NAND3_X1  g0797(.A1(new_n700), .A2(new_n973), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n997), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n701), .B2(new_n967), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n996), .A2(new_n694), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n963), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n991), .A2(new_n992), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n986), .B1(new_n1004), .B2(new_n743), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n747), .A2(new_n207), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n985), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n762), .B1(new_n211), .B2(new_n438), .C1(new_n242), .C2(new_n755), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT111), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n749), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1010), .B2(new_n1009), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n771), .A2(G137), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n607), .B1(new_n789), .B2(G150), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n798), .A2(new_n203), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G143), .B2(new_n792), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n773), .A2(new_n220), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n783), .A2(new_n201), .B1(new_n785), .B2(new_n202), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G159), .C2(new_n777), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n771), .A2(G317), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n785), .A2(new_n480), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(KEYINPUT46), .A2(new_n1022), .B1(new_n789), .B2(G303), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1022), .A2(KEYINPUT46), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G311), .B2(new_n792), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n341), .B1(new_n773), .B2(new_n486), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G294), .B2(new_n777), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(G283), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n798), .A2(new_n560), .B1(new_n783), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1020), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1012), .B1(new_n1033), .B2(new_n761), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n817), .B2(new_n971), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1008), .A2(new_n1035), .ZN(G387));
  AOI21_X1  g0836(.A(new_n708), .B1(new_n989), .B2(new_n743), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n743), .B2(new_n989), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n684), .A2(new_n817), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n771), .A2(G150), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n372), .B1(new_n773), .B2(new_n486), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n592), .B2(new_n797), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G50), .A2(new_n789), .B1(new_n792), .B2(G159), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n777), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1044), .A2(new_n364), .B1(new_n203), .B2(new_n783), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G77), .B2(new_n786), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n372), .B1(new_n774), .B2(G116), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n798), .A2(new_n1029), .B1(new_n799), .B2(new_n785), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G311), .A2(new_n777), .B1(new_n784), .B2(G303), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n778), .B2(new_n790), .C1(new_n791), .C2(new_n793), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT48), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT49), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1048), .B1(new_n794), .B2(new_n770), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1047), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n761), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n274), .A2(new_n211), .A3(new_n707), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(G107), .B2(new_n211), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n237), .A2(G45), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n364), .A2(G50), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT50), .ZN(new_n1064));
  AOI211_X1 g0864(.A(G45), .B(new_n707), .C1(G68), .C2(G77), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n755), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1061), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n763), .B1(new_n1067), .B2(KEYINPUT113), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(KEYINPUT113), .B2(new_n1067), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1059), .A2(new_n748), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT114), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n989), .A2(new_n1007), .B1(new_n1039), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1038), .A2(new_n1072), .ZN(G393));
  NAND2_X1  g0873(.A1(new_n1003), .A2(new_n1001), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n989), .A2(new_n743), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1004), .A2(new_n704), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT115), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1004), .A2(KEYINPUT115), .A3(new_n704), .A4(new_n1076), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1074), .A2(new_n1006), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n973), .A2(new_n760), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n762), .B1(new_n486), .B2(new_n211), .C1(new_n755), .C2(new_n250), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n748), .A2(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G150), .A2(new_n792), .B1(new_n789), .B2(G159), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT51), .Z(new_n1087));
  OAI21_X1  g0887(.A(new_n372), .B1(new_n773), .B2(new_n222), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G77), .B2(new_n797), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n771), .A2(G143), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n1044), .A2(new_n201), .B1(new_n203), .B2(new_n785), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(new_n365), .B2(new_n784), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1044), .A2(new_n469), .B1(new_n799), .B2(new_n783), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n808), .B(new_n1094), .C1(G283), .C2(new_n786), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n274), .B1(G116), .B2(new_n797), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n791), .C2(new_n770), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G311), .A2(new_n789), .B1(new_n792), .B2(G317), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1093), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1085), .B1(new_n1100), .B2(new_n761), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1082), .B1(new_n1083), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1081), .A2(new_n1102), .ZN(G390));
  NAND3_X1  g0903(.A1(new_n464), .A2(G330), .A3(new_n953), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n668), .A3(new_n937), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n929), .B1(new_n741), .B2(new_n942), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n941), .A2(new_n945), .A3(G330), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n930), .B1(new_n829), .B2(new_n831), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n742), .A2(new_n825), .A3(new_n941), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n930), .B1(new_n723), .B2(new_n825), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n945), .A2(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n929), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1105), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n875), .B1(new_n1109), .B2(new_n929), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n908), .A2(new_n1118), .A3(new_n922), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n950), .B(new_n875), .C1(new_n929), .C2(new_n1113), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n1120), .A3(new_n1112), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1117), .B(new_n1121), .C1(new_n1122), .C2(new_n1107), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1105), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1119), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1107), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1129), .A3(new_n704), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(KEYINPUT116), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n1127), .A2(new_n1128), .A3(new_n1006), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n908), .A2(new_n758), .A3(new_n922), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n748), .B1(new_n365), .B2(new_n839), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1044), .A2(new_n843), .B1(new_n783), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n773), .A2(new_n201), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G150), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n785), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT53), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1139), .B(new_n1142), .C1(new_n1143), .C2(new_n770), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n792), .A2(G128), .B1(G159), .B2(new_n797), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n607), .B1(new_n789), .B2(G132), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G116), .A2(new_n789), .B1(new_n792), .B2(G283), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1148), .B(new_n607), .C1(new_n220), .C2(new_n798), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n786), .A2(G87), .B1(new_n774), .B2(G68), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G107), .A2(new_n777), .B1(new_n784), .B2(G97), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n770), .C2(new_n799), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1144), .A2(new_n1147), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1135), .B1(new_n1153), .B2(new_n761), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1134), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1133), .A2(KEYINPUT117), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1123), .A2(new_n1129), .A3(new_n1157), .A4(new_n704), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT117), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1155), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1159), .B1(new_n1132), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1131), .A2(new_n1156), .A3(new_n1158), .A4(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT57), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n906), .B1(new_n915), .B2(KEYINPUT106), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n918), .A2(new_n919), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n951), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n895), .A2(new_n876), .A3(new_n897), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(KEYINPUT105), .B2(new_n898), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n946), .B1(new_n1168), .B2(new_n901), .ZN(new_n1169));
  OAI211_X1 g0969(.A(G330), .B(new_n1166), .C1(new_n1169), .C2(KEYINPUT40), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1171));
  OR2_X1    g0971(.A1(new_n433), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n433), .A2(new_n1171), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n676), .A2(new_n422), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1170), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n923), .A2(new_n935), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT40), .B1(new_n907), .B2(new_n947), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1177), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(G330), .A3(new_n1166), .A4(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1178), .A2(new_n1179), .A3(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1179), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1105), .B1(new_n1187), .B2(new_n1125), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1163), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1182), .B1(new_n952), .B2(G330), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n941), .A2(new_n945), .A3(KEYINPUT40), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1167), .B1(new_n919), .B2(new_n918), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(new_n916), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1180), .A2(new_n1194), .A3(new_n1177), .A4(new_n940), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n936), .B1(new_n1191), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1178), .A2(new_n1183), .A3(new_n1179), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1190), .A2(new_n1198), .A3(KEYINPUT57), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1189), .A2(new_n704), .A3(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1006), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1177), .A2(new_n758), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n748), .B1(G50), .B2(new_n839), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G50), .B1(new_n272), .B2(new_n472), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n777), .A2(G97), .B1(new_n774), .B2(G58), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n438), .B2(new_n783), .C1(new_n770), .C2(new_n1029), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n472), .B(new_n341), .C1(new_n785), .C2(new_n220), .ZN(new_n1207));
  XOR2_X1   g1007(.A(new_n1207), .B(KEYINPUT118), .Z(new_n1208));
  AOI21_X1  g1008(.A(new_n1015), .B1(G107), .B2(new_n789), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n480), .B2(new_n793), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT58), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n783), .A2(new_n843), .B1(new_n785), .B2(new_n1136), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G132), .B2(new_n777), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n789), .A2(G128), .B1(G150), .B2(new_n797), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(new_n1143), .C2(new_n793), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT59), .Z(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT119), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n771), .A2(G124), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n774), .C2(G159), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT119), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n1222), .C1(new_n1218), .C2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1213), .B1(new_n1212), .B2(new_n1211), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1203), .B1(new_n1225), .B2(new_n761), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1202), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1201), .A2(new_n1228), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1200), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(G375));
  NAND2_X1  g1031(.A1(new_n929), .A2(new_n758), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n748), .B1(G68), .B2(new_n839), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n1044), .A2(new_n480), .B1(new_n560), .B2(new_n783), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1017), .B(new_n1234), .C1(G97), .C2(new_n786), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n274), .B1(new_n592), .B2(new_n797), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G283), .A2(new_n789), .B1(new_n792), .B2(G294), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n771), .A2(G303), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n786), .A2(G159), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n1140), .B2(new_n783), .C1(new_n1044), .C2(new_n1136), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n771), .B2(G128), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n790), .A2(new_n843), .B1(new_n201), .B2(new_n798), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G132), .B2(new_n792), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n372), .B1(new_n773), .B2(new_n202), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT120), .Z(new_n1247));
  OAI21_X1  g1047(.A(new_n1239), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1233), .B1(new_n1248), .B2(new_n761), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1125), .A2(new_n1007), .B1(new_n1232), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n986), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1126), .A2(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT121), .ZN(G381));
  NAND4_X1  g1055(.A1(new_n1081), .A2(new_n1008), .A3(new_n1035), .A4(new_n1102), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1156), .A2(new_n1130), .A3(new_n1161), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1038), .A2(new_n819), .A3(new_n1072), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(G381), .A2(G384), .A3(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1257), .A2(new_n1230), .A3(new_n1258), .A4(new_n1260), .ZN(G407));
  INV_X1    g1061(.A(G213), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1262), .A2(G343), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1230), .A2(new_n1258), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(G213), .A3(new_n1264), .ZN(G409));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1105), .A2(new_n1111), .A3(KEYINPUT60), .A4(new_n1116), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1268), .A2(new_n704), .A3(new_n1126), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1250), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n864), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(KEYINPUT123), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1271), .A2(new_n1274), .A3(new_n864), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(G384), .A3(new_n1250), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1200), .A2(G378), .A3(new_n1229), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT122), .B1(new_n1201), .B2(new_n1228), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1007), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT122), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1227), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1190), .A2(new_n1198), .A3(new_n1251), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1279), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1258), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1263), .B(new_n1277), .C1(new_n1278), .C2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1266), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1278), .A2(new_n1285), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1263), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1277), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1263), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1277), .B(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1288), .A2(new_n1293), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G390), .A2(G387), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1256), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G393), .A2(G396), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1259), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT125), .ZN(new_n1303));
  XOR2_X1   g1103(.A(new_n1300), .B(new_n1303), .Z(new_n1304));
  NAND2_X1  g1104(.A1(new_n1298), .A2(new_n1304), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1300), .B(new_n1303), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  OAI21_X1  g1107(.A(KEYINPUT63), .B1(new_n1286), .B2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1292), .A2(KEYINPUT124), .A3(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1308), .A3(new_n1297), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1305), .A2(new_n1311), .ZN(G405));
  INV_X1    g1112(.A(new_n1258), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1278), .B1(new_n1230), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT127), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT127), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1316), .B(new_n1278), .C1(new_n1230), .C2(new_n1313), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1315), .A2(new_n1291), .A3(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1314), .A2(KEYINPUT127), .A3(new_n1277), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(new_n1306), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1304), .A2(new_n1319), .A3(new_n1318), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(G402));
endmodule


