//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT76), .B(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n224), .A3(KEYINPUT79), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT2), .B1(new_n215), .B2(new_n217), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n214), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n217), .A3(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n222), .B1(new_n221), .B2(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(KEYINPUT3), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n213), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n238));
  INV_X1    g037(.A(G228gat), .ZN(new_n239));
  INV_X1    g038(.A(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT29), .B1(new_n210), .B2(new_n211), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244));
  OR2_X1    g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n244), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n225), .A2(new_n228), .B1(new_n234), .B2(new_n233), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n242), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n229), .A2(KEYINPUT81), .A3(new_n235), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT81), .B1(new_n229), .B2(new_n235), .ZN(new_n252));
  OAI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n241), .B1(new_n253), .B2(new_n238), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT84), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n256));
  AOI211_X1 g055(.A(new_n256), .B(new_n241), .C1(new_n238), .C2(new_n253), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n250), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT31), .B(G50gat), .Z(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n259), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n250), .B(new_n261), .C1(new_n255), .C2(new_n257), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n265), .A3(new_n262), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G226gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n270), .A2(new_n240), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT24), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n273), .A2(G183gat), .A3(G190gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G183gat), .B(G190gat), .ZN(new_n275));
  OAI211_X1 g074(.A(KEYINPUT25), .B(new_n274), .C1(new_n275), .C2(new_n273), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT23), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(G169gat), .B2(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT66), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G190gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n285), .B1(new_n290), .B2(KEYINPUT24), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n279), .B1(new_n277), .B2(KEYINPUT23), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n280), .A2(G169gat), .A3(G176gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n291), .A2(new_n294), .A3(new_n295), .A4(KEYINPUT25), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n283), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n292), .B2(new_n293), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n278), .A2(KEYINPUT65), .A3(new_n281), .A4(new_n279), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n291), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(G183gat), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n306), .B2(G183gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n286), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(KEYINPUT68), .A3(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n320));
  OR3_X1    g119(.A1(new_n319), .A2(new_n277), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n277), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(new_n319), .B2(new_n277), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n325), .A2(new_n284), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n298), .A2(new_n304), .B1(new_n318), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n272), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT77), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n304), .A2(new_n283), .A3(new_n296), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n318), .A2(new_n326), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(new_n271), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT77), .B(new_n272), .C1(new_n330), .C2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n328), .B(new_n212), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n327), .A2(new_n272), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n271), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n213), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n335), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT78), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n335), .A2(new_n339), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n335), .A2(new_n339), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT30), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n335), .A2(new_n339), .A3(new_n351), .A4(new_n344), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362));
  AND2_X1   g161(.A1(G113gat), .A2(G120gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(G113gat), .A2(G120gat), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n363), .A2(new_n364), .A3(KEYINPUT1), .ZN(new_n365));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT71), .B1(new_n363), .B2(new_n364), .ZN(new_n368));
  INV_X1    g167(.A(G113gat), .ZN(new_n369));
  INV_X1    g168(.A(G120gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g171(.A1(G113gat), .A2(G120gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT1), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n374), .A3(new_n375), .A4(new_n366), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n375), .A3(new_n373), .ZN(new_n377));
  INV_X1    g176(.A(G134gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G127gat), .ZN(new_n379));
  INV_X1    g178(.A(G127gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G134gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(KEYINPUT70), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n376), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n249), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n361), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n249), .B2(new_n246), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n237), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(KEYINPUT72), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT72), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n367), .A2(new_n376), .A3(new_n392), .A4(new_n383), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR4_X1   g193(.A1(new_n394), .A2(new_n251), .A3(new_n252), .A4(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n236), .A2(new_n384), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n360), .B1(new_n397), .B2(new_n386), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT5), .B1(new_n398), .B2(KEYINPUT82), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n400), .B(new_n360), .C1(new_n397), .C2(new_n386), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT83), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n249), .B(new_n384), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(new_n360), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(KEYINPUT82), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .A4(KEYINPUT5), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n396), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n251), .A2(new_n252), .ZN(new_n409));
  INV_X1    g208(.A(new_n394), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n387), .ZN(new_n412));
  OAI22_X1  g211(.A1(new_n237), .A2(new_n389), .B1(new_n386), .B2(new_n387), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n415), .A2(KEYINPUT5), .A3(new_n361), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n359), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT40), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n360), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT39), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n415), .B2(new_n361), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT39), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT4), .B1(new_n409), .B2(new_n410), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(new_n361), .C1(new_n423), .C2(new_n413), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n358), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n418), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n423), .A2(new_n413), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT39), .B(new_n419), .C1(new_n427), .C2(new_n360), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n428), .A2(KEYINPUT40), .A3(new_n358), .A4(new_n424), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n417), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n354), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n348), .A2(new_n353), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n426), .A2(new_n429), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n417), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n269), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n345), .B1(new_n340), .B2(KEYINPUT37), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n213), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n439), .A2(new_n213), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n328), .B(new_n212), .C1(new_n272), .C2(new_n327), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT87), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT37), .B(new_n441), .C1(new_n442), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n438), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT88), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n438), .A2(new_n445), .A3(new_n449), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n402), .A2(new_n407), .ZN(new_n452));
  INV_X1    g251(.A(new_n396), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n415), .A2(KEYINPUT5), .A3(new_n361), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(new_n358), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n417), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT6), .B(new_n359), .C1(new_n408), .C2(new_n416), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(new_n459), .A3(new_n349), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n341), .A2(KEYINPUT37), .A3(new_n347), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT38), .B1(new_n461), .B2(new_n437), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n451), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n436), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n466));
  NAND2_X1  g265(.A1(G227gat), .A2(G233gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT64), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n332), .A2(new_n394), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n330), .A2(new_n331), .A3(new_n391), .A4(new_n393), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT32), .ZN(new_n473));
  XOR2_X1   g272(.A(G71gat), .B(G99gat), .Z(new_n474));
  XNOR2_X1  g273(.A(G15gat), .B(G43gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n476), .B2(KEYINPUT33), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n302), .A2(new_n303), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n297), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n325), .A2(new_n284), .ZN(new_n482));
  INV_X1    g281(.A(new_n317), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n312), .B2(new_n313), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(new_n315), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n481), .A2(new_n394), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n330), .A2(new_n331), .B1(new_n391), .B2(new_n393), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n468), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n477), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n473), .A2(KEYINPUT33), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n479), .A2(new_n489), .B1(new_n491), .B2(new_n476), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n469), .A3(new_n471), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT34), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n465), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n492), .B2(KEYINPUT74), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n489), .ZN(new_n498));
  INV_X1    g297(.A(new_n490), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n476), .B1(new_n472), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n498), .A2(KEYINPUT74), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(KEYINPUT75), .B(new_n496), .C1(new_n497), .C2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT73), .B1(new_n488), .B2(new_n477), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n472), .A2(new_n466), .A3(new_n478), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n500), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n505), .A2(new_n494), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n492), .A2(new_n495), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n465), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT74), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n492), .A2(KEYINPUT74), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(new_n494), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT75), .B1(new_n513), .B2(new_n496), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n458), .A2(new_n459), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n354), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n509), .A2(new_n515), .B1(new_n517), .B2(new_n269), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n432), .B1(new_n458), .B2(new_n459), .ZN(new_n519));
  INV_X1    g318(.A(new_n268), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n265), .B1(new_n260), .B2(new_n262), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n492), .A2(new_n495), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n519), .A2(new_n522), .A3(new_n513), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n494), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n523), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n269), .A2(KEYINPUT35), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n519), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n464), .A2(new_n518), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT14), .ZN(new_n532));
  OR2_X1    g331(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(KEYINPUT91), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  OR2_X1    g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G43gat), .A2(G50gat), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G29gat), .ZN(new_n539));
  INV_X1    g338(.A(G36gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT90), .B(G50gat), .Z(new_n543));
  OAI211_X1 g342(.A(new_n535), .B(new_n537), .C1(new_n543), .C2(G43gat), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n533), .A2(new_n534), .A3(new_n542), .A4(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n538), .B1(new_n532), .B2(new_n541), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT17), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT16), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(G1gat), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(G1gat), .B2(new_n549), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G8gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n548), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n547), .A2(new_n553), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT18), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n547), .B(new_n553), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n556), .B(KEYINPUT13), .Z(new_n562));
  AOI22_X1  g361(.A1(new_n558), .A2(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G169gat), .B(G197gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT12), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n560), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n560), .B2(new_n563), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT94), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT96), .B(G92gat), .Z(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT8), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT95), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(KEYINPUT95), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT98), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n590), .A2(new_n597), .A3(new_n592), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(new_n594), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT99), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n603), .A3(new_n591), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n548), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(KEYINPUT100), .A3(new_n548), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT101), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n605), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n614), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(new_n610), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n580), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n612), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n613), .A3(new_n615), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n579), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G57gat), .B(G64gat), .Z(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(KEYINPUT92), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(KEYINPUT9), .B2(new_n624), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(G231gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n380), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n553), .B1(KEYINPUT21), .B2(new_n630), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT93), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G155gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n636), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n630), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n605), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n596), .B2(new_n598), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n601), .A2(KEYINPUT102), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n601), .A2(KEYINPUT102), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n645), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n647), .A2(KEYINPUT10), .A3(new_n602), .A4(new_n604), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n645), .A2(new_n650), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n655), .A2(new_n658), .A3(new_n662), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR4_X1   g465(.A1(new_n530), .A2(new_n573), .A3(new_n643), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n516), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g469(.A(KEYINPUT16), .B(G8gat), .Z(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(new_n432), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n667), .ZN(new_n673));
  OAI21_X1  g472(.A(G8gat), .B1(new_n673), .B2(new_n354), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n672), .ZN(new_n675));
  MUX2_X1   g474(.A(new_n672), .B(new_n675), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g475(.A(new_n527), .ZN(new_n677));
  AOI21_X1  g476(.A(G15gat), .B1(new_n667), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n502), .A2(new_n508), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n514), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n667), .A2(G15gat), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n679), .A2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n269), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT43), .B(G22gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  OAI22_X1  g485(.A1(new_n680), .A2(new_n514), .B1(new_n519), .B2(new_n522), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n687), .B1(new_n463), .B2(new_n436), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n524), .A2(KEYINPUT35), .B1(new_n528), .B2(new_n519), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT104), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n464), .A2(new_n518), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n525), .A2(new_n529), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n623), .A2(KEYINPUT44), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n690), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n530), .B2(new_n623), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n666), .A2(new_n642), .ZN(new_n699));
  INV_X1    g498(.A(new_n573), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n698), .A2(KEYINPUT105), .A3(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n516), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n530), .A2(new_n623), .A3(new_n701), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(new_n539), .A3(new_n668), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1328gat));
  OAI21_X1  g511(.A(G36gat), .B1(new_n707), .B2(new_n354), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n709), .A2(new_n540), .A3(new_n432), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(G1329gat));
  AOI21_X1  g515(.A(KEYINPUT105), .B1(new_n698), .B2(new_n702), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n704), .B(new_n701), .C1(new_n696), .C2(new_n697), .ZN(new_n718));
  INV_X1    g517(.A(new_n681), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT107), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n681), .A3(new_n706), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(G43gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n709), .A2(new_n721), .A3(new_n677), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G43gat), .B1(new_n703), .B2(new_n719), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(new_n543), .B1(new_n703), .B2(new_n522), .ZN(new_n733));
  INV_X1    g532(.A(new_n623), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n522), .A2(new_n543), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n699), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n530), .A2(new_n573), .A3(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n705), .A2(new_n269), .A3(new_n706), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(new_n741), .B2(new_n543), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n690), .A2(new_n694), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n664), .A2(new_n665), .ZN(new_n745));
  NOR4_X1   g544(.A1(new_n744), .A2(new_n700), .A3(new_n643), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n668), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  INV_X1    g547(.A(new_n746), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n432), .B(KEYINPUT108), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n749), .A2(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n750), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT49), .B(G64gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n746), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT109), .Z(G1333gat));
  OAI21_X1  g555(.A(G71gat), .B1(new_n749), .B2(new_n719), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n527), .A2(G71gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n749), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n269), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT111), .B(G78gat), .Z(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n642), .A2(new_n700), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n698), .A2(new_n666), .A3(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(new_n668), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n734), .B(new_n765), .C1(new_n688), .C2(new_n689), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n666), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n668), .A2(new_n582), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n767), .A2(new_n582), .B1(new_n772), .B2(new_n773), .ZN(G1336gat));
  AOI21_X1  g573(.A(new_n581), .B1(new_n766), .B2(new_n432), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n750), .A2(G92gat), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n775), .A2(KEYINPUT112), .B1(new_n772), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n775), .A2(KEYINPUT112), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT52), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n766), .A2(new_n752), .ZN(new_n781));
  OAI221_X1 g580(.A(new_n780), .B1(new_n772), .B2(new_n776), .C1(new_n781), .C2(new_n581), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1337gat));
  AND2_X1   g582(.A1(new_n766), .A2(new_n681), .ZN(new_n784));
  INV_X1    g583(.A(G99gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n677), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n784), .A2(new_n785), .B1(new_n772), .B2(new_n786), .ZN(G1338gat));
  AND2_X1   g586(.A1(new_n766), .A2(new_n269), .ZN(new_n788));
  INV_X1    g587(.A(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n269), .A2(new_n789), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n788), .A2(new_n789), .B1(new_n772), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g591(.A(new_n642), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n651), .A2(new_n657), .A3(new_n652), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n657), .B1(new_n651), .B2(new_n652), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n653), .A2(new_n797), .A3(new_n654), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n663), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n794), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n651), .A2(new_n657), .A3(new_n652), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n655), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n662), .B1(new_n796), .B2(new_n797), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n801), .A2(new_n700), .A3(new_n665), .A4(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n561), .A2(new_n562), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n568), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT114), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(KEYINPUT114), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n570), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n664), .B2(new_n665), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n734), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n805), .A2(new_n665), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT55), .B1(new_n803), .B2(new_n804), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n816), .A2(new_n623), .A3(new_n817), .A4(new_n812), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n793), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n623), .A2(new_n642), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n573), .A4(new_n745), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n745), .A2(new_n623), .A3(new_n573), .A4(new_n642), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n516), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n522), .A2(new_n513), .A3(new_n523), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n750), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n700), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n269), .B(new_n527), .C1(new_n819), .C2(new_n825), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n668), .A3(new_n750), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT115), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n573), .A2(new_n369), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n831), .B1(new_n835), .B2(new_n836), .ZN(G1340gat));
  AOI21_X1  g636(.A(G120gat), .B1(new_n830), .B2(new_n666), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n745), .A2(new_n370), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n835), .B2(new_n839), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n834), .B2(new_n793), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n830), .A2(new_n380), .A3(new_n642), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NAND4_X1  g642(.A1(new_n829), .A2(new_n378), .A3(new_n354), .A4(new_n734), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n834), .B2(new_n623), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  NAND2_X1  g646(.A1(new_n819), .A2(new_n825), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n269), .ZN(new_n849));
  XNOR2_X1  g648(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n853), .A3(new_n269), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n752), .A2(new_n681), .A3(new_n516), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(new_n700), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT58), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n681), .A2(new_n522), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n826), .A2(new_n858), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(KEYINPUT118), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n752), .A2(G141gat), .A3(new_n573), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g663(.A1(KEYINPUT119), .A2(new_n860), .A3(new_n863), .A4(new_n861), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n857), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n859), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n856), .A2(G141gat), .B1(new_n867), .B2(new_n863), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n869), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n866), .B1(new_n872), .B2(new_n873), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n860), .A2(new_n861), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n752), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n216), .A3(new_n666), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n745), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(KEYINPUT59), .A3(new_n216), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT59), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n522), .B(new_n850), .C1(new_n819), .C2(new_n825), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n848), .A2(new_n269), .A3(new_n851), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT121), .ZN(new_n886));
  INV_X1    g685(.A(new_n823), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n805), .A2(new_n665), .ZN(new_n888));
  INV_X1    g687(.A(new_n812), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n888), .A2(new_n734), .A3(new_n889), .A4(new_n801), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n803), .A2(new_n804), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n573), .B1(new_n891), .B2(new_n794), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n813), .B1(new_n888), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(new_n734), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n887), .B1(new_n894), .B2(new_n793), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n853), .B1(new_n895), .B2(new_n522), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n884), .A2(new_n886), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n666), .B1(new_n855), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n898), .B2(new_n855), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n881), .B1(new_n901), .B2(G148gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n877), .B1(new_n880), .B2(new_n902), .ZN(G1345gat));
  INV_X1    g702(.A(G155gat), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n876), .A2(new_n904), .A3(new_n642), .ZN(new_n905));
  OAI21_X1  g704(.A(G155gat), .B1(new_n878), .B2(new_n793), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1346gat));
  OAI21_X1  g706(.A(G162gat), .B1(new_n878), .B2(new_n623), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n623), .A2(G162gat), .A3(new_n432), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n875), .B2(new_n909), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n668), .A2(new_n354), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n832), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(G169gat), .A3(new_n700), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n668), .B(new_n750), .C1(new_n819), .C2(new_n825), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n914), .A2(new_n828), .ZN(new_n915));
  AOI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n700), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(new_n916), .ZN(G1348gat));
  INV_X1    g716(.A(G176gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n918), .A3(new_n666), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n832), .A2(new_n911), .ZN(new_n920));
  OAI21_X1  g719(.A(G176gat), .B1(new_n920), .B2(new_n745), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1349gat));
  NAND2_X1  g721(.A1(new_n306), .A2(G183gat), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n915), .A2(new_n316), .A3(new_n923), .A4(new_n642), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n920), .B2(new_n793), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(G183gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n920), .A2(new_n925), .A3(new_n793), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n920), .B2(new_n623), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n288), .A3(new_n734), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n914), .A2(new_n858), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(KEYINPUT123), .B(G197gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n700), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n719), .A2(new_n911), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n819), .A2(new_n823), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT57), .B1(new_n940), .B2(new_n269), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n941), .B1(KEYINPUT121), .B2(new_n885), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n939), .B1(new_n942), .B2(new_n884), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(KEYINPUT124), .A3(new_n700), .ZN(new_n944));
  INV_X1    g743(.A(new_n937), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(KEYINPUT124), .B1(new_n943), .B2(new_n700), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n938), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n943), .A2(new_n666), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n914), .A2(new_n951), .A3(new_n666), .A4(new_n858), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n954), .A3(KEYINPUT125), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT125), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n951), .B1(new_n943), .B2(new_n666), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n953), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n955), .A2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n936), .A2(new_n204), .A3(new_n642), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n642), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  INV_X1    g763(.A(G218gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n965), .B1(new_n935), .B2(new_n623), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  INV_X1    g766(.A(new_n939), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n896), .B1(new_n882), .B2(new_n883), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n885), .A2(KEYINPUT121), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n967), .B(new_n968), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n623), .A2(new_n203), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n967), .B1(new_n897), .B2(new_n968), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n966), .C1(new_n973), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1355gat));
endmodule


