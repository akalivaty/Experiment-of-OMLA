

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  NAND2_X1 U323 ( .A1(n525), .A2(n489), .ZN(n450) );
  NAND2_X1 U324 ( .A1(n541), .A2(n543), .ZN(n374) );
  NAND2_X1 U325 ( .A1(n538), .A2(n520), .ZN(n524) );
  INV_X1 U326 ( .A(n578), .ZN(n444) );
  INV_X1 U327 ( .A(n516), .ZN(n525) );
  NOR2_X1 U328 ( .A1(n455), .A2(n510), .ZN(n538) );
  XOR2_X2 U329 ( .A(n441), .B(n440), .Z(n516) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n426) );
  XOR2_X1 U331 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n319) );
  XNOR2_X1 U332 ( .A(n307), .B(n306), .ZN(n308) );
  INV_X1 U333 ( .A(n353), .ZN(n306) );
  NOR2_X1 U334 ( .A1(n585), .A2(n462), .ZN(n463) );
  XNOR2_X1 U335 ( .A(n402), .B(n401), .ZN(n537) );
  XNOR2_X1 U336 ( .A(n314), .B(n313), .ZN(n315) );
  INV_X1 U337 ( .A(KEYINPUT87), .ZN(n313) );
  XNOR2_X1 U338 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U339 ( .A(n425), .B(KEYINPUT55), .ZN(n442) );
  XNOR2_X1 U340 ( .A(n574), .B(n373), .ZN(n543) );
  XOR2_X1 U341 ( .A(KEYINPUT94), .B(n466), .Z(n493) );
  XOR2_X1 U342 ( .A(G64GAT), .B(G92GAT), .Z(n291) );
  XOR2_X1 U343 ( .A(KEYINPUT89), .B(n449), .Z(n292) );
  XNOR2_X1 U344 ( .A(G29GAT), .B(G134GAT), .ZN(n301) );
  NOR2_X1 U345 ( .A1(n549), .A2(n394), .ZN(n395) );
  INV_X1 U346 ( .A(KEYINPUT115), .ZN(n404) );
  XNOR2_X1 U347 ( .A(n404), .B(KEYINPUT54), .ZN(n405) );
  XNOR2_X1 U348 ( .A(n376), .B(n315), .ZN(n317) );
  XNOR2_X1 U349 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U350 ( .A(KEYINPUT41), .ZN(n373) );
  NOR2_X1 U351 ( .A1(n292), .A2(n460), .ZN(n474) );
  INV_X1 U352 ( .A(n543), .ZN(n555) );
  XOR2_X1 U353 ( .A(KEYINPUT86), .B(n458), .Z(n510) );
  INV_X1 U354 ( .A(G183GAT), .ZN(n445) );
  XNOR2_X1 U355 ( .A(n443), .B(KEYINPUT116), .ZN(n559) );
  INV_X1 U356 ( .A(G43GAT), .ZN(n467) );
  XOR2_X1 U357 ( .A(n408), .B(n323), .Z(n513) );
  XNOR2_X1 U358 ( .A(n445), .B(KEYINPUT118), .ZN(n446) );
  XNOR2_X1 U359 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U360 ( .A(n447), .B(n446), .ZN(G1350GAT) );
  XNOR2_X1 U361 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U362 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n294) );
  XNOR2_X1 U363 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n293) );
  XNOR2_X1 U364 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U365 ( .A(n295), .B(G155GAT), .Z(n297) );
  XNOR2_X1 U366 ( .A(G141GAT), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U367 ( .A(n297), .B(n296), .ZN(n414) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(KEYINPUT85), .Z(n299) );
  XNOR2_X1 U369 ( .A(KEYINPUT6), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U370 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U371 ( .A(n414), .B(n300), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n301), .B(G85GAT), .ZN(n339) );
  XOR2_X1 U373 ( .A(n339), .B(KEYINPUT84), .Z(n303) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U375 ( .A(n303), .B(n302), .ZN(n309) );
  XOR2_X1 U376 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n305) );
  XOR2_X1 U377 ( .A(KEYINPUT0), .B(G127GAT), .Z(n427) );
  XOR2_X1 U378 ( .A(G120GAT), .B(G57GAT), .Z(n370) );
  XNOR2_X1 U379 ( .A(n427), .B(n370), .ZN(n304) );
  XNOR2_X1 U380 ( .A(n305), .B(n304), .ZN(n307) );
  XOR2_X1 U381 ( .A(G113GAT), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U382 ( .A(n311), .B(n310), .ZN(n458) );
  INV_X1 U383 ( .A(n510), .ZN(n485) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n312) );
  XNOR2_X1 U385 ( .A(n312), .B(G211GAT), .ZN(n408) );
  XOR2_X1 U386 ( .A(G8GAT), .B(G183GAT), .Z(n376) );
  NAND2_X1 U387 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U389 ( .A(n316), .B(G218GAT), .ZN(n336) );
  XOR2_X1 U390 ( .A(n317), .B(n336), .Z(n322) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n318) );
  XNOR2_X1 U392 ( .A(G176GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U393 ( .A(n291), .B(n320), .ZN(n362) );
  XNOR2_X1 U394 ( .A(n426), .B(n362), .ZN(n321) );
  XNOR2_X1 U395 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U396 ( .A(n513), .B(KEYINPUT114), .Z(n403) );
  XNOR2_X1 U397 ( .A(KEYINPUT108), .B(KEYINPUT48), .ZN(n402) );
  XOR2_X1 U398 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n325) );
  XNOR2_X1 U399 ( .A(G162GAT), .B(G92GAT), .ZN(n324) );
  XNOR2_X1 U400 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U401 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n327) );
  XNOR2_X1 U402 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n326) );
  XNOR2_X1 U403 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U404 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n331) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U407 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U408 ( .A(KEYINPUT10), .B(n332), .ZN(n333) );
  XNOR2_X1 U409 ( .A(n334), .B(n333), .ZN(n343) );
  XNOR2_X1 U410 ( .A(G99GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U411 ( .A(n335), .B(KEYINPUT69), .ZN(n363) );
  XOR2_X1 U412 ( .A(n336), .B(n363), .Z(n341) );
  XOR2_X1 U413 ( .A(G43GAT), .B(G50GAT), .Z(n338) );
  XNOR2_X1 U414 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U415 ( .A(n338), .B(n337), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n350), .B(n339), .ZN(n340) );
  XNOR2_X1 U417 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U418 ( .A(n343), .B(n342), .Z(n560) );
  INV_X1 U419 ( .A(n560), .ZN(n549) );
  XOR2_X1 U420 ( .A(G22GAT), .B(G141GAT), .Z(n345) );
  XNOR2_X1 U421 ( .A(G169GAT), .B(G15GAT), .ZN(n344) );
  XNOR2_X1 U422 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U423 ( .A(G8GAT), .B(KEYINPUT30), .Z(n347) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(KEYINPUT67), .ZN(n346) );
  XNOR2_X1 U425 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U426 ( .A(n349), .B(n348), .ZN(n358) );
  XOR2_X1 U427 ( .A(n350), .B(KEYINPUT29), .Z(n352) );
  NAND2_X1 U428 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U429 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U430 ( .A(n354), .B(n353), .Z(n356) );
  XNOR2_X1 U431 ( .A(G36GAT), .B(G29GAT), .ZN(n355) );
  XNOR2_X1 U432 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U433 ( .A(n358), .B(n357), .ZN(n541) );
  XOR2_X1 U434 ( .A(KEYINPUT32), .B(KEYINPUT68), .Z(n360) );
  NAND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U436 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U437 ( .A(n361), .B(KEYINPUT31), .Z(n365) );
  XNOR2_X1 U438 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U439 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(G85GAT), .Z(n367) );
  XNOR2_X1 U441 ( .A(G148GAT), .B(G78GAT), .ZN(n366) );
  XNOR2_X1 U442 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U443 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U444 ( .A(G71GAT), .B(KEYINPUT13), .Z(n375) );
  XNOR2_X1 U445 ( .A(n370), .B(n375), .ZN(n371) );
  XNOR2_X1 U446 ( .A(n372), .B(n371), .ZN(n574) );
  XNOR2_X1 U447 ( .A(n374), .B(KEYINPUT46), .ZN(n393) );
  XOR2_X1 U448 ( .A(n376), .B(n375), .Z(n378) );
  XNOR2_X1 U449 ( .A(G15GAT), .B(G127GAT), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U451 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n380) );
  NAND2_X1 U452 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U453 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U454 ( .A(n382), .B(n381), .Z(n384) );
  XOR2_X1 U455 ( .A(G22GAT), .B(G78GAT), .Z(n418) );
  XNOR2_X1 U456 ( .A(n418), .B(KEYINPUT75), .ZN(n383) );
  XNOR2_X1 U457 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U458 ( .A(G57GAT), .B(G211GAT), .Z(n386) );
  XNOR2_X1 U459 ( .A(G1GAT), .B(G155GAT), .ZN(n385) );
  XNOR2_X1 U460 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U461 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n388) );
  XNOR2_X1 U462 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n387) );
  XNOR2_X1 U463 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U464 ( .A(n390), .B(n389), .Z(n391) );
  XOR2_X1 U465 ( .A(n392), .B(n391), .Z(n578) );
  NAND2_X1 U466 ( .A1(n393), .A2(n444), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n395), .B(KEYINPUT47), .ZN(n400) );
  XOR2_X1 U468 ( .A(KEYINPUT36), .B(n549), .Z(n585) );
  NOR2_X1 U469 ( .A1(n585), .A2(n444), .ZN(n396) );
  XOR2_X1 U470 ( .A(KEYINPUT45), .B(n396), .Z(n397) );
  NOR2_X1 U471 ( .A1(n574), .A2(n397), .ZN(n398) );
  INV_X1 U472 ( .A(n541), .ZN(n569) );
  NAND2_X1 U473 ( .A1(n398), .A2(n569), .ZN(n399) );
  NAND2_X1 U474 ( .A1(n400), .A2(n399), .ZN(n401) );
  NAND2_X1 U475 ( .A1(n403), .A2(n537), .ZN(n406) );
  NOR2_X1 U476 ( .A1(n485), .A2(n407), .ZN(n568) );
  XOR2_X1 U477 ( .A(KEYINPUT81), .B(n408), .Z(n410) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n424) );
  XOR2_X1 U480 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n412) );
  XNOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U483 ( .A(n414), .B(n413), .ZN(n422) );
  XOR2_X1 U484 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n416) );
  XNOR2_X1 U485 ( .A(G218GAT), .B(G106GAT), .ZN(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U487 ( .A(n417), .B(G204GAT), .Z(n420) );
  XNOR2_X1 U488 ( .A(G50GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U489 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U490 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U491 ( .A(n424), .B(n423), .ZN(n453) );
  NAND2_X1 U492 ( .A1(n568), .A2(n453), .ZN(n425) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U495 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U496 ( .A(KEYINPUT64), .B(G71GAT), .Z(n431) );
  XNOR2_X1 U497 ( .A(G113GAT), .B(G15GAT), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n441) );
  XOR2_X1 U500 ( .A(G134GAT), .B(G190GAT), .Z(n435) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U503 ( .A(G120GAT), .B(G176GAT), .Z(n437) );
  XNOR2_X1 U504 ( .A(KEYINPUT20), .B(G183GAT), .ZN(n436) );
  XNOR2_X1 U505 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U506 ( .A(n439), .B(n438), .Z(n440) );
  NAND2_X1 U507 ( .A1(n442), .A2(n525), .ZN(n443) );
  NOR2_X1 U508 ( .A1(n559), .A2(n444), .ZN(n447) );
  XOR2_X1 U509 ( .A(KEYINPUT95), .B(KEYINPUT38), .Z(n465) );
  NOR2_X1 U510 ( .A1(n574), .A2(n569), .ZN(n475) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(KEYINPUT88), .Z(n448) );
  XOR2_X1 U512 ( .A(n513), .B(n448), .Z(n455) );
  XOR2_X1 U513 ( .A(KEYINPUT28), .B(n453), .Z(n492) );
  INV_X1 U514 ( .A(n492), .ZN(n520) );
  NOR2_X1 U515 ( .A1(n525), .A2(n524), .ZN(n449) );
  INV_X1 U516 ( .A(n513), .ZN(n489) );
  XNOR2_X1 U517 ( .A(n450), .B(KEYINPUT90), .ZN(n451) );
  NAND2_X1 U518 ( .A1(n451), .A2(n453), .ZN(n452) );
  XNOR2_X1 U519 ( .A(n452), .B(KEYINPUT25), .ZN(n457) );
  NOR2_X1 U520 ( .A1(n525), .A2(n453), .ZN(n454) );
  XOR2_X1 U521 ( .A(KEYINPUT26), .B(n454), .Z(n566) );
  NOR2_X1 U522 ( .A1(n566), .A2(n455), .ZN(n456) );
  NOR2_X1 U523 ( .A1(n457), .A2(n456), .ZN(n459) );
  NOR2_X1 U524 ( .A1(n459), .A2(n458), .ZN(n460) );
  NOR2_X1 U525 ( .A1(n578), .A2(n474), .ZN(n461) );
  XNOR2_X1 U526 ( .A(n461), .B(KEYINPUT93), .ZN(n462) );
  XOR2_X1 U527 ( .A(KEYINPUT37), .B(n463), .Z(n509) );
  NAND2_X1 U528 ( .A1(n475), .A2(n509), .ZN(n464) );
  XNOR2_X1 U529 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n493), .A2(n525), .ZN(n470) );
  XOR2_X1 U531 ( .A(KEYINPUT98), .B(KEYINPUT40), .Z(n468) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(KEYINPUT77), .Z(n472) );
  NAND2_X1 U533 ( .A1(n578), .A2(n560), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n497) );
  NAND2_X1 U536 ( .A1(n475), .A2(n497), .ZN(n482) );
  NOR2_X1 U537 ( .A1(n510), .A2(n482), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT34), .B(n476), .Z(n477) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n513), .A2(n482), .ZN(n479) );
  XNOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT91), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(G1325GAT) );
  NOR2_X1 U543 ( .A1(n516), .A2(n482), .ZN(n481) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U546 ( .A1(n520), .A2(n482), .ZN(n483) );
  XOR2_X1 U547 ( .A(KEYINPUT92), .B(n483), .Z(n484) );
  XNOR2_X1 U548 ( .A(G22GAT), .B(n484), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n485), .A2(n493), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n486) );
  XNOR2_X1 U551 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n488), .B(G29GAT), .ZN(G1328GAT) );
  XOR2_X1 U553 ( .A(G36GAT), .B(KEYINPUT97), .Z(n491) );
  NAND2_X1 U554 ( .A1(n493), .A2(n489), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT99), .Z(n495) );
  NAND2_X1 U557 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(G1331GAT) );
  NOR2_X1 U559 ( .A1(n555), .A2(n541), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT100), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n497), .A2(n508), .ZN(n504) );
  NOR2_X1 U562 ( .A1(n510), .A2(n504), .ZN(n499) );
  XNOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT101), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n513), .A2(n504), .ZN(n501) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(n501), .Z(n502) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n502), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n516), .A2(n504), .ZN(n503) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n503), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n520), .A2(n504), .ZN(n506) );
  XNOR2_X1 U572 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n505) );
  XNOR2_X1 U573 ( .A(n506), .B(n505), .ZN(n507) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n507), .Z(G1335GAT) );
  NAND2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n510), .A2(n519), .ZN(n511) );
  XOR2_X1 U577 ( .A(n511), .B(KEYINPUT104), .Z(n512) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n512), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n519), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(n517), .Z(n518) );
  XNOR2_X1 U584 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XOR2_X1 U589 ( .A(G113GAT), .B(KEYINPUT109), .Z(n528) );
  NAND2_X1 U590 ( .A1(n525), .A2(n537), .ZN(n526) );
  NOR2_X1 U591 ( .A1(n524), .A2(n526), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n534), .A2(n541), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT49), .B(KEYINPUT110), .Z(n530) );
  NAND2_X1 U595 ( .A1(n534), .A2(n543), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n578), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n532), .B(KEYINPUT50), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n549), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U605 ( .A1(n566), .A2(n539), .ZN(n540) );
  XOR2_X1 U606 ( .A(KEYINPUT111), .B(n540), .Z(n550) );
  NAND2_X1 U607 ( .A1(n550), .A2(n541), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U610 ( .A1(n550), .A2(n543), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n578), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT112), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n548), .ZN(G1346GAT) );
  XOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT113), .Z(n552) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1347GAT) );
  NOR2_X1 U619 ( .A1(n559), .A2(n569), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(KEYINPUT117), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  NOR2_X1 U622 ( .A1(n559), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(n558), .ZN(G1349GAT) );
  XNOR2_X1 U626 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n573) );
  INV_X1 U633 ( .A(n566), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n569), .A2(n584), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n576) );
  INV_X1 U640 ( .A(n584), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT124), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n583) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

