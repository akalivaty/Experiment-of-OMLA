

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XOR2_X1 U323 ( .A(n364), .B(n363), .Z(n527) );
  XOR2_X1 U324 ( .A(n442), .B(n356), .Z(n291) );
  INV_X1 U325 ( .A(KEYINPUT101), .ZN(n382) );
  XNOR2_X1 U326 ( .A(n382), .B(KEYINPUT25), .ZN(n383) );
  XNOR2_X1 U327 ( .A(n384), .B(n383), .ZN(n388) );
  XNOR2_X1 U328 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n474) );
  INV_X1 U329 ( .A(n448), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U332 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n414) );
  XNOR2_X1 U333 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U334 ( .A(n415), .B(n414), .ZN(n498) );
  INV_X1 U335 ( .A(G190GAT), .ZN(n480) );
  INV_X1 U336 ( .A(G106GAT), .ZN(n457) );
  XNOR2_X1 U337 ( .A(n379), .B(n378), .ZN(n534) );
  XNOR2_X1 U338 ( .A(n480), .B(KEYINPUT58), .ZN(n481) );
  XNOR2_X1 U339 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U340 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(G15GAT), .B(G1GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n292), .B(KEYINPUT71), .ZN(n422) );
  XNOR2_X1 U343 ( .A(G8GAT), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n293), .B(KEYINPUT78), .ZN(n356) );
  XNOR2_X1 U345 ( .A(n422), .B(n356), .ZN(n312) );
  XOR2_X1 U346 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n295) );
  XNOR2_X1 U347 ( .A(G22GAT), .B(G211GAT), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U349 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n297) );
  XNOR2_X1 U350 ( .A(KEYINPUT80), .B(KEYINPUT82), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U352 ( .A(n299), .B(n298), .Z(n310) );
  XOR2_X1 U353 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n301) );
  XNOR2_X1 U354 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n308) );
  XOR2_X1 U356 ( .A(KEYINPUT13), .B(G57GAT), .Z(n443) );
  XOR2_X1 U357 ( .A(G78GAT), .B(G155GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(G127GAT), .B(G71GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U360 ( .A(n443), .B(n304), .Z(n306) );
  NAND2_X1 U361 ( .A1(G231GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U363 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n578) );
  INV_X1 U366 ( .A(n578), .ZN(n566) );
  XOR2_X1 U367 ( .A(KEYINPUT92), .B(KEYINPUT95), .Z(n314) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n314), .B(n313), .ZN(n323) );
  XOR2_X1 U370 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n321) );
  XOR2_X1 U371 ( .A(KEYINPUT0), .B(G134GAT), .Z(n316) );
  XNOR2_X1 U372 ( .A(KEYINPUT85), .B(G127GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U374 ( .A(G113GAT), .B(n317), .Z(n365) );
  XOR2_X1 U375 ( .A(G155GAT), .B(KEYINPUT2), .Z(n319) );
  XNOR2_X1 U376 ( .A(KEYINPUT3), .B(KEYINPUT91), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n338) );
  XNOR2_X1 U378 ( .A(n365), .B(n338), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n335) );
  NAND2_X1 U381 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XOR2_X1 U382 ( .A(G148GAT), .B(G162GAT), .Z(n325) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(G120GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U385 ( .A(G29GAT), .B(G85GAT), .Z(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U387 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U388 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n331) );
  XNOR2_X1 U389 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n525) );
  XOR2_X1 U393 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n337) );
  XNOR2_X1 U394 ( .A(G218GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n346) );
  XOR2_X1 U396 ( .A(G148GAT), .B(G78GAT), .Z(n446) );
  XOR2_X1 U397 ( .A(n446), .B(n338), .Z(n344) );
  XOR2_X1 U398 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n339), .B(G162GAT), .ZN(n400) );
  XOR2_X1 U401 ( .A(n400), .B(KEYINPUT23), .Z(n341) );
  NAND2_X1 U402 ( .A1(G228GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U403 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n419), .B(n342), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n351) );
  XNOR2_X1 U407 ( .A(G211GAT), .B(KEYINPUT90), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n347), .B(KEYINPUT89), .ZN(n348) );
  XOR2_X1 U409 ( .A(n348), .B(KEYINPUT21), .Z(n350) );
  XNOR2_X1 U410 ( .A(G197GAT), .B(G204GAT), .ZN(n349) );
  XOR2_X1 U411 ( .A(n350), .B(n349), .Z(n355) );
  XNOR2_X1 U412 ( .A(n351), .B(n355), .ZN(n477) );
  XOR2_X1 U413 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n353) );
  XNOR2_X1 U414 ( .A(KEYINPUT18), .B(KEYINPUT86), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U416 ( .A(G169GAT), .B(n354), .Z(n366) );
  XOR2_X1 U417 ( .A(n366), .B(n355), .Z(n364) );
  XOR2_X1 U418 ( .A(G176GAT), .B(G64GAT), .Z(n442) );
  NAND2_X1 U419 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n291), .B(n357), .ZN(n358) );
  XOR2_X1 U421 ( .A(n358), .B(KEYINPUT97), .Z(n362) );
  XOR2_X1 U422 ( .A(G92GAT), .B(G218GAT), .Z(n360) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(G190GAT), .ZN(n359) );
  XNOR2_X1 U424 ( .A(n360), .B(n359), .ZN(n397) );
  XNOR2_X1 U425 ( .A(n397), .B(KEYINPUT96), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n379) );
  XOR2_X1 U428 ( .A(KEYINPUT87), .B(G99GAT), .Z(n368) );
  XNOR2_X1 U429 ( .A(G43GAT), .B(G190GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U431 ( .A(KEYINPUT20), .B(KEYINPUT64), .Z(n370) );
  XNOR2_X1 U432 ( .A(G15GAT), .B(KEYINPUT88), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U434 ( .A(n372), .B(n371), .Z(n377) );
  XOR2_X1 U435 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XOR2_X1 U436 ( .A(G183GAT), .B(G176GAT), .Z(n374) );
  NAND2_X1 U437 ( .A1(G227GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n447), .B(n375), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n378) );
  AND2_X1 U441 ( .A1(n527), .A2(n534), .ZN(n380) );
  XOR2_X1 U442 ( .A(KEYINPUT100), .B(n380), .Z(n381) );
  NAND2_X1 U443 ( .A1(n477), .A2(n381), .ZN(n384) );
  XNOR2_X1 U444 ( .A(n527), .B(KEYINPUT27), .ZN(n390) );
  NOR2_X1 U445 ( .A1(n477), .A2(n534), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U447 ( .A1(n390), .A2(n568), .ZN(n386) );
  XNOR2_X1 U448 ( .A(KEYINPUT99), .B(n386), .ZN(n387) );
  NOR2_X1 U449 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U450 ( .A1(n525), .A2(n389), .ZN(n394) );
  XNOR2_X1 U451 ( .A(KEYINPUT28), .B(n477), .ZN(n537) );
  NAND2_X1 U452 ( .A1(n525), .A2(n390), .ZN(n531) );
  NOR2_X1 U453 ( .A1(n534), .A2(n531), .ZN(n391) );
  NAND2_X1 U454 ( .A1(n537), .A2(n391), .ZN(n392) );
  XOR2_X1 U455 ( .A(KEYINPUT98), .B(n392), .Z(n393) );
  NOR2_X1 U456 ( .A1(n394), .A2(n393), .ZN(n486) );
  XOR2_X1 U457 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n396) );
  XNOR2_X1 U458 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n398) );
  XOR2_X1 U460 ( .A(n398), .B(n397), .Z(n402) );
  XNOR2_X1 U461 ( .A(G99GAT), .B(G106GAT), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n399), .B(G85GAT), .ZN(n448) );
  XNOR2_X1 U463 ( .A(n400), .B(n448), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U465 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n404) );
  NAND2_X1 U466 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U468 ( .A(n406), .B(n405), .Z(n412) );
  XNOR2_X1 U469 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n407), .B(G29GAT), .ZN(n408) );
  XOR2_X1 U471 ( .A(n408), .B(KEYINPUT70), .Z(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n430) );
  XNOR2_X1 U474 ( .A(n430), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n557) );
  XOR2_X1 U476 ( .A(KEYINPUT77), .B(n557), .Z(n544) );
  XNOR2_X1 U477 ( .A(KEYINPUT36), .B(n544), .ZN(n583) );
  NOR2_X1 U478 ( .A1(n486), .A2(n583), .ZN(n413) );
  NAND2_X1 U479 ( .A1(n566), .A2(n413), .ZN(n415) );
  XOR2_X1 U480 ( .A(G8GAT), .B(G197GAT), .Z(n417) );
  XNOR2_X1 U481 ( .A(G36GAT), .B(G50GAT), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U483 ( .A(n418), .B(G113GAT), .Z(n421) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n426) );
  XOR2_X1 U486 ( .A(n422), .B(KEYINPUT30), .Z(n424) );
  NAND2_X1 U487 ( .A1(G229GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U489 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U490 ( .A(KEYINPUT68), .B(KEYINPUT72), .Z(n428) );
  XNOR2_X1 U491 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n570) );
  INV_X1 U495 ( .A(n570), .ZN(n455) );
  XOR2_X1 U496 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n434) );
  XNOR2_X1 U497 ( .A(G204GAT), .B(G92GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n454) );
  XNOR2_X1 U499 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n436) );
  AND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  NAND2_X1 U502 ( .A1(n437), .A2(KEYINPUT74), .ZN(n441) );
  INV_X1 U503 ( .A(n437), .ZN(n439) );
  INV_X1 U504 ( .A(KEYINPUT74), .ZN(n438) );
  NAND2_X1 U505 ( .A1(n439), .A2(n438), .ZN(n440) );
  NAND2_X1 U506 ( .A1(n441), .A2(n440), .ZN(n445) );
  XOR2_X1 U507 ( .A(n443), .B(n442), .Z(n444) );
  XNOR2_X1 U508 ( .A(n445), .B(n444), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n450) );
  XOR2_X1 U510 ( .A(n454), .B(n453), .Z(n574) );
  XNOR2_X1 U511 ( .A(n574), .B(KEYINPUT41), .ZN(n562) );
  NOR2_X1 U512 ( .A1(n455), .A2(n562), .ZN(n509) );
  NAND2_X1 U513 ( .A1(n498), .A2(n509), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT113), .ZN(n529) );
  INV_X1 U515 ( .A(n537), .ZN(n521) );
  NAND2_X1 U516 ( .A1(n529), .A2(n521), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT114), .B(KEYINPUT44), .Z(n458) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(G1339GAT) );
  XOR2_X1 U519 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n462) );
  NOR2_X1 U520 ( .A1(n570), .A2(n562), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n463), .A2(n578), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT116), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n465), .A2(n557), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT47), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n583), .A2(n566), .ZN(n467) );
  XNOR2_X1 U527 ( .A(KEYINPUT45), .B(n467), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n468), .A2(n570), .ZN(n469) );
  NOR2_X1 U529 ( .A1(n469), .A2(n574), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT48), .ZN(n532) );
  XOR2_X1 U532 ( .A(n527), .B(KEYINPUT122), .Z(n473) );
  NOR2_X1 U533 ( .A1(n532), .A2(n473), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n525), .A2(n476), .ZN(n569) );
  NAND2_X1 U535 ( .A1(n569), .A2(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT55), .B(n478), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n479), .A2(n534), .ZN(n565) );
  NOR2_X1 U538 ( .A1(n544), .A2(n565), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT103), .ZN(n490) );
  NAND2_X1 U541 ( .A1(n544), .A2(n578), .ZN(n484) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n484), .ZN(n485) );
  NOR2_X1 U543 ( .A1(n486), .A2(n485), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT102), .B(n487), .Z(n511) );
  NOR2_X1 U545 ( .A1(n570), .A2(n574), .ZN(n497) );
  INV_X1 U546 ( .A(n497), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n511), .A2(n488), .ZN(n495) );
  NAND2_X1 U548 ( .A1(n495), .A2(n525), .ZN(n489) );
  XOR2_X1 U549 ( .A(n490), .B(n489), .Z(G1324GAT) );
  NAND2_X1 U550 ( .A1(n527), .A2(n495), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n492), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n494) );
  NAND2_X1 U554 ( .A1(n495), .A2(n534), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n521), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n499) );
  XOR2_X1 U559 ( .A(KEYINPUT38), .B(n499), .Z(n507) );
  NAND2_X1 U560 ( .A1(n507), .A2(n525), .ZN(n502) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT107), .Z(n504) );
  NAND2_X1 U565 ( .A1(n507), .A2(n527), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n534), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U570 ( .A1(n521), .A2(n507), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  INV_X1 U572 ( .A(n509), .ZN(n510) );
  NOR2_X1 U573 ( .A1(n511), .A2(n510), .ZN(n522) );
  NAND2_X1 U574 ( .A1(n522), .A2(n525), .ZN(n514) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(KEYINPUT108), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n527), .A2(n522), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U580 ( .A(G71GAT), .B(KEYINPUT109), .Z(n517) );
  NAND2_X1 U581 ( .A1(n522), .A2(n534), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT110), .B(n520), .Z(n524) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n529), .A2(n525), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n527), .A2(n529), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n529), .A2(n534), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U596 ( .A(n533), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U597 ( .A1(n534), .A2(n548), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(n535), .Z(n536) );
  NAND2_X1 U599 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n570), .A2(n543), .ZN(n538) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  NOR2_X1 U602 ( .A1(n562), .A2(n543), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n566), .A2(n543), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n541), .Z(n542) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U609 ( .A(KEYINPUT119), .B(KEYINPUT51), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n568), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n570), .A2(n556), .ZN(n549) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n562), .A2(n556), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n566), .A2(n556), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NOR2_X1 U625 ( .A1(n570), .A2(n565), .ZN(n559) );
  XOR2_X1 U626 ( .A(G169GAT), .B(n559), .Z(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n561) );
  XNOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n562), .A2(n565), .ZN(n563) );
  XOR2_X1 U631 ( .A(n564), .B(n563), .Z(G1349GAT) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(G183GAT), .B(n567), .Z(G1350GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n582) );
  NOR2_X1 U635 ( .A1(n570), .A2(n582), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U640 ( .A(n582), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n579), .A2(n574), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

