//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(KEYINPUT81), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G113gat), .B2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT72), .B(G120gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n209), .B(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G113gat), .A2(G120gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n207), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G127gat), .ZN(new_n219));
  INV_X1    g018(.A(G127gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G134gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n217), .A2(KEYINPUT71), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT71), .B1(new_n217), .B2(new_n222), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n213), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G155gat), .ZN(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G141gat), .B(G148gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g031(.A(G155gat), .B(G162gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT79), .ZN(new_n234));
  INV_X1    g033(.A(G141gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(new_n235), .A3(G148gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(G148gat), .ZN(new_n237));
  INV_X1    g036(.A(G148gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G141gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n233), .B(new_n236), .C1(new_n240), .C2(new_n234), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(KEYINPUT80), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT80), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G162gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n246), .B2(G155gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n232), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n250));
  INV_X1    g049(.A(new_n216), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n208), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n252), .B2(new_n210), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n217), .A2(KEYINPUT71), .A3(new_n222), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT80), .B(G162gat), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT2), .B1(new_n256), .B2(new_n228), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n231), .A2(KEYINPUT79), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n236), .A2(new_n227), .A3(new_n229), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(new_n260), .A3(new_n213), .A4(new_n232), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n249), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n206), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI211_X1 g064(.A(KEYINPUT81), .B(new_n263), .C1(new_n249), .C2(new_n261), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n260), .A2(new_n269), .A3(new_n232), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n225), .A3(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n225), .A2(new_n248), .A3(KEYINPUT4), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n211), .A2(new_n212), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n222), .A2(new_n208), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n253), .A2(new_n254), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n233), .B1(new_n242), .B2(new_n240), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT79), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n236), .A2(new_n227), .A3(new_n229), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n280), .B2(new_n257), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n273), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n271), .B(new_n263), .C1(new_n272), .C2(new_n282), .ZN(new_n283));
  XOR2_X1   g082(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT83), .B1(new_n267), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n248), .A2(KEYINPUT3), .B1(new_n255), .B2(new_n213), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n264), .B1(new_n288), .B2(new_n270), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n261), .A2(KEYINPUT4), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n276), .A2(new_n281), .A3(new_n273), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n284), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT83), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n293), .B(new_n294), .C1(new_n265), .C2(new_n266), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n295), .ZN(new_n296));
  MUX2_X1   g095(.A(new_n292), .B(new_n290), .S(KEYINPUT84), .Z(new_n297));
  AND2_X1   g096(.A1(new_n289), .A2(new_n284), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n205), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT89), .B1(new_n300), .B2(KEYINPUT6), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n287), .A2(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT6), .ZN(new_n304));
  NOR4_X1   g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n205), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G176gat), .ZN(new_n310));
  INV_X1    g109(.A(G169gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT65), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT65), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G169gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT23), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(KEYINPUT64), .ZN(new_n326));
  INV_X1    g125(.A(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n325), .A2(new_n326), .A3(new_n329), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n320), .A3(KEYINPUT66), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n323), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(new_n330), .B2(KEYINPUT67), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(KEYINPUT67), .B2(new_n330), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n327), .A3(new_n328), .ZN(new_n344));
  OAI21_X1  g143(.A(KEYINPUT68), .B1(G183gat), .B2(G190gat), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n344), .A2(new_n324), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n340), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n328), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n351), .B(KEYINPUT28), .Z(new_n352));
  INV_X1    g151(.A(KEYINPUT26), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n316), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n319), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n355), .A2(KEYINPUT70), .B1(new_n353), .B2(new_n338), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(KEYINPUT70), .B2(new_n355), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(new_n357), .A3(new_n330), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n307), .B(new_n308), .C1(new_n359), .C2(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT69), .B1(new_n337), .B2(new_n348), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n362), .B(new_n347), .C1(new_n335), .C2(new_n336), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n308), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT29), .B1(new_n349), .B2(new_n358), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT76), .B1(new_n367), .B2(new_n365), .ZN(new_n368));
  XNOR2_X1  g167(.A(G197gat), .B(G204gat), .ZN(new_n369));
  INV_X1    g168(.A(G211gat), .ZN(new_n370));
  INV_X1    g169(.A(G218gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(KEYINPUT22), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G211gat), .B(G218gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n366), .A3(new_n368), .A4(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n365), .A2(KEYINPUT29), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n364), .A2(new_n378), .B1(new_n359), .B2(new_n365), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n375), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT37), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(G8gat), .B(G36gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT77), .ZN(new_n386));
  XOR2_X1   g185(.A(G64gat), .B(G92gat), .Z(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n381), .B2(KEYINPUT37), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT38), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n382), .A2(new_n383), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT38), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n383), .B1(new_n379), .B2(new_n376), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n360), .A2(new_n368), .A3(new_n366), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n393), .B1(new_n376), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n391), .A2(new_n392), .A3(new_n388), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n388), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n267), .A2(new_n286), .A3(KEYINPUT83), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n262), .A2(new_n264), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n262), .A2(new_n206), .A3(new_n264), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n294), .B1(new_n402), .B2(new_n293), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n299), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n205), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT6), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n302), .A2(new_n205), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n397), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n306), .A2(new_n390), .A3(new_n396), .A4(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n269), .B1(new_n375), .B2(KEYINPUT29), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n248), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT29), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n270), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n375), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n270), .A2(KEYINPUT85), .A3(new_n412), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT85), .B1(new_n270), .B2(new_n412), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n419), .A2(new_n376), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n411), .A2(G228gat), .A3(G233gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(KEYINPUT86), .B(G22gat), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OR2_X1    g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n427), .A3(new_n425), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n423), .B2(new_n425), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G78gat), .B(G106gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT31), .B(G50gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n423), .A2(G22gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n381), .B2(new_n388), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n440), .B(new_n443), .C1(new_n381), .C2(new_n388), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n381), .A2(new_n388), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n282), .A2(KEYINPUT84), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n271), .B(new_n447), .C1(new_n292), .C2(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n264), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(KEYINPUT39), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(new_n405), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT39), .B1(new_n262), .B2(new_n264), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT88), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n452), .A2(KEYINPUT88), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n449), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n451), .A2(KEYINPUT40), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT40), .B1(new_n451), .B2(new_n455), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(new_n300), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n446), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n409), .A2(new_n439), .A3(new_n459), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n406), .A2(new_n407), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n300), .A2(KEYINPUT6), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n439), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT36), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n276), .B(new_n358), .C1(new_n361), .C2(new_n363), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n315), .A2(new_n320), .A3(KEYINPUT66), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT66), .B1(new_n315), .B2(new_n320), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT25), .B1(new_n476), .B2(new_n333), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n362), .B1(new_n477), .B2(new_n347), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n337), .A2(KEYINPUT69), .A3(new_n348), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n276), .A4(new_n358), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n364), .A2(new_n225), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n487));
  XNOR2_X1  g286(.A(G15gat), .B(G43gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G99gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n491), .B2(KEYINPUT33), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n470), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n492), .ZN(new_n494));
  AOI211_X1 g293(.A(KEYINPUT74), .B(new_n494), .C1(new_n483), .C2(new_n485), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n483), .A2(new_n485), .B1(new_n487), .B2(KEYINPUT33), .ZN(new_n496));
  OAI22_X1  g295(.A1(new_n493), .A2(new_n495), .B1(new_n496), .B2(new_n490), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n473), .A2(new_n481), .A3(new_n484), .A4(new_n482), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  OAI221_X1 g301(.A(new_n500), .B1(new_n496), .B2(new_n490), .C1(new_n493), .C2(new_n495), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n469), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT75), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT75), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n506), .A3(new_n501), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n504), .B1(new_n508), .B2(new_n469), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n502), .A2(new_n503), .A3(new_n439), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT35), .B1(new_n465), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n463), .A2(new_n303), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n300), .A2(KEYINPUT89), .A3(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n462), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT35), .B1(new_n435), .B2(new_n438), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n461), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n468), .A2(new_n509), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT13), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT16), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n524), .B(KEYINPUT91), .C1(G1gat), .C2(new_n521), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n521), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n527), .A3(G8gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT92), .B(G8gat), .Z(new_n529));
  OAI211_X1 g328(.A(new_n524), .B(new_n529), .C1(G1gat), .C2(new_n521), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G43gat), .B(G50gat), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n534));
  INV_X1    g333(.A(G29gat), .ZN(new_n535));
  INV_X1    g334(.A(G36gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT14), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G29gat), .B2(G36gat), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(KEYINPUT15), .ZN(new_n541));
  NAND2_X1  g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT90), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n534), .A2(new_n540), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n539), .A3(new_n542), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT15), .A3(new_n533), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n520), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(KEYINPUT17), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n545), .A2(new_n554), .A3(new_n547), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n531), .A2(KEYINPUT93), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT93), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n558), .A3(new_n530), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(new_n519), .A3(new_n551), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n552), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g362(.A1(new_n528), .A2(new_n558), .A3(new_n530), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n558), .B1(new_n528), .B2(new_n530), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n566), .A2(new_n556), .B1(new_n550), .B2(new_n531), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT18), .A4(new_n519), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n560), .A2(KEYINPUT18), .A3(new_n519), .A4(new_n551), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT94), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G197gat), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT11), .B(G169gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT12), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n569), .A3(new_n571), .A4(new_n577), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n518), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  OAI21_X1  g386(.A(G92gat), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n589), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n588), .A2(new_n590), .B1(new_n586), .B2(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT8), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT98), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n594), .B2(new_n593), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(G99gat), .A2(G106gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(new_n593), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT99), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n601), .A3(new_n593), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n591), .A2(new_n596), .B1(new_n600), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n585), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n603), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n591), .A2(new_n596), .A3(new_n600), .A4(new_n602), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(KEYINPUT100), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n548), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n584), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n604), .A2(new_n605), .A3(new_n585), .ZN(new_n614));
  AOI21_X1  g413(.A(KEYINPUT100), .B1(new_n607), .B2(new_n608), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n550), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(KEYINPUT102), .A3(new_n611), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  INV_X1    g418(.A(new_n555), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n554), .B1(new_n545), .B2(new_n547), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n609), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n556), .A2(KEYINPUT101), .A3(new_n609), .A4(new_n606), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G190gat), .B(G218gat), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n618), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n618), .B2(new_n626), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT97), .ZN(new_n633));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n618), .A2(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n627), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n618), .A2(new_n626), .A3(new_n628), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n635), .B(new_n631), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G57gat), .B(G64gat), .Z(new_n643));
  INV_X1    g442(.A(KEYINPUT9), .ZN(new_n644));
  INV_X1    g443(.A(G71gat), .ZN(new_n645));
  INV_X1    g444(.A(G78gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(G71gat), .B(G78gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n643), .A2(new_n649), .A3(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT96), .B(KEYINPUT19), .Z(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  OAI21_X1  g456(.A(new_n532), .B1(new_n654), .B2(new_n653), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G127gat), .B(G155gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT20), .ZN(new_n661));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT95), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n661), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n659), .B(new_n666), .ZN(new_n667));
  OR3_X1    g466(.A1(new_n642), .A2(KEYINPUT104), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT104), .B1(new_n642), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(G230gat), .ZN(new_n671));
  INV_X1    g470(.A(G233gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n653), .B1(new_n604), .B2(new_n605), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n607), .A2(new_n652), .A3(new_n651), .A4(new_n608), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT10), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n651), .A2(KEYINPUT10), .A3(new_n652), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n606), .B2(new_n609), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n674), .B1(new_n677), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n675), .A2(new_n676), .A3(new_n673), .ZN(new_n682));
  XNOR2_X1  g481(.A(G120gat), .B(G148gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT105), .ZN(new_n684));
  XNOR2_X1  g483(.A(G176gat), .B(G204gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n681), .B2(new_n682), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n583), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n464), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n522), .ZN(G1324gat));
  OAI21_X1  g493(.A(G8gat), .B1(new_n692), .B2(new_n461), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n696));
  INV_X1    g495(.A(new_n692), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT16), .B(G8gat), .Z(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n446), .A3(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n699), .A2(KEYINPUT106), .A3(new_n696), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT106), .B1(new_n699), .B2(new_n696), .ZN(new_n701));
  OAI221_X1 g500(.A(new_n695), .B1(new_n696), .B2(new_n699), .C1(new_n700), .C2(new_n701), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n692), .B2(new_n509), .ZN(new_n703));
  INV_X1    g502(.A(G15gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n508), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n692), .B2(new_n705), .ZN(G1326gat));
  OR3_X1    g505(.A1(new_n692), .A2(KEYINPUT107), .A3(new_n439), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n692), .B2(new_n439), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT43), .B(G22gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  INV_X1    g511(.A(new_n642), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n518), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n460), .A2(new_n467), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT36), .B1(new_n505), .B2(new_n507), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n504), .A3(new_n716), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n517), .A2(new_n511), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n642), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n667), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n582), .A2(new_n721), .A3(new_n690), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n464), .ZN(new_n724));
  INV_X1    g523(.A(new_n464), .ZN(new_n725));
  INV_X1    g524(.A(new_n690), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n642), .A2(new_n726), .A3(new_n667), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT108), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n583), .A2(new_n535), .A3(new_n725), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT109), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n724), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1328gat));
  OAI21_X1  g534(.A(G36gat), .B1(new_n723), .B2(new_n461), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n737));
  AOI211_X1 g536(.A(G36gat), .B(new_n461), .C1(new_n737), .C2(KEYINPUT46), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n583), .A2(new_n728), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n737), .A2(KEYINPUT46), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(G43gat), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n583), .A2(new_n743), .A3(new_n508), .A4(new_n728), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT111), .ZN(new_n745));
  INV_X1    g544(.A(new_n509), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n714), .A2(new_n719), .A3(new_n746), .A4(new_n722), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1330gat));
  NAND2_X1  g550(.A1(new_n466), .A2(G50gat), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n583), .A2(new_n466), .A3(new_n728), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n723), .A2(new_n752), .B1(G50gat), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g554(.A1(new_n518), .A2(new_n581), .A3(new_n670), .A4(new_n726), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n725), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G57gat), .ZN(G1332gat));
  INV_X1    g557(.A(KEYINPUT49), .ZN(new_n759));
  INV_X1    g558(.A(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n446), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT112), .Z(new_n762));
  NAND2_X1  g561(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n760), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n763), .B(new_n764), .ZN(G1333gat));
  NAND3_X1  g564(.A1(new_n756), .A2(new_n645), .A3(new_n508), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n756), .A2(new_n746), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n645), .ZN(new_n768));
  XOR2_X1   g567(.A(new_n768), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n466), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n721), .A2(new_n581), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n726), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n720), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775), .B2(new_n464), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n773), .B1(KEYINPUT113), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n642), .B(new_n778), .C1(new_n717), .C2(new_n718), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n777), .A2(KEYINPUT113), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n517), .A2(new_n511), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n746), .B2(new_n715), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(new_n642), .A3(new_n778), .A4(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n725), .A2(new_n587), .A3(new_n690), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n776), .B1(new_n787), .B2(new_n788), .ZN(G1336gat));
  NOR3_X1   g588(.A1(new_n461), .A2(G92gat), .A3(new_n726), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n781), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n714), .A2(new_n719), .A3(new_n446), .A4(new_n774), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(new_n794), .B2(G92gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n781), .A2(KEYINPUT114), .A3(new_n785), .A4(new_n790), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT115), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n794), .A2(G92gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n775), .A2(new_n509), .ZN(new_n806));
  XOR2_X1   g605(.A(KEYINPUT116), .B(G99gat), .Z(new_n807));
  NAND3_X1  g606(.A1(new_n508), .A2(new_n690), .A3(new_n807), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n806), .A2(new_n807), .B1(new_n787), .B2(new_n808), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n720), .A2(new_n466), .A3(new_n774), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n439), .A2(G106gat), .A3(new_n726), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n811), .B(new_n812), .C1(new_n787), .C2(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n813), .B(KEYINPUT117), .Z(new_n815));
  AOI22_X1  g614(.A1(new_n810), .A2(G106gat), .B1(new_n786), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n812), .ZN(G1339gat));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n567), .A2(new_n519), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n549), .A2(new_n551), .A3(new_n520), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n576), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n580), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n642), .A2(new_n822), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n677), .A2(new_n679), .A3(new_n674), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(KEYINPUT54), .A3(new_n680), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n826), .B(new_n674), .C1(new_n677), .C2(new_n679), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n827), .A2(new_n828), .A3(new_n686), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n827), .B2(new_n686), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n687), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT55), .B(new_n825), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n818), .B1(new_n823), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n580), .A2(new_n821), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n641), .B2(new_n636), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n838), .A2(KEYINPUT119), .A3(new_n834), .A4(new_n833), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n581), .A2(new_n833), .A3(new_n834), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n690), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n642), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n667), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n668), .A2(new_n582), .A3(new_n669), .A4(new_n726), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(new_n439), .A3(new_n508), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n464), .A2(new_n446), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n212), .A3(new_n582), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n846), .A2(new_n725), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n446), .A3(new_n510), .ZN(new_n852));
  AOI21_X1  g651(.A(G113gat), .B1(new_n852), .B2(new_n581), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n850), .A2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n849), .B2(new_n726), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n211), .A3(new_n690), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n849), .B2(new_n667), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n852), .A2(new_n220), .A3(new_n721), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n218), .A3(new_n642), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  OAI21_X1  g661(.A(G134gat), .B1(new_n849), .B2(new_n713), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  AND2_X1   g664(.A1(new_n509), .A2(new_n848), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n846), .B2(new_n466), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n868), .B(new_n439), .C1(new_n844), .C2(new_n845), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n870), .B2(new_n582), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n509), .A2(new_n466), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n851), .A2(new_n873), .A3(KEYINPUT121), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n851), .B2(new_n873), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n461), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n582), .A2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n871), .B(new_n872), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n851), .A2(new_n873), .A3(new_n446), .A4(new_n878), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n870), .A2(KEYINPUT120), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n882), .B(new_n866), .C1(new_n867), .C2(new_n869), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(new_n581), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n884), .B2(G141gat), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n879), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g687(.A(KEYINPUT122), .B(new_n879), .C1(new_n885), .C2(new_n872), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(new_n876), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n238), .A3(new_n690), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n823), .A2(new_n835), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT123), .B1(new_n843), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n667), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n843), .A2(new_n894), .A3(KEYINPUT123), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n845), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n466), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n899), .A2(new_n869), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n690), .A3(new_n866), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(G148gat), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n893), .B1(new_n902), .B2(KEYINPUT59), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT124), .B(new_n904), .C1(new_n901), .C2(G148gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n881), .A2(new_n883), .ZN(new_n907));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n238), .C1(new_n907), .C2(new_n690), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n892), .B1(new_n906), .B2(new_n908), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n891), .A2(new_n228), .A3(new_n721), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n907), .A2(new_n721), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n228), .ZN(G1346gat));
  AOI21_X1  g711(.A(new_n246), .B1(new_n891), .B2(new_n642), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n713), .A2(new_n256), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n907), .B2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n725), .A2(new_n461), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n847), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n582), .ZN(new_n918));
  INV_X1    g717(.A(new_n510), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n846), .A2(new_n919), .A3(new_n916), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n581), .A2(new_n312), .A3(new_n314), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1348gat));
  OAI21_X1  g721(.A(G176gat), .B1(new_n917), .B2(new_n726), .ZN(new_n923));
  INV_X1    g722(.A(new_n920), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n318), .A3(new_n690), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n917), .B2(new_n667), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n721), .A2(new_n350), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n924), .A2(KEYINPUT125), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT125), .B1(new_n924), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n917), .B2(new_n713), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n924), .A2(new_n328), .A3(new_n642), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT126), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n934), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G1351gat));
  AND2_X1   g738(.A1(new_n509), .A2(new_n916), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(new_n466), .A3(new_n846), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n581), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n900), .A2(new_n940), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n581), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n943), .B2(new_n690), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n941), .A2(new_n946), .A3(new_n690), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n947), .A2(new_n949), .ZN(G1353gat));
  NAND3_X1  g749(.A1(new_n941), .A2(new_n370), .A3(new_n721), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n721), .B(new_n940), .C1(new_n899), .C2(new_n869), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT127), .Z(G1354gat));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n371), .A3(new_n642), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n943), .A2(new_n642), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n371), .ZN(G1355gat));
endmodule


