

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X2 U322 ( .A(KEYINPUT41), .B(n571), .ZN(n494) );
  XNOR2_X1 U323 ( .A(n374), .B(n290), .ZN(n375) );
  XNOR2_X1 U324 ( .A(KEYINPUT38), .B(n439), .ZN(n490) );
  XNOR2_X1 U325 ( .A(n360), .B(n359), .ZN(n513) );
  AND2_X1 U326 ( .A1(G231GAT), .A2(G233GAT), .ZN(n290) );
  AND2_X1 U327 ( .A1(n578), .A2(n575), .ZN(n450) );
  XOR2_X1 U328 ( .A(G176GAT), .B(G64GAT), .Z(n433) );
  INV_X1 U329 ( .A(KEYINPUT89), .ZN(n352) );
  XNOR2_X1 U330 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U331 ( .A(n458), .B(KEYINPUT48), .ZN(n459) );
  XNOR2_X1 U332 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U333 ( .A(n460), .B(n459), .ZN(n538) );
  XNOR2_X1 U334 ( .A(n355), .B(n354), .ZN(n358) );
  XNOR2_X1 U335 ( .A(n387), .B(n386), .ZN(n575) );
  INV_X1 U336 ( .A(G29GAT), .ZN(n440) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n469) );
  XNOR2_X1 U338 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U339 ( .A(n470), .B(n469), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n443), .B(n442), .ZN(G1328GAT) );
  XOR2_X1 U341 ( .A(G57GAT), .B(G148GAT), .Z(n292) );
  XNOR2_X1 U342 ( .A(G1GAT), .B(G155GAT), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U344 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n294) );
  XNOR2_X1 U345 ( .A(KEYINPUT84), .B(KEYINPUT6), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(n296), .B(n295), .Z(n301) );
  XOR2_X1 U348 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n298) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(KEYINPUT5), .B(n299), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U353 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n303) );
  XNOR2_X1 U354 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n320) );
  XOR2_X1 U356 ( .A(G85GAT), .B(n320), .Z(n305) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U359 ( .A(n307), .B(n306), .Z(n313) );
  XNOR2_X1 U360 ( .A(G127GAT), .B(KEYINPUT77), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n308), .B(KEYINPUT0), .ZN(n309) );
  XOR2_X1 U362 ( .A(n309), .B(KEYINPUT76), .Z(n311) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n343) );
  XNOR2_X1 U365 ( .A(n343), .B(G120GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n563) );
  XOR2_X1 U367 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n408) );
  INV_X1 U368 ( .A(n563), .ZN(n497) );
  XOR2_X1 U369 ( .A(G162GAT), .B(KEYINPUT71), .Z(n315) );
  XNOR2_X1 U370 ( .A(G50GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n400) );
  XOR2_X1 U372 ( .A(G211GAT), .B(KEYINPUT82), .Z(n317) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n317), .B(n316), .ZN(n356) );
  XNOR2_X1 U375 ( .A(n400), .B(n356), .ZN(n329) );
  XOR2_X1 U376 ( .A(G78GAT), .B(G148GAT), .Z(n319) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n430) );
  XNOR2_X1 U379 ( .A(n320), .B(n430), .ZN(n327) );
  XOR2_X1 U380 ( .A(G22GAT), .B(G155GAT), .Z(n374) );
  XOR2_X1 U381 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n322) );
  XNOR2_X1 U382 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U384 ( .A(n374), .B(n323), .Z(n325) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U388 ( .A(n329), .B(n328), .ZN(n462) );
  XOR2_X1 U389 ( .A(G120GAT), .B(G71GAT), .Z(n425) );
  XOR2_X1 U390 ( .A(G176GAT), .B(G99GAT), .Z(n331) );
  XNOR2_X1 U391 ( .A(G43GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U393 ( .A(n425), .B(n332), .Z(n334) );
  NAND2_X1 U394 ( .A1(G227GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U396 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n336) );
  XNOR2_X1 U397 ( .A(G15GAT), .B(KEYINPUT78), .ZN(n335) );
  XNOR2_X1 U398 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U399 ( .A(n338), .B(n337), .Z(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n339) );
  XNOR2_X1 U401 ( .A(n339), .B(KEYINPUT17), .ZN(n340) );
  XOR2_X1 U402 ( .A(n340), .B(KEYINPUT79), .Z(n342) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U404 ( .A(n342), .B(n341), .ZN(n360) );
  XNOR2_X1 U405 ( .A(n343), .B(n360), .ZN(n344) );
  XNOR2_X1 U406 ( .A(n345), .B(n344), .ZN(n525) );
  INV_X1 U407 ( .A(n525), .ZN(n516) );
  XOR2_X1 U408 ( .A(KEYINPUT87), .B(KEYINPUT90), .Z(n347) );
  XNOR2_X1 U409 ( .A(G8GAT), .B(G204GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U411 ( .A(n433), .B(G92GAT), .Z(n349) );
  XOR2_X1 U412 ( .A(G36GAT), .B(G190GAT), .Z(n389) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(n389), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U415 ( .A(n351), .B(n350), .Z(n355) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n356), .B(KEYINPUT88), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  NOR2_X1 U419 ( .A1(n516), .A2(n513), .ZN(n361) );
  NOR2_X1 U420 ( .A1(n462), .A2(n361), .ZN(n362) );
  XOR2_X1 U421 ( .A(KEYINPUT25), .B(n362), .Z(n366) );
  XNOR2_X1 U422 ( .A(KEYINPUT27), .B(n513), .ZN(n368) );
  XOR2_X1 U423 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n364) );
  NAND2_X1 U424 ( .A1(n462), .A2(n516), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n566) );
  NOR2_X1 U426 ( .A1(n368), .A2(n566), .ZN(n365) );
  NOR2_X1 U427 ( .A1(n366), .A2(n365), .ZN(n367) );
  NOR2_X1 U428 ( .A1(n497), .A2(n367), .ZN(n372) );
  NOR2_X1 U429 ( .A1(n563), .A2(n368), .ZN(n369) );
  XOR2_X1 U430 ( .A(KEYINPUT91), .B(n369), .Z(n540) );
  XOR2_X1 U431 ( .A(n462), .B(KEYINPUT28), .Z(n519) );
  NAND2_X1 U432 ( .A1(n540), .A2(n519), .ZN(n523) );
  NOR2_X1 U433 ( .A1(n525), .A2(n523), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n370), .B(KEYINPUT92), .ZN(n371) );
  NOR2_X1 U435 ( .A1(n372), .A2(n371), .ZN(n474) );
  XOR2_X1 U436 ( .A(G15GAT), .B(G1GAT), .Z(n373) );
  XNOR2_X1 U437 ( .A(n373), .B(G8GAT), .ZN(n409) );
  INV_X1 U438 ( .A(n409), .ZN(n376) );
  XOR2_X1 U439 ( .A(G57GAT), .B(KEYINPUT13), .Z(n424) );
  XOR2_X1 U440 ( .A(n377), .B(n424), .Z(n379) );
  XNOR2_X1 U441 ( .A(G127GAT), .B(G183GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U443 ( .A(G64GAT), .B(G78GAT), .Z(n381) );
  XNOR2_X1 U444 ( .A(G71GAT), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U446 ( .A(KEYINPUT15), .B(KEYINPUT74), .Z(n383) );
  XNOR2_X1 U447 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U449 ( .A(n385), .B(n384), .Z(n386) );
  NOR2_X1 U450 ( .A1(n474), .A2(n575), .ZN(n406) );
  XNOR2_X1 U451 ( .A(KEYINPUT36), .B(KEYINPUT96), .ZN(n405) );
  XNOR2_X1 U452 ( .A(G99GAT), .B(G85GAT), .ZN(n388) );
  XNOR2_X1 U453 ( .A(n388), .B(G92GAT), .ZN(n429) );
  XOR2_X1 U454 ( .A(n429), .B(n389), .Z(n391) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n391), .B(n390), .ZN(n404) );
  XOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n393) );
  XNOR2_X1 U458 ( .A(KEYINPUT9), .B(KEYINPUT73), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U460 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n395) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(G106GAT), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(n397), .B(n396), .Z(n402) );
  XOR2_X1 U464 ( .A(G29GAT), .B(G43GAT), .Z(n399) );
  XNOR2_X1 U465 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n410), .B(n400), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U469 ( .A(n404), .B(n403), .Z(n553) );
  INV_X1 U470 ( .A(n553), .ZN(n468) );
  XNOR2_X1 U471 ( .A(n405), .B(n468), .ZN(n578) );
  NAND2_X1 U472 ( .A1(n406), .A2(n578), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n511) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n423) );
  XOR2_X1 U475 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n412) );
  NAND2_X1 U476 ( .A1(G229GAT), .A2(G233GAT), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U478 ( .A(n413), .B(KEYINPUT67), .Z(n421) );
  XOR2_X1 U479 ( .A(G113GAT), .B(G50GAT), .Z(n415) );
  XNOR2_X1 U480 ( .A(G169GAT), .B(G36GAT), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U482 ( .A(KEYINPUT68), .B(G141GAT), .Z(n417) );
  XNOR2_X1 U483 ( .A(G22GAT), .B(G197GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n567) );
  INV_X1 U488 ( .A(n567), .ZN(n541) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n438) );
  XOR2_X1 U490 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n427) );
  NAND2_X1 U491 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n428), .B(KEYINPUT33), .Z(n432) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U496 ( .A(n434), .B(n433), .Z(n436) );
  XNOR2_X1 U497 ( .A(KEYINPUT70), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U499 ( .A(n438), .B(n437), .ZN(n571) );
  NOR2_X1 U500 ( .A1(n541), .A2(n571), .ZN(n475) );
  NAND2_X1 U501 ( .A1(n511), .A2(n475), .ZN(n439) );
  NOR2_X1 U502 ( .A1(n563), .A2(n490), .ZN(n443) );
  XNOR2_X1 U503 ( .A(KEYINPUT95), .B(KEYINPUT39), .ZN(n441) );
  INV_X1 U504 ( .A(KEYINPUT122), .ZN(n467) );
  XOR2_X1 U505 ( .A(KEYINPUT47), .B(KEYINPUT109), .Z(n448) );
  NOR2_X1 U506 ( .A1(n541), .A2(n494), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n444), .B(KEYINPUT46), .ZN(n445) );
  NOR2_X1 U508 ( .A1(n575), .A2(n445), .ZN(n446) );
  NAND2_X1 U509 ( .A1(n446), .A2(n553), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n449) );
  XNOR2_X1 U512 ( .A(KEYINPUT66), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U514 ( .A1(n452), .A2(n571), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT111), .ZN(n454) );
  NOR2_X1 U516 ( .A1(n454), .A2(n567), .ZN(n455) );
  XNOR2_X1 U517 ( .A(n455), .B(KEYINPUT112), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n457), .A2(n456), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n458) );
  NOR2_X1 U520 ( .A1(n538), .A2(n513), .ZN(n461) );
  XNOR2_X1 U521 ( .A(KEYINPUT54), .B(n461), .ZN(n564) );
  NOR2_X1 U522 ( .A1(n462), .A2(n497), .ZN(n463) );
  AND2_X1 U523 ( .A1(n564), .A2(n463), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT55), .B(n464), .Z(n465) );
  NAND2_X1 U525 ( .A1(n465), .A2(n525), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n561) );
  NAND2_X1 U527 ( .A1(n561), .A2(n468), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(KEYINPUT75), .Z(n472) );
  NAND2_X1 U529 ( .A1(n553), .A2(n575), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n495) );
  NAND2_X1 U532 ( .A1(n475), .A2(n495), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n563), .A2(n481), .ZN(n476) );
  XOR2_X1 U534 ( .A(G1GAT), .B(n476), .Z(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U536 ( .A1(n513), .A2(n481), .ZN(n478) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n478), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n516), .A2(n481), .ZN(n480) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n519), .A2(n481), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT94), .B(n482), .Z(n483) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  NOR2_X1 U544 ( .A1(n490), .A2(n513), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G36GAT), .B(n486), .ZN(G1329GAT) );
  NOR2_X1 U548 ( .A1(n490), .A2(n516), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U551 ( .A(G43GAT), .B(n489), .Z(G1330GAT) );
  XNOR2_X1 U552 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n492) );
  NOR2_X1 U553 ( .A1(n519), .A2(n490), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n493), .ZN(G1331GAT) );
  NOR2_X1 U556 ( .A1(n567), .A2(n494), .ZN(n510) );
  NAND2_X1 U557 ( .A1(n495), .A2(n510), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(KEYINPUT103), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n497), .A2(n506), .ZN(n501) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n499) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1332GAT) );
  INV_X1 U564 ( .A(n513), .ZN(n502) );
  NAND2_X1 U565 ( .A1(n502), .A2(n506), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n503), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n506), .A2(n525), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n508) );
  INV_X1 U570 ( .A(n519), .ZN(n505) );
  NAND2_X1 U571 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U575 ( .A1(n563), .A2(n518), .ZN(n512) );
  XOR2_X1 U576 ( .A(G85GAT), .B(n512), .Z(G1336GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n518), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1337GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n518), .ZN(n517) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U583 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n522), .Z(G1339GAT) );
  NOR2_X1 U586 ( .A1(n538), .A2(n523), .ZN(n524) );
  NAND2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n534) );
  NOR2_X1 U588 ( .A1(n541), .A2(n534), .ZN(n526) );
  XOR2_X1 U589 ( .A(G113GAT), .B(n526), .Z(G1340GAT) );
  NOR2_X1 U590 ( .A1(n534), .A2(n494), .ZN(n530) );
  XOR2_X1 U591 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n528) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  INV_X1 U595 ( .A(n575), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n549), .A2(n534), .ZN(n532) );
  XNOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n533), .Z(G1342GAT) );
  NOR2_X1 U600 ( .A1(n553), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U603 ( .A(G134GAT), .B(n537), .Z(G1343GAT) );
  NOR2_X1 U604 ( .A1(n538), .A2(n566), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n540), .A2(n539), .ZN(n552) );
  NOR2_X1 U606 ( .A1(n541), .A2(n552), .ZN(n542) );
  XOR2_X1 U607 ( .A(KEYINPUT118), .B(n542), .Z(n543) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U609 ( .A1(n494), .A2(n552), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n545) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT119), .B(n546), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n552), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U620 ( .A1(n561), .A2(n567), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 U622 ( .A(n494), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n556), .A2(n561), .ZN(n558) );
  XOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT123), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n575), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n579) );
  NAND2_X1 U633 ( .A1(n579), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n579), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .Z(n577) );
  NAND2_X1 U641 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n581) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1355GAT) );
endmodule

