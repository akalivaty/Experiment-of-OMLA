

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588;

  INV_X1 U320 ( .A(KEYINPUT98), .ZN(n423) );
  XNOR2_X1 U321 ( .A(n462), .B(n461), .ZN(n468) );
  XOR2_X1 U322 ( .A(n303), .B(n302), .Z(n522) );
  XNOR2_X1 U323 ( .A(KEYINPUT109), .B(KEYINPUT47), .ZN(n461) );
  INV_X1 U324 ( .A(KEYINPUT95), .ZN(n290) );
  INV_X1 U325 ( .A(KEYINPUT117), .ZN(n473) );
  XNOR2_X1 U326 ( .A(n291), .B(n290), .ZN(n292) );
  XNOR2_X1 U327 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  XNOR2_X1 U328 ( .A(n340), .B(n292), .ZN(n293) );
  XNOR2_X1 U329 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n476) );
  OR2_X1 U331 ( .A1(n451), .A2(n581), .ZN(n452) );
  XNOR2_X1 U332 ( .A(n344), .B(n343), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n452), .B(KEYINPUT37), .ZN(n519) );
  INV_X1 U334 ( .A(G190GAT), .ZN(n480) );
  XOR2_X1 U335 ( .A(n477), .B(KEYINPUT28), .Z(n533) );
  XOR2_X1 U336 ( .A(KEYINPUT38), .B(n453), .Z(n504) );
  XNOR2_X1 U337 ( .A(n480), .B(KEYINPUT58), .ZN(n481) );
  XNOR2_X1 U338 ( .A(n454), .B(G36GAT), .ZN(n455) );
  XNOR2_X1 U339 ( .A(n482), .B(n481), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n456), .B(n455), .ZN(G1329GAT) );
  XOR2_X1 U341 ( .A(G64GAT), .B(G92GAT), .Z(n289) );
  XNOR2_X1 U342 ( .A(G176GAT), .B(G204GAT), .ZN(n288) );
  XNOR2_X1 U343 ( .A(n289), .B(n288), .ZN(n340) );
  NAND2_X1 U344 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U345 ( .A(G8GAT), .B(G183GAT), .Z(n430) );
  XOR2_X1 U346 ( .A(n293), .B(n430), .Z(n298) );
  XOR2_X1 U347 ( .A(KEYINPUT89), .B(G218GAT), .Z(n295) );
  XNOR2_X1 U348 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(G197GAT), .B(n296), .Z(n396) );
  XOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .Z(n345) );
  XNOR2_X1 U352 ( .A(n396), .B(n345), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n303) );
  XOR2_X1 U354 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n300) );
  XNOR2_X1 U355 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(n301), .ZN(n402) );
  INV_X1 U358 ( .A(n402), .ZN(n302) );
  XOR2_X1 U359 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n305) );
  XNOR2_X1 U360 ( .A(G8GAT), .B(KEYINPUT30), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n305), .B(n304), .ZN(n323) );
  XOR2_X1 U362 ( .A(G197GAT), .B(G141GAT), .Z(n307) );
  XNOR2_X1 U363 ( .A(G36GAT), .B(G50GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .Z(n309) );
  XNOR2_X1 U366 ( .A(G169GAT), .B(G22GAT), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U368 ( .A(n311), .B(n310), .Z(n321) );
  XOR2_X1 U369 ( .A(KEYINPUT65), .B(KEYINPUT68), .Z(n313) );
  XNOR2_X1 U370 ( .A(KEYINPUT67), .B(KEYINPUT70), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n319) );
  XOR2_X1 U372 ( .A(G29GAT), .B(G43GAT), .Z(n315) );
  XNOR2_X1 U373 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n349) );
  XOR2_X1 U375 ( .A(KEYINPUT69), .B(G1GAT), .Z(n431) );
  XOR2_X1 U376 ( .A(n349), .B(n431), .Z(n317) );
  NAND2_X1 U377 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n534) );
  INV_X1 U382 ( .A(n534), .ZN(n572) );
  XOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .Z(n346) );
  XOR2_X1 U384 ( .A(KEYINPUT75), .B(KEYINPUT77), .Z(n324) );
  XNOR2_X1 U385 ( .A(n346), .B(n324), .ZN(n325) );
  XOR2_X1 U386 ( .A(G120GAT), .B(G71GAT), .Z(n404) );
  XNOR2_X1 U387 ( .A(n325), .B(n404), .ZN(n329) );
  XOR2_X1 U388 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n327) );
  XNOR2_X1 U389 ( .A(KEYINPUT76), .B(KEYINPUT33), .ZN(n326) );
  XOR2_X1 U390 ( .A(n327), .B(n326), .Z(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n333) );
  INV_X1 U392 ( .A(n333), .ZN(n331) );
  NAND2_X1 U393 ( .A1(G230GAT), .A2(G233GAT), .ZN(n332) );
  INV_X1 U394 ( .A(n332), .ZN(n330) );
  NAND2_X1 U395 ( .A1(n331), .A2(n330), .ZN(n335) );
  NAND2_X1 U396 ( .A1(n333), .A2(n332), .ZN(n334) );
  NAND2_X1 U397 ( .A1(n335), .A2(n334), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n336), .B(KEYINPUT74), .ZN(n344) );
  XNOR2_X1 U399 ( .A(G106GAT), .B(G78GAT), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n337), .B(G148GAT), .ZN(n393) );
  XOR2_X1 U401 ( .A(n393), .B(KEYINPUT31), .Z(n342) );
  XOR2_X1 U402 ( .A(G57GAT), .B(KEYINPUT71), .Z(n339) );
  XNOR2_X1 U403 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n440) );
  XNOR2_X1 U405 ( .A(n440), .B(n340), .ZN(n341) );
  NOR2_X1 U406 ( .A1(n572), .A2(n457), .ZN(n490) );
  XOR2_X1 U407 ( .A(n346), .B(n345), .Z(n348) );
  XOR2_X1 U408 ( .A(G50GAT), .B(G162GAT), .Z(n386) );
  XOR2_X1 U409 ( .A(G134GAT), .B(KEYINPUT80), .Z(n370) );
  XNOR2_X1 U410 ( .A(n386), .B(n370), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U412 ( .A(n349), .B(KEYINPUT9), .Z(n351) );
  NAND2_X1 U413 ( .A1(G232GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U415 ( .A(n353), .B(n352), .Z(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n355) );
  XNOR2_X1 U417 ( .A(G218GAT), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT64), .Z(n357) );
  XNOR2_X1 U420 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U423 ( .A(n361), .B(n360), .Z(n543) );
  XNOR2_X1 U424 ( .A(n543), .B(KEYINPUT36), .ZN(n584) );
  XOR2_X1 U425 ( .A(KEYINPUT4), .B(G57GAT), .Z(n363) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G120GAT), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U428 ( .A(G155GAT), .B(G162GAT), .Z(n365) );
  XNOR2_X1 U429 ( .A(G127GAT), .B(G148GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n383) );
  XOR2_X1 U432 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n369) );
  XNOR2_X1 U433 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U435 ( .A(G85GAT), .B(n370), .Z(n372) );
  XOR2_X1 U436 ( .A(G113GAT), .B(KEYINPUT0), .Z(n403) );
  XNOR2_X1 U437 ( .A(G29GAT), .B(n403), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U439 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n377), .B(KEYINPUT5), .Z(n381) );
  XOR2_X1 U443 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n379) );
  XNOR2_X1 U444 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n395) );
  XNOR2_X1 U446 ( .A(n395), .B(KEYINPUT6), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n520) );
  XOR2_X1 U449 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n385) );
  XNOR2_X1 U450 ( .A(KEYINPUT23), .B(KEYINPUT88), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U452 ( .A(KEYINPUT22), .B(G204GAT), .Z(n388) );
  XOR2_X1 U453 ( .A(G22GAT), .B(G155GAT), .Z(n442) );
  XNOR2_X1 U454 ( .A(n386), .B(n442), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U456 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U457 ( .A1(G228GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U459 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n477) );
  XOR2_X1 U462 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n400) );
  XNOR2_X1 U463 ( .A(G43GAT), .B(G99GAT), .ZN(n399) );
  XNOR2_X1 U464 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U465 ( .A(n402), .B(n401), .Z(n414) );
  XOR2_X1 U466 ( .A(G190GAT), .B(G134GAT), .Z(n406) );
  XNOR2_X1 U467 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U469 ( .A(G15GAT), .B(G127GAT), .Z(n443) );
  XOR2_X1 U470 ( .A(n407), .B(n443), .Z(n412) );
  XOR2_X1 U471 ( .A(G176GAT), .B(G183GAT), .Z(n409) );
  NAND2_X1 U472 ( .A1(G227GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U474 ( .A(KEYINPUT85), .B(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U476 ( .A(n414), .B(n413), .ZN(n531) );
  NAND2_X1 U477 ( .A1(n531), .A2(n522), .ZN(n415) );
  XOR2_X1 U478 ( .A(KEYINPUT97), .B(n415), .Z(n416) );
  NAND2_X1 U479 ( .A1(n477), .A2(n416), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n417), .B(KEYINPUT25), .ZN(n421) );
  XOR2_X1 U481 ( .A(n522), .B(KEYINPUT96), .Z(n418) );
  XOR2_X1 U482 ( .A(KEYINPUT27), .B(n418), .Z(n425) );
  NOR2_X1 U483 ( .A1(n531), .A2(n477), .ZN(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT26), .B(n419), .ZN(n570) );
  AND2_X1 U485 ( .A1(n425), .A2(n570), .ZN(n420) );
  NOR2_X1 U486 ( .A1(n421), .A2(n420), .ZN(n422) );
  NOR2_X1 U487 ( .A1(n520), .A2(n422), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n429) );
  NAND2_X1 U489 ( .A1(n520), .A2(n425), .ZN(n529) );
  NOR2_X1 U490 ( .A1(n531), .A2(n529), .ZN(n427) );
  INV_X1 U491 ( .A(n533), .ZN(n426) );
  NAND2_X1 U492 ( .A1(n427), .A2(n426), .ZN(n428) );
  NAND2_X1 U493 ( .A1(n429), .A2(n428), .ZN(n488) );
  NAND2_X1 U494 ( .A1(n584), .A2(n488), .ZN(n451) );
  XOR2_X1 U495 ( .A(n430), .B(G78GAT), .Z(n433) );
  XNOR2_X1 U496 ( .A(n431), .B(G211GAT), .ZN(n432) );
  XNOR2_X1 U497 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U498 ( .A(n434), .B(G64GAT), .Z(n439) );
  XOR2_X1 U499 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n436) );
  XNOR2_X1 U500 ( .A(KEYINPUT15), .B(KEYINPUT82), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U502 ( .A(G71GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U504 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n450) );
  XOR2_X1 U507 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n447) );
  NAND2_X1 U508 ( .A1(G231GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U509 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U510 ( .A(KEYINPUT81), .B(n448), .Z(n449) );
  XOR2_X1 U511 ( .A(n450), .B(n449), .Z(n554) );
  INV_X1 U512 ( .A(n554), .ZN(n581) );
  NAND2_X1 U513 ( .A1(n490), .A2(n519), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n522), .A2(n504), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n454) );
  INV_X1 U516 ( .A(n543), .ZN(n557) );
  XOR2_X1 U517 ( .A(KEYINPUT41), .B(n457), .Z(n536) );
  AND2_X1 U518 ( .A1(n536), .A2(n534), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT46), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n581), .A2(n459), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n460), .A2(n557), .ZN(n462) );
  NAND2_X1 U522 ( .A1(n581), .A2(n584), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n463), .B(KEYINPUT110), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n464), .B(KEYINPUT45), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n465), .A2(n457), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n572), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n470) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n530) );
  INV_X1 U530 ( .A(n530), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT116), .B(n522), .ZN(n471) );
  NAND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n520), .A2(n476), .ZN(n571) );
  NAND2_X1 U534 ( .A1(n477), .A2(n571), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n479), .A2(n531), .ZN(n563) );
  NOR2_X1 U537 ( .A1(n557), .A2(n563), .ZN(n482) );
  INV_X1 U538 ( .A(G183GAT), .ZN(n485) );
  NOR2_X1 U539 ( .A1(n563), .A2(n554), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT122), .B(n483), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1350GAT) );
  NAND2_X1 U542 ( .A1(n557), .A2(n581), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  NAND2_X1 U544 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n489), .B(KEYINPUT99), .ZN(n507) );
  AND2_X1 U546 ( .A1(n490), .A2(n507), .ZN(n496) );
  NAND2_X1 U547 ( .A1(n520), .A2(n496), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(n491), .ZN(n492) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n496), .A2(n522), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U553 ( .A1(n496), .A2(n531), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U555 ( .A1(n496), .A2(n533), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(KEYINPUT100), .ZN(n498) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n498), .ZN(G1327GAT) );
  NAND2_X1 U558 ( .A1(n504), .A2(n520), .ZN(n501) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT101), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n531), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n533), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  INV_X1 U568 ( .A(n536), .ZN(n564) );
  NOR2_X1 U569 ( .A1(n564), .A2(n534), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT104), .ZN(n518) );
  AND2_X1 U571 ( .A1(n507), .A2(n518), .ZN(n514) );
  NAND2_X1 U572 ( .A1(n520), .A2(n514), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT105), .Z(n511) );
  NAND2_X1 U575 ( .A1(n514), .A2(n522), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n514), .A2(n531), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n533), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  AND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n526), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT108), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n524), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n526), .A2(n531), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n526), .A2(n533), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n548) );
  NAND2_X1 U596 ( .A1(n531), .A2(n548), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n533), .A2(n532), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n544), .A2(n534), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U601 ( .A1(n544), .A2(n536), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n541) );
  NAND2_X1 U605 ( .A1(n544), .A2(n581), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n570), .ZN(n556) );
  NOR2_X1 U613 ( .A1(n572), .A2(n556), .ZN(n549) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n549), .Z(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT114), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n564), .A2(n556), .ZN(n552) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n554), .A2(n556), .ZN(n555) );
  XOR2_X1 U621 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n559) );
  XNOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT115), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n562) );
  NOR2_X1 U626 ( .A1(n563), .A2(n572), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(KEYINPUT119), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n566) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n571), .A2(n570), .ZN(n578) );
  NOR2_X1 U636 ( .A1(n572), .A2(n578), .ZN(n577) );
  XOR2_X1 U637 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT123), .B(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n578), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n457), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n587) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

