//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n211), .A2(G20), .A3(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n206), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT65), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT66), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT76), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(new_n216), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G58), .A2(G68), .ZN(new_n250));
  OAI21_X1  g0050(.A(G20), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G159), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(KEYINPUT16), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT75), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n204), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT7), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT7), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n257), .A2(new_n261), .A3(new_n204), .A4(new_n258), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n216), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n255), .B1(new_n263), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n212), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n260), .A2(G68), .A3(new_n262), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n251), .A2(new_n253), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT16), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n247), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n273), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n275), .A2(new_n267), .A3(KEYINPUT76), .A4(new_n269), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(G274), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G232), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT78), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G87), .ZN(new_n288));
  OR2_X1    g0088(.A1(G223), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n288), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT78), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n283), .A2(new_n285), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n287), .A2(new_n298), .A3(new_n299), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n257), .A2(new_n258), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(new_n289), .A3(new_n291), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n282), .B1(new_n305), .B2(new_n288), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n306), .B2(new_n286), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT79), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n307), .A3(KEYINPUT79), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT80), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n269), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n203), .A2(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n317), .A2(new_n321), .B1(new_n319), .B2(new_n314), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n277), .A2(new_n312), .A3(new_n313), .A4(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT17), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n322), .B1(new_n274), .B2(new_n276), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n327), .A2(new_n313), .A3(KEYINPUT17), .A4(new_n312), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n269), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n261), .B1(new_n295), .B2(new_n204), .ZN(new_n331));
  NOR4_X1   g0131(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT7), .A4(G20), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT75), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n265), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n334), .B2(new_n255), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT76), .B1(new_n335), .B2(new_n275), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n254), .B1(new_n333), .B2(new_n265), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n337), .A2(new_n273), .A3(new_n247), .A4(new_n330), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n323), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT77), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n327), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(G179), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n287), .A2(new_n298), .A3(new_n343), .A4(new_n301), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n306), .B2(new_n286), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n340), .A2(new_n342), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n329), .B1(KEYINPUT18), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n340), .A2(new_n342), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n204), .A2(G33), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n222), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(new_n269), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n356), .A2(KEYINPUT11), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n315), .A2(new_n216), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT12), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(KEYINPUT11), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n316), .A2(G68), .A3(new_n320), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n357), .A2(new_n359), .A3(new_n360), .A4(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(G232), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  OAI211_X1 g0164(.A(G226), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n365));
  INV_X1    g0165(.A(G33), .ZN(new_n366));
  INV_X1    g0166(.A(G97), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n363), .B(new_n365), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n297), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT13), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n282), .A2(new_n284), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G274), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n373), .B1(new_n213), .B2(new_n281), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n372), .A2(G238), .B1(new_n374), .B2(new_n280), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n370), .B1(new_n369), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT74), .B1(new_n378), .B2(G179), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .A4(new_n343), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(KEYINPUT73), .A2(G169), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT14), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT14), .ZN(new_n385));
  INV_X1    g0185(.A(new_n383), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(new_n376), .C2(new_n377), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n362), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n283), .B1(new_n290), .B2(new_n371), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n304), .A2(G222), .A3(new_n364), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n304), .A2(G1698), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT67), .B(G223), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n391), .B1(new_n222), .B2(new_n304), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n394), .B2(new_n297), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n395), .A2(KEYINPUT72), .A3(G190), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT72), .B1(new_n395), .B2(G190), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G150), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n204), .A2(new_n366), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n318), .A2(new_n354), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G50), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n204), .B1(new_n250), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n269), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n402), .B1(new_n203), .B2(G20), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n316), .A2(new_n405), .B1(new_n402), .B2(new_n315), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT9), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT9), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n409), .A3(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n303), .B2(new_n395), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT10), .B1(new_n398), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n394), .A2(new_n297), .ZN(new_n414));
  INV_X1    g0214(.A(new_n390), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(G200), .B1(new_n408), .B2(new_n410), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n397), .C2(new_n396), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n416), .A2(G179), .ZN(new_n421));
  OR2_X1    g0221(.A1(new_n421), .A2(KEYINPUT69), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n407), .B1(new_n395), .B2(G169), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT68), .ZN(new_n424));
  OR2_X1    g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(KEYINPUT69), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n422), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n319), .A2(KEYINPUT71), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT71), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n318), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n400), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n433), .A2(new_n354), .B1(new_n204), .B2(new_n222), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n269), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n320), .A2(G77), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n316), .A2(new_n437), .B1(new_n222), .B2(new_n315), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n283), .B1(new_n223), .B2(new_n371), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n304), .A2(G232), .A3(new_n364), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT70), .A2(G107), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT70), .A2(G107), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(new_n295), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n441), .B(new_n445), .C1(new_n392), .C2(new_n217), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n440), .B1(new_n446), .B2(new_n297), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n439), .B1(G169), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n343), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n435), .B(new_n438), .C1(new_n447), .C2(new_n303), .ZN(new_n451));
  INV_X1    g0251(.A(new_n447), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n299), .ZN(new_n453));
  OAI22_X1  g0253(.A1(new_n448), .A2(new_n450), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g0254(.A(G200), .B1(new_n376), .B2(new_n377), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n362), .B1(new_n378), .B2(G190), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n389), .A2(new_n420), .A3(new_n428), .A4(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n350), .A2(new_n352), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT90), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n204), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n462), .A2(KEYINPUT87), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n304), .A2(new_n204), .A3(G87), .A4(new_n463), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G116), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT88), .B1(new_n469), .B2(G20), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT88), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(new_n204), .A3(G33), .A4(G116), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n468), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n442), .A2(G20), .A3(new_n443), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n475));
  NOR2_X1   g0275(.A1(KEYINPUT89), .A2(KEYINPUT23), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT24), .B1(new_n467), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n473), .A2(new_n478), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT24), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n465), .A2(new_n466), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n330), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n314), .B2(G107), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n314), .A2(new_n486), .A3(G107), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n203), .A2(G33), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n314), .A2(new_n490), .A3(new_n212), .A4(new_n268), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n488), .A2(new_n489), .B1(new_n224), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n460), .B1(new_n485), .B2(new_n492), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n467), .A2(KEYINPUT24), .A3(new_n479), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n269), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n492), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(KEYINPUT90), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n279), .A2(G1), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n374), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n499), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n282), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n503), .B2(new_n225), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n304), .A2(G257), .A3(G1698), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n304), .A2(G250), .A3(new_n364), .ZN(new_n506));
  INV_X1    g0306(.A(G294), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n506), .C1(new_n366), .C2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n504), .B1(new_n297), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G179), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n345), .B2(new_n509), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n493), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(G190), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n496), .A3(new_n497), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n502), .A2(G270), .A3(new_n282), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n501), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n304), .A2(G264), .A3(G1698), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n304), .A2(G257), .A3(new_n364), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n295), .A2(G303), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n297), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n345), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G283), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n204), .C1(G33), .C2(new_n367), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n269), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n491), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(KEYINPUT85), .A3(G116), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n491), .B2(new_n530), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n314), .A2(G116), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT86), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n534), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n527), .A2(new_n542), .A3(KEYINPUT21), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n520), .B1(new_n297), .B2(new_n525), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n544), .A3(G179), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT21), .B1(new_n527), .B2(new_n542), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n521), .A2(new_n526), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n542), .B1(G200), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n299), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT82), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT81), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n400), .B2(new_n222), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n252), .A2(KEYINPUT81), .A3(G77), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  AND2_X1   g0359(.A1(G97), .A2(G107), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G97), .A2(G107), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n558), .B1(G20), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n260), .A2(new_n262), .A3(new_n444), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n330), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n314), .A2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n535), .B2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n554), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n564), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(new_n558), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n566), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n269), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(KEYINPUT82), .A3(new_n569), .ZN(new_n576));
  AND2_X1   g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n502), .A2(G257), .A3(new_n282), .ZN(new_n578));
  OAI211_X1 g0378(.A(G244), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n304), .A2(KEYINPUT4), .A3(G244), .A4(new_n364), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n304), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n528), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n578), .B1(new_n584), .B2(new_n297), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(new_n299), .A3(new_n501), .ZN(new_n586));
  INV_X1    g0386(.A(new_n501), .ZN(new_n587));
  AOI211_X1 g0387(.A(new_n587), .B(new_n578), .C1(new_n584), .C2(new_n297), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n588), .B2(G200), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(G179), .A3(new_n501), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n588), .B2(new_n345), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n575), .A2(new_n569), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n577), .A2(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n354), .A2(KEYINPUT19), .A3(new_n367), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G87), .A2(G97), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n442), .A2(new_n595), .A3(new_n443), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n204), .B1(new_n366), .B2(new_n367), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n594), .B1(new_n598), .B2(KEYINPUT19), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n204), .B(G68), .C1(new_n293), .C2(new_n294), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT83), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n304), .A2(KEYINPUT83), .A3(new_n204), .A4(G68), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n269), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n433), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n314), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n535), .A2(new_n606), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n605), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  OAI211_X1 g0410(.A(G238), .B(new_n364), .C1(new_n293), .C2(new_n294), .ZN(new_n611));
  OAI211_X1 g0411(.A(G244), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n612), .A3(new_n469), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n297), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n499), .A2(new_n219), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n374), .A2(new_n499), .B1(new_n615), .B2(new_n282), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n343), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n616), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n345), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n610), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT19), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n596), .B2(new_n597), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n602), .B(new_n603), .C1(new_n623), .C2(new_n594), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n607), .B1(new_n624), .B2(new_n269), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n619), .A2(G200), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n614), .A2(G190), .A3(new_n616), .ZN(new_n627));
  OR3_X1    g0427(.A1(new_n491), .A2(KEYINPUT84), .A3(new_n218), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT84), .B1(new_n491), .B2(new_n218), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n625), .A2(new_n626), .A3(new_n627), .A4(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n621), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n593), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n459), .A2(new_n518), .A3(new_n553), .A4(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n428), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT18), .B1(new_n327), .B2(new_n347), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n339), .A2(new_n351), .A3(new_n348), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n452), .A2(new_n345), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(new_n449), .A3(new_n439), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n640), .A2(KEYINPUT93), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(KEYINPUT93), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n456), .A2(new_n455), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n384), .B(new_n387), .C1(new_n379), .C2(new_n381), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n644), .A2(new_n645), .B1(new_n362), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n638), .B1(new_n647), .B2(new_n329), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n635), .B1(new_n648), .B2(new_n420), .ZN(new_n649));
  INV_X1    g0449(.A(new_n459), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n610), .A2(new_n618), .A3(new_n620), .ZN(new_n651));
  INV_X1    g0451(.A(new_n627), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT91), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n625), .A2(new_n626), .A3(KEYINPUT91), .A4(new_n630), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n651), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n593), .A2(new_n657), .A3(new_n516), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n496), .A2(new_n497), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n511), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n547), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n545), .A3(new_n543), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n621), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n584), .A2(new_n297), .ZN(new_n665));
  INV_X1    g0465(.A(new_n578), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n501), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G169), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n668), .A2(new_n590), .B1(new_n571), .B2(new_n576), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT26), .B1(new_n657), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n591), .A2(new_n631), .A3(new_n621), .A4(new_n592), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n664), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n649), .B1(new_n650), .B2(new_n676), .ZN(G369));
  NAND3_X1  g0477(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(G213), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n493), .A2(new_n498), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n518), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n512), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n683), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT94), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n548), .B2(new_n683), .ZN(new_n689));
  INV_X1    g0489(.A(new_n683), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n662), .A2(KEYINPUT94), .A3(new_n690), .ZN(new_n691));
  AOI22_X1  g0491(.A1(new_n685), .A2(new_n687), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n660), .A2(new_n690), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n542), .A2(new_n683), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n662), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n552), .B2(new_n696), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n687), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n695), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n207), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n596), .A2(G116), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n210), .B2(new_n706), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n710));
  XNOR2_X1  g0510(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n509), .A2(new_n617), .A3(new_n585), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n544), .A2(G179), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n508), .A2(new_n297), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n716), .A2(new_n504), .A3(new_n619), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n549), .A2(new_n343), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n544), .A2(new_n617), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n513), .A3(new_n343), .A4(new_n667), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n715), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n683), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT31), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n633), .A2(new_n518), .A3(new_n553), .A4(new_n690), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n690), .B1(new_n664), .B2(new_n674), .ZN(new_n730));
  XNOR2_X1  g0530(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n605), .A2(new_n608), .A3(new_n630), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n303), .B1(new_n614), .B2(new_n616), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n654), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(new_n627), .A3(new_n656), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n669), .A3(KEYINPUT26), .A4(new_n621), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n671), .A2(new_n672), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n512), .A2(new_n548), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n621), .C1(new_n658), .C2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT29), .A3(new_n690), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n729), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n711), .B1(new_n745), .B2(G1), .ZN(G364));
  INV_X1    g0546(.A(G13), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n203), .B1(new_n748), .B2(G45), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n706), .A2(KEYINPUT97), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT97), .ZN(new_n751));
  INV_X1    g0551(.A(new_n749), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n705), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n207), .A2(new_n304), .ZN(new_n756));
  INV_X1    g0556(.A(G355), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n756), .A2(new_n757), .B1(G116), .B2(new_n207), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n704), .A2(new_n304), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(new_n211), .B2(new_n279), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n245), .A2(G45), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n212), .B1(G20), .B2(new_n345), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n755), .B1(new_n763), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n204), .B1(new_n771), .B2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n367), .ZN(new_n773));
  NAND3_X1  g0573(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n299), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n402), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(G190), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n773), .B(new_n777), .C1(G68), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n204), .A2(new_n299), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n343), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n304), .B1(new_n782), .B2(new_n248), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n204), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n781), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(G77), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n784), .A2(new_n771), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT98), .B(KEYINPUT32), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OR3_X1    g0592(.A1(new_n303), .A2(KEYINPUT99), .A3(G179), .ZN(new_n793));
  OAI21_X1  g0593(.A(KEYINPUT99), .B1(new_n303), .B2(G179), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n793), .A2(new_n780), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n793), .A2(new_n784), .A3(new_n794), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G87), .A2(new_n796), .B1(new_n798), .B2(G107), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n779), .A2(new_n787), .A3(new_n792), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n295), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT100), .Z(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n782), .A2(new_n804), .B1(new_n785), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n797), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n788), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n806), .B(new_n808), .C1(G329), .C2(new_n809), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT33), .B(G317), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n778), .ZN(new_n812));
  INV_X1    g0612(.A(new_n772), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G294), .B1(G326), .B2(new_n775), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n810), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n800), .B1(new_n803), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n770), .B1(new_n816), .B2(new_n767), .ZN(new_n817));
  INV_X1    g0617(.A(new_n766), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n698), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n699), .A2(new_n754), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n698), .A2(G330), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n439), .A2(new_n683), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n640), .B(new_n823), .C1(new_n453), .C2(new_n451), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n643), .B2(new_n823), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n730), .B(new_n825), .Z(new_n826));
  AOI21_X1  g0626(.A(new_n755), .B1(new_n826), .B2(new_n729), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n729), .B2(new_n826), .ZN(new_n828));
  INV_X1    g0628(.A(new_n767), .ZN(new_n829));
  INV_X1    g0629(.A(new_n782), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G143), .A2(new_n830), .B1(new_n786), .B2(G159), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n775), .A2(G137), .ZN(new_n832));
  INV_X1    g0632(.A(new_n778), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n832), .C1(new_n399), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT34), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n835), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n797), .A2(new_n216), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n304), .B1(new_n772), .B2(new_n248), .C1(new_n840), .C2(new_n788), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G50), .B2(new_n796), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n836), .A2(new_n837), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n295), .B1(new_n788), .B2(new_n805), .C1(new_n507), .C2(new_n782), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n773), .B(new_n844), .C1(G303), .C2(new_n775), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n798), .A2(G87), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n796), .A2(G107), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n833), .A2(new_n807), .B1(new_n785), .B2(new_n530), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n845), .A2(new_n846), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n829), .B1(new_n843), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n767), .A2(new_n764), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n754), .B(new_n851), .C1(new_n222), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n825), .B2(new_n765), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n828), .A2(new_n854), .ZN(G384));
  NOR2_X1   g0655(.A1(new_n748), .A2(new_n203), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT103), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n389), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n646), .A2(KEYINPUT103), .A3(new_n362), .ZN(new_n860));
  INV_X1    g0660(.A(new_n645), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n362), .A2(new_n683), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n861), .B2(new_n646), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT31), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT105), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n722), .A2(new_n683), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n868), .B1(new_n722), .B2(new_n683), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n725), .A2(new_n871), .ZN(new_n872));
  AND4_X1   g0672(.A1(new_n857), .A2(new_n866), .A3(new_n825), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(new_n681), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n340), .A2(new_n342), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n327), .B2(new_n312), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n349), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n272), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n333), .B2(new_n265), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n880), .A2(KEYINPUT104), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT16), .B1(new_n880), .B2(KEYINPUT104), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n270), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n875), .B1(new_n883), .B2(new_n322), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n348), .B1(new_n883), .B2(new_n322), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n327), .A2(new_n312), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n326), .A2(new_n328), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n349), .A2(KEYINPUT18), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n890), .A3(new_n352), .ZN(new_n891));
  INV_X1    g0691(.A(new_n884), .ZN(new_n892));
  AOI221_X4 g0692(.A(new_n874), .B1(new_n878), .B2(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n878), .A2(new_n888), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n873), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n866), .A2(new_n825), .A3(new_n872), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n326), .A2(new_n328), .A3(new_n636), .A4(new_n637), .ZN(new_n900));
  INV_X1    g0700(.A(new_n876), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n349), .A2(new_n876), .A3(new_n877), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n339), .A2(new_n348), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n886), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n904), .B1(new_n906), .B2(new_n876), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n874), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n898), .B1(new_n899), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n897), .B1(new_n857), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n872), .A2(new_n352), .A3(new_n350), .A4(new_n458), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(G330), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(KEYINPUT106), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(KEYINPUT106), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n894), .A2(new_n895), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n874), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n899), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n905), .A2(new_n886), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n878), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n923), .B2(new_n902), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n920), .B1(new_n893), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n683), .B1(new_n859), .B2(new_n860), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n638), .A2(new_n875), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n893), .A2(new_n896), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n690), .B(new_n825), .C1(new_n664), .C2(new_n674), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n640), .A2(new_n683), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n866), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n459), .A2(new_n732), .A3(new_n742), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n649), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n935), .B(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n856), .B1(new_n916), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n938), .B2(new_n916), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n212), .A2(new_n204), .A3(new_n530), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n564), .B(KEYINPUT102), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT35), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n944), .B2(new_n943), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT36), .Z(new_n947));
  NOR3_X1   g0747(.A1(new_n249), .A2(new_n210), .A3(new_n222), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n216), .A2(G50), .ZN(new_n949));
  OAI211_X1 g0749(.A(G1), .B(new_n747), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n591), .A2(new_n592), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n593), .B1(new_n577), .B2(new_n690), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n669), .A2(new_n683), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n952), .B1(new_n956), .B2(new_n512), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n690), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n692), .A2(KEYINPUT42), .A3(new_n955), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT42), .B1(new_n692), .B2(new_n955), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n733), .A2(new_n683), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n621), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n657), .B2(new_n963), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT108), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n692), .A2(new_n955), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT42), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n959), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT108), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n966), .A2(new_n967), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n958), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n969), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n962), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n702), .A2(new_n956), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n977), .A2(KEYINPUT109), .A3(new_n979), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n983), .ZN(new_n986));
  AOI221_X4 g0786(.A(new_n981), .B1(new_n962), .B2(new_n978), .C1(new_n969), .C2(new_n976), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT109), .B1(new_n977), .B2(new_n979), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n705), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n695), .B2(new_n955), .ZN(new_n992));
  OAI211_X1 g0792(.A(KEYINPUT44), .B(new_n956), .C1(new_n692), .C2(new_n694), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n689), .A2(new_n691), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n701), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n693), .A3(new_n955), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n994), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n700), .A3(new_n701), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n699), .A2(new_n685), .A3(new_n687), .ZN(new_n1004));
  AND4_X1   g0804(.A1(new_n702), .A2(new_n689), .A3(new_n691), .A4(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n702), .A2(new_n1004), .B1(new_n689), .B2(new_n691), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(new_n744), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n994), .A2(new_n1001), .A3(new_n702), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1003), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n990), .B1(new_n1010), .B2(new_n745), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n985), .B(new_n989), .C1(new_n752), .C2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n768), .B1(new_n207), .B2(new_n433), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n233), .B2(new_n759), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n782), .A2(new_n399), .B1(new_n785), .B2(new_n402), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n295), .B(new_n1016), .C1(G137), .C2(new_n809), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n772), .A2(new_n216), .ZN(new_n1018));
  INV_X1    g0818(.A(G143), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n776), .A2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1018), .B(new_n1020), .C1(G159), .C2(new_n778), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n796), .A2(G58), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n798), .A2(G77), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G317), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n782), .A2(new_n801), .B1(new_n788), .B2(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n304), .B(new_n1026), .C1(G283), .C2(new_n786), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n778), .A2(G294), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n813), .A2(new_n444), .B1(G311), .B2(new_n775), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n798), .A2(G97), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n795), .A2(new_n530), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT46), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n754), .B(new_n1015), .C1(new_n1035), .C2(new_n767), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n818), .B2(new_n966), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT111), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1012), .A2(new_n1038), .ZN(G387));
  INV_X1    g0839(.A(new_n1007), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n685), .A2(new_n687), .A3(new_n766), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n756), .A2(new_n707), .B1(G107), .B2(new_n207), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n429), .A2(new_n431), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n402), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT50), .Z(new_n1045));
  OAI211_X1 g0845(.A(new_n707), .B(new_n279), .C1(new_n216), .C2(new_n222), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT112), .Z(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n760), .B1(new_n237), .B2(G45), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1042), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n755), .B1(new_n1050), .B2(new_n769), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n782), .A2(new_n402), .B1(new_n788), .B2(new_n399), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n295), .B(new_n1052), .C1(G68), .C2(new_n786), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n789), .A2(new_n776), .B1(new_n833), .B2(new_n318), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n772), .A2(new_n433), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n796), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1053), .A2(new_n1030), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n782), .A2(new_n1025), .B1(new_n785), .B2(new_n801), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(KEYINPUT113), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n778), .A2(G311), .B1(new_n775), .B2(G322), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT48), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n795), .A2(new_n507), .B1(new_n807), .B2(new_n772), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n304), .B1(new_n809), .B2(G326), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n530), .C2(new_n797), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT49), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1058), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1051), .B1(new_n1072), .B2(new_n767), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1040), .A2(new_n752), .B1(new_n1041), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1008), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n705), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1040), .A2(new_n745), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  INV_X1    g0878(.A(KEYINPUT114), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1003), .A2(new_n1079), .A3(new_n1009), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n994), .A2(new_n1001), .A3(new_n702), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(KEYINPUT114), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1075), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n702), .B1(new_n994), .B2(new_n1001), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n706), .B1(new_n1085), .B2(new_n1008), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n752), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n242), .A2(new_n760), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n768), .B1(new_n367), .B2(new_n207), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n755), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n295), .B1(new_n785), .B2(new_n507), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n833), .A2(new_n801), .B1(new_n772), .B2(new_n530), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G322), .C2(new_n809), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n1095), .B1(new_n224), .B2(new_n797), .C1(new_n807), .C2(new_n795), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n830), .A2(G311), .B1(G317), .B2(new_n775), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n830), .A2(G159), .B1(G150), .B2(new_n775), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n772), .A2(new_n222), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n304), .B1(new_n788), .B2(new_n1019), .C1(new_n833), .C2(new_n402), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(KEYINPUT51), .B2(new_n1099), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1043), .A2(new_n786), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1105), .B(new_n846), .C1(new_n216), .C2(new_n795), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1096), .A2(new_n1098), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1107), .B2(new_n767), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n955), .B2(new_n818), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1087), .A2(new_n1089), .A3(new_n1109), .ZN(G390));
  NAND3_X1  g0910(.A1(new_n872), .A2(G330), .A3(new_n825), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n866), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n926), .B1(new_n933), .B2(new_n866), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n919), .B2(new_n925), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n741), .A2(new_n690), .A3(new_n825), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n932), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n866), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n926), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1118), .B(new_n1119), .C1(new_n893), .C2(new_n924), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1113), .B1(new_n1115), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT116), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n912), .B2(new_n727), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n459), .A2(KEYINPUT116), .A3(G330), .A4(new_n872), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n936), .A4(new_n649), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n825), .A2(G330), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n724), .B2(new_n725), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n866), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n933), .B1(new_n1113), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n866), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n932), .A4(new_n1116), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT115), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1114), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n893), .A2(new_n896), .A3(new_n920), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT39), .B1(new_n899), .B2(new_n909), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1120), .A2(new_n1133), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1138), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1120), .A2(new_n1133), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1115), .A2(new_n1145), .A3(KEYINPUT115), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1122), .B(new_n1137), .C1(new_n1144), .C2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1136), .B(KEYINPUT117), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1142), .A2(new_n1143), .A3(new_n1138), .ZN(new_n1149));
  OAI21_X1  g0949(.A(KEYINPUT115), .B1(new_n1115), .B2(new_n1145), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1142), .A2(new_n1120), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1149), .A2(new_n1150), .B1(new_n1151), .B2(new_n1113), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1147), .B(new_n705), .C1(new_n1148), .C2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1141), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(new_n765), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n852), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n304), .B1(new_n809), .B2(G294), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n367), .B2(new_n785), .C1(new_n530), .C2(new_n782), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n838), .B(new_n1158), .C1(G87), .C2(new_n796), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n776), .A2(new_n807), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1101), .B(new_n1160), .C1(new_n444), .C2(new_n778), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n813), .A2(G159), .B1(G137), .B2(new_n778), .ZN(new_n1162));
  INV_X1    g0962(.A(G128), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1162), .B1(new_n1163), .B2(new_n776), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n797), .A2(new_n402), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n304), .B1(new_n785), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(G125), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n782), .A2(new_n840), .B1(new_n788), .B2(new_n1168), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n795), .A2(new_n399), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT53), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1159), .A2(new_n1161), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n755), .B1(new_n319), .B2(new_n1156), .C1(new_n1173), .C2(new_n829), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(new_n1152), .B2(new_n752), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1153), .A2(new_n1176), .ZN(G378));
  AND2_X1   g0977(.A1(new_n420), .A2(new_n428), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n407), .A2(new_n875), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1178), .B(new_n1179), .Z(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n899), .A2(new_n909), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n898), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n857), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n866), .A2(new_n872), .A3(new_n857), .A4(new_n825), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n918), .B2(new_n899), .ZN(new_n1187));
  OAI211_X1 g0987(.A(G330), .B(new_n1182), .C1(new_n1185), .C2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1182), .B1(new_n911), .B2(G330), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n935), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(G330), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1182), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n928), .B1(new_n929), .B2(new_n934), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1154), .B2(new_n926), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1196), .A3(new_n1188), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1191), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT57), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1126), .B1(new_n1152), .B2(new_n1137), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n705), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1147), .A2(new_n1127), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1198), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1193), .A2(new_n764), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n304), .A2(G41), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n402), .B1(G33), .B2(G41), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n782), .A2(new_n224), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT118), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1208), .B1(new_n807), .B2(new_n788), .C1(new_n433), .C2(new_n785), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1018), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n833), .A2(new_n367), .B1(new_n776), .B2(new_n530), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(KEYINPUT118), .B2(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n798), .A2(G58), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1057), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1210), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1166), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n796), .A2(new_n1223), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G128), .A2(new_n830), .B1(new_n786), .B2(G137), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n778), .A2(G132), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n813), .A2(G150), .B1(G125), .B2(new_n775), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n798), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n767), .B1(new_n1222), .B2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT119), .Z(new_n1236));
  AOI211_X1 g1036(.A(new_n754), .B(new_n1236), .C1(new_n402), .C2(new_n852), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1198), .A2(new_n752), .B1(new_n1207), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1206), .A2(new_n1238), .ZN(G375));
  INV_X1    g1039(.A(new_n1148), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n990), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(new_n1135), .C2(new_n1127), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n444), .A2(new_n786), .B1(new_n809), .B2(G303), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n304), .B1(new_n830), .B2(G283), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1023), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1055), .B1(new_n778), .B2(G116), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n507), .B2(new_n776), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1245), .B(new_n1247), .C1(G97), .C2(new_n796), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(KEYINPUT120), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n795), .A2(new_n789), .B1(new_n1163), .B2(new_n788), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT121), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n776), .A2(new_n840), .B1(new_n772), .B2(new_n402), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n778), .B2(new_n1223), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n304), .B1(new_n785), .B2(new_n399), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G137), .B2(new_n830), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1252), .A2(new_n1218), .A3(new_n1254), .A4(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT120), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1248), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n767), .B1(new_n1250), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1260), .B(new_n755), .C1(G68), .C2(new_n1156), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1112), .B2(new_n764), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1135), .B2(new_n752), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1242), .A2(new_n1263), .ZN(G381));
  NOR4_X1   g1064(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1263), .A3(new_n1242), .ZN(new_n1266));
  OR4_X1    g1066(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1266), .ZN(G407));
  AND2_X1   g1067(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n682), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G407), .B(G213), .C1(G375), .C2(new_n1271), .ZN(G409));
  OAI211_X1 g1072(.A(G378), .B(new_n1238), .C1(new_n1201), .C2(new_n1204), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n990), .B1(new_n1191), .B2(new_n1197), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT122), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1203), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1203), .B2(new_n1274), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1198), .A2(new_n752), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1207), .A2(new_n1237), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1276), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1273), .B1(new_n1281), .B2(G378), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1269), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT123), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1285), .A2(new_n1286), .A3(KEYINPUT60), .A4(new_n1126), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1126), .A2(KEYINPUT60), .A3(new_n1131), .A4(new_n1134), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT123), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT60), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n706), .B1(new_n1127), .B2(new_n1135), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1287), .A2(new_n1289), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1293), .A2(G384), .A3(new_n1263), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1293), .B2(new_n1263), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1284), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1263), .ZN(new_n1297));
  INV_X1    g1097(.A(G384), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1293), .A2(G384), .A3(new_n1263), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(KEYINPUT124), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1270), .A2(G2897), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(G2897), .A3(new_n1270), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1283), .A2(KEYINPUT126), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1198), .A2(new_n1241), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT122), .B1(new_n1311), .B2(new_n1200), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1203), .A2(new_n1274), .A3(new_n1275), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1312), .A2(new_n1238), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1268), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1270), .B1(new_n1315), .B2(new_n1273), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1310), .B1(new_n1316), .B2(new_n1307), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1309), .A2(new_n1317), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1012), .A2(G390), .A3(new_n1038), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G390), .B1(new_n1012), .B2(new_n1038), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT127), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(G393), .B(G396), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT61), .ZN(new_n1325));
  OAI211_X1 g1125(.A(KEYINPUT127), .B(new_n1322), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1328));
  AOI211_X1 g1128(.A(new_n1270), .B(new_n1328), .C1(new_n1315), .C2(new_n1273), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1327), .B1(new_n1329), .B2(KEYINPUT63), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1329), .B2(KEYINPUT63), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  OAI211_X1 g1133(.A(KEYINPUT125), .B(new_n1333), .C1(new_n1283), .C2(new_n1328), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1318), .A2(new_n1330), .A3(new_n1332), .A4(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1282), .A2(new_n1337), .A3(new_n1269), .A4(new_n1302), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1338), .B(new_n1325), .C1(new_n1316), .C2(new_n1307), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1329), .A2(new_n1337), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1336), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1335), .A2(new_n1341), .ZN(G405));
  AOI21_X1  g1142(.A(G378), .B1(new_n1206), .B2(new_n1238), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1273), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1305), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1302), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1346), .A2(new_n1336), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1336), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(G402));
endmodule


