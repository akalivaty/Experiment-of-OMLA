//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G43gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(KEYINPUT33), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G113gat), .B2(G120gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G127gat), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n209), .B(new_n217), .C1(new_n212), .C2(new_n214), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G134gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(G134gat), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G169gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G169gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n225), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(KEYINPUT69), .A2(G169gat), .A3(G176gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n224), .B(KEYINPUT68), .C1(G169gat), .C2(G176gat), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT24), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(G183gat), .A3(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  OR3_X1    g050(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n245), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT70), .B1(new_n254), .B2(new_n255), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT71), .B(G183gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT72), .B(G190gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n250), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n238), .A2(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n244), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n225), .A2(new_n226), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT25), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n262), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n256), .A2(new_n257), .A3(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT26), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n240), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n246), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n258), .B2(KEYINPUT27), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(new_n259), .ZN(new_n276));
  INV_X1    g075(.A(new_n259), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT27), .B(G183gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT28), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n272), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n223), .B1(new_n268), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT64), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n244), .A3(new_n263), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT67), .B1(new_n233), .B2(new_n225), .ZN(new_n285));
  AND4_X1   g084(.A1(KEYINPUT67), .A2(new_n225), .A3(new_n227), .A4(new_n229), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n255), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n255), .ZN(new_n291));
  INV_X1    g090(.A(new_n267), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n223), .ZN(new_n294));
  INV_X1    g093(.A(new_n280), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n281), .A2(new_n283), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n283), .A4(new_n296), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n208), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n202), .A2(KEYINPUT33), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n267), .B1(new_n288), .B2(new_n289), .ZN(new_n303));
  AOI211_X1 g102(.A(new_n223), .B(new_n280), .C1(new_n303), .C2(new_n291), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n294), .B1(new_n293), .B2(new_n295), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT74), .B1(new_n306), .B2(new_n283), .ZN(new_n307));
  INV_X1    g106(.A(new_n300), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n301), .B1(new_n309), .B2(new_n206), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n281), .A2(new_n296), .B1(G227gat), .B2(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT34), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n283), .A2(KEYINPUT34), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n311), .A2(new_n312), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n300), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n207), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n205), .B1(new_n317), .B2(new_n302), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n310), .A2(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G228gat), .A2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323));
  AND2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(KEYINPUT22), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G211gat), .B(G218gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT77), .B(KEYINPUT2), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n335), .B(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  AOI211_X1 g137(.A(new_n333), .B(new_n332), .C1(KEYINPUT2), .C2(new_n329), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n328), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n322), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n327), .B2(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(new_n340), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n345), .A2(new_n349), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G22gat), .ZN(new_n353));
  INV_X1    g152(.A(G22gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT83), .A4(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n362), .A2(new_n358), .B1(new_n353), .B2(new_n355), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n321), .A2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT0), .ZN(new_n367));
  XNOR2_X1  g166(.A(G57gat), .B(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n335), .B(KEYINPUT78), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(new_n339), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n223), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n374), .A3(new_n223), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n223), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n341), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT5), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT81), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n376), .A2(new_n384), .A3(new_n378), .A4(new_n381), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n373), .A2(new_n387), .A3(new_n375), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n375), .A2(new_n387), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n379), .A4(new_n378), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n294), .A2(new_n347), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(new_n372), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT80), .B(KEYINPUT5), .C1(new_n392), .C2(new_n379), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n379), .B1(new_n391), .B2(new_n372), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n369), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT6), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n386), .A2(new_n369), .A3(new_n398), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT6), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n400), .B1(new_n403), .B2(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n293), .A2(new_n295), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(new_n342), .B1(G226gat), .B2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(G226gat), .A3(G233gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n328), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n327), .B1(new_n410), .B2(new_n406), .ZN(new_n411));
  XNOR2_X1  g210(.A(G8gat), .B(G36gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413));
  XOR2_X1   g212(.A(new_n412), .B(new_n413), .Z(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(new_n414), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT30), .A4(new_n414), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n417), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n365), .A2(new_n404), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT76), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n426), .B1(new_n310), .B2(new_n316), .ZN(new_n427));
  OAI211_X1 g226(.A(KEYINPUT76), .B(new_n315), .C1(new_n320), .C2(new_n301), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n319), .A2(new_n429), .A3(new_n320), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n309), .A2(new_n206), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n301), .A2(new_n315), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT75), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n427), .B(new_n428), .C1(new_n430), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT86), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n319), .B2(new_n320), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT75), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n427), .A4(new_n428), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n383), .A2(new_n385), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT6), .B1(new_n443), .B2(new_n369), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n369), .B(KEYINPUT84), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n441), .B2(new_n442), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n444), .A2(new_n446), .B1(KEYINPUT6), .B2(new_n399), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT35), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n360), .B2(new_n363), .ZN(new_n449));
  NOR3_X1   g248(.A1(new_n447), .A2(new_n449), .A3(new_n422), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n440), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n438), .A2(new_n452), .A3(new_n427), .A4(new_n428), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n362), .A2(new_n358), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n353), .A2(new_n355), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n359), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n404), .B2(new_n423), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT37), .B1(new_n418), .B2(KEYINPUT85), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT37), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n409), .A2(new_n411), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(new_n419), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT38), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n461), .A2(new_n467), .A3(new_n419), .A4(new_n464), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n447), .A2(new_n466), .A3(new_n415), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n446), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n376), .A2(new_n378), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n380), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT39), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n473), .B1(new_n392), .B2(new_n379), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n445), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n473), .A3(new_n380), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n475), .A2(KEYINPUT40), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT40), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n364), .B1(new_n479), .B2(new_n422), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n460), .B1(new_n469), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n425), .A2(new_n451), .B1(new_n455), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  INV_X1    g282(.A(G1gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT16), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(G1gat), .B2(new_n483), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(G8gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT15), .ZN(new_n491));
  INV_X1    g290(.A(G29gat), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT14), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G29gat), .A2(G36gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n491), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n490), .B2(KEYINPUT15), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n490), .A2(new_n500), .A3(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n494), .A2(new_n496), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n505), .A2(new_n506), .B1(G29gat), .B2(G36gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n497), .A2(KEYINPUT87), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n491), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR3_X1   g308(.A1(new_n504), .A2(KEYINPUT17), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  INV_X1    g311(.A(new_n491), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n490), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  XOR2_X1   g314(.A(G43gat), .B(G50gat), .Z(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT88), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n497), .B(new_n515), .C1(new_n518), .C2(new_n502), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n511), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n489), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n488), .B1(new_n509), .B2(new_n504), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT89), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(KEYINPUT18), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n504), .A2(new_n509), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n489), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n522), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n524), .B(KEYINPUT13), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT18), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n522), .A4(new_n525), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539));
  INV_X1    g338(.A(G197gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT11), .B(G169gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n543), .B(KEYINPUT12), .Z(new_n544));
  INV_X1    g343(.A(KEYINPUT91), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n544), .B1(new_n533), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n538), .A2(new_n546), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550));
  INV_X1    g349(.A(G85gat), .ZN(new_n551));
  INV_X1    g350(.A(G92gat), .ZN(new_n552));
  OAI211_X1 g351(.A(KEYINPUT98), .B(KEYINPUT7), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(KEYINPUT98), .A2(KEYINPUT7), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(G85gat), .A3(G92gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(KEYINPUT8), .A2(new_n559), .B1(new_n551), .B2(new_n552), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n559), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(KEYINPUT99), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(KEYINPUT99), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n556), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT17), .B1(new_n504), .B2(new_n509), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n514), .A2(new_n511), .A3(new_n519), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n568), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT41), .ZN(new_n573));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT97), .Z(new_n575));
  OAI22_X1  g374(.A1(new_n527), .A2(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n550), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n578), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n571), .A2(new_n576), .A3(new_n550), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n575), .A2(new_n573), .ZN(new_n582));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n577), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n584), .ZN(new_n589));
  AOI211_X1 g388(.A(KEYINPUT100), .B(new_n585), .C1(new_n581), .C2(new_n577), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G64gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G57gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n593), .A2(G57gat), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT9), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT92), .B(G57gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n595), .B1(new_n604), .B2(G64gat), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(KEYINPUT9), .B2(new_n601), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT21), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n489), .B1(new_n615), .B2(new_n607), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT94), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n618), .A2(new_n623), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n614), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n613), .A3(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G230gat), .ZN(new_n631));
  INV_X1    g430(.A(G233gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n604), .A2(G64gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(new_n594), .ZN(new_n635));
  INV_X1    g434(.A(new_n606), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n635), .A2(new_n636), .B1(new_n597), .B2(new_n602), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n566), .B1(new_n565), .B2(new_n556), .ZN(new_n638));
  AND4_X1   g437(.A1(new_n566), .A2(new_n556), .A3(new_n560), .A4(new_n561), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n607), .A2(new_n564), .A3(new_n567), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n568), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n633), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n633), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(G176gat), .B(G204gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n648), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n592), .A2(new_n630), .A3(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n482), .A2(new_n549), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n404), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n484), .ZN(G1324gat));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n423), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT16), .B(G8gat), .Z(new_n663));
  AND2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(KEYINPUT42), .ZN(new_n666));
  INV_X1    g465(.A(G8gat), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n665), .B(new_n666), .C1(new_n667), .C2(new_n662), .ZN(G1325gat));
  XNOR2_X1  g467(.A(new_n455), .B(KEYINPUT102), .ZN(new_n669));
  OAI21_X1  g468(.A(G15gat), .B1(new_n659), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n435), .A2(new_n440), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n671), .A2(G15gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n659), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n659), .A2(new_n459), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  NAND2_X1  g475(.A1(new_n451), .A2(new_n425), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n469), .A2(new_n480), .ZN(new_n678));
  INV_X1    g477(.A(new_n460), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n678), .A2(new_n454), .A3(new_n453), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n591), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n549), .A2(new_n630), .A3(new_n656), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n404), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n492), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT45), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT44), .B1(new_n482), .B2(new_n592), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n690));
  NAND3_X1  g489(.A1(new_n681), .A2(new_n591), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n684), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n692), .A2(new_n686), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n492), .B2(new_n693), .ZN(G1328gat));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n422), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n493), .B1(new_n695), .B2(KEYINPUT104), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(KEYINPUT104), .B2(new_n695), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n685), .A2(new_n493), .A3(new_n422), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(G1329gat));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n455), .B(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n692), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n592), .B1(new_n677), .B2(new_n680), .ZN(new_n707));
  INV_X1    g506(.A(new_n671), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n707), .A2(new_n702), .A3(new_n708), .A4(new_n683), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n705), .B2(KEYINPUT105), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n701), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n455), .B(new_n684), .C1(new_n689), .C2(new_n691), .ZN(new_n713));
  OAI211_X1 g512(.A(KEYINPUT47), .B(new_n709), .C1(new_n713), .C2(new_n702), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(G1330gat));
  INV_X1    g514(.A(G50gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n692), .B2(new_n364), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n459), .A2(G50gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT107), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n685), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n717), .A2(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1331gat));
  NAND4_X1  g524(.A1(new_n592), .A2(new_n549), .A3(new_n630), .A4(new_n656), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n482), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n686), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(new_n604), .Z(G1332gat));
  NOR3_X1   g528(.A1(new_n482), .A2(new_n423), .A3(new_n726), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  NAND3_X1  g533(.A1(new_n727), .A2(G71gat), .A3(new_n704), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n482), .A2(new_n671), .A3(new_n726), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n598), .B1(new_n736), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n735), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n364), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  INV_X1    g542(.A(new_n549), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n630), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n657), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n681), .B2(new_n591), .ZN(new_n749));
  INV_X1    g548(.A(new_n690), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n592), .B(new_n750), .C1(new_n677), .C2(new_n680), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT110), .B(new_n747), .C1(new_n749), .C2(new_n751), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n755), .A2(new_n757), .A3(new_n404), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n745), .B1(new_n707), .B2(KEYINPUT111), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n482), .A2(new_n761), .A3(new_n592), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n482), .B2(new_n592), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n707), .A2(KEYINPUT111), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n764), .A2(new_n765), .A3(KEYINPUT51), .A4(new_n745), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n686), .A2(new_n551), .A3(new_n656), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n758), .A2(new_n551), .B1(new_n768), .B2(new_n769), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n422), .A3(new_n756), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n657), .A2(G92gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n422), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n763), .B2(new_n766), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n771), .A2(G92gat), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(KEYINPUT52), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n752), .A2(new_n423), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(G92gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n776), .A2(new_n777), .B1(new_n774), .B2(new_n781), .ZN(G1337gat));
  INV_X1    g581(.A(G99gat), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n783), .A3(new_n708), .A4(new_n656), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n755), .A2(new_n757), .A3(new_n669), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n783), .ZN(G1338gat));
  OAI211_X1 g585(.A(new_n364), .B(new_n747), .C1(new_n749), .C2(new_n751), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n459), .A2(G106gat), .A3(new_n657), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n792), .B1(new_n763), .B2(new_n766), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n790), .A2(new_n793), .A3(KEYINPUT113), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n746), .B1(new_n682), .B2(new_n761), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT51), .B1(new_n796), .B2(new_n765), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n760), .A2(new_n762), .A3(new_n759), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n787), .B2(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n795), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n754), .A2(new_n364), .A3(new_n756), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n793), .B1(new_n802), .B2(G106gat), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n794), .A2(new_n801), .B1(new_n803), .B2(new_n789), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  INV_X1    g604(.A(new_n630), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n643), .A2(new_n644), .A3(new_n633), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n646), .A2(KEYINPUT54), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n652), .B1(new_n645), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n808), .A2(KEYINPUT55), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT55), .B1(new_n808), .B2(new_n810), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n649), .A2(new_n653), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n815), .B(new_n818), .C1(new_n547), .C2(new_n548), .ZN(new_n819));
  INV_X1    g618(.A(new_n544), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n529), .A2(new_n531), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n525), .B1(new_n521), .B2(new_n522), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n538), .A2(new_n820), .B1(new_n543), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n656), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n591), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  AND4_X1   g625(.A1(new_n591), .A2(new_n824), .A3(new_n815), .A4(new_n818), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n806), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n658), .A2(new_n744), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(KEYINPUT115), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT115), .B1(new_n828), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n805), .B1(new_n832), .B2(new_n364), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT116), .B(new_n459), .C1(new_n830), .C2(new_n831), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n671), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n404), .A2(new_n422), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n549), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n832), .A2(new_n404), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n423), .A3(new_n365), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n744), .A2(new_n210), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT117), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n840), .B2(new_n842), .ZN(G1340gat));
  OAI21_X1  g642(.A(new_n211), .B1(new_n840), .B2(new_n657), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n657), .A2(new_n211), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  XOR2_X1   g646(.A(new_n847), .B(KEYINPUT118), .Z(G1341gat));
  NAND4_X1  g647(.A1(new_n835), .A2(G127gat), .A3(new_n630), .A4(new_n836), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n217), .B1(new_n840), .B2(new_n806), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n850), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1342gat));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n365), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n423), .A2(new_n591), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(G134gat), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT56), .ZN(new_n858));
  OAI21_X1  g657(.A(G134gat), .B1(new_n837), .B2(new_n592), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1343gat));
  AND2_X1   g659(.A1(new_n455), .A2(new_n836), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n832), .A2(new_n459), .ZN(new_n862));
  XNOR2_X1  g661(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n459), .B1(new_n828), .B2(new_n829), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n861), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(new_n549), .ZN(new_n869));
  NAND2_X1  g668(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n704), .A2(new_n459), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n549), .A2(G141gat), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n871), .A2(new_n423), .A3(new_n839), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n874), .B(new_n876), .ZN(G1344gat));
  NAND2_X1  g676(.A1(new_n828), .A2(new_n829), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n828), .A2(KEYINPUT115), .A3(new_n829), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n364), .A3(new_n863), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(KEYINPUT57), .B2(new_n865), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n656), .A3(new_n861), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(G148gat), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(KEYINPUT59), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n887), .B1(new_n886), .B2(KEYINPUT59), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n656), .B(new_n861), .C1(new_n864), .C2(new_n867), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n891), .A2(new_n890), .A3(new_n893), .ZN(new_n895));
  OAI22_X1  g694(.A1(new_n888), .A2(new_n889), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n871), .A2(new_n839), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n422), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n892), .A3(new_n656), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(G1345gat));
  INV_X1    g699(.A(G155gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n901), .A3(new_n630), .ZN(new_n902));
  OAI21_X1  g701(.A(G155gat), .B1(new_n868), .B2(new_n806), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n868), .B2(new_n592), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n856), .A2(G162gat), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n905), .B1(new_n897), .B2(new_n906), .ZN(G1347gat));
  NOR2_X1   g706(.A1(new_n686), .A2(new_n423), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n908), .A2(new_n365), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n882), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n233), .A3(new_n744), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT116), .B1(new_n882), .B2(new_n459), .ZN(new_n912));
  INV_X1    g711(.A(new_n834), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n708), .B(new_n908), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT124), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n833), .A2(new_n834), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n916), .A2(new_n917), .A3(new_n708), .A4(new_n908), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n915), .A2(new_n744), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n911), .B1(new_n919), .B2(new_n226), .ZN(G1348gat));
  INV_X1    g719(.A(G176gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n910), .A2(new_n921), .A3(new_n656), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n915), .A2(new_n656), .A3(new_n918), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n921), .ZN(G1349gat));
  NAND3_X1  g723(.A1(new_n915), .A2(new_n630), .A3(new_n918), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n258), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n910), .A2(new_n278), .A3(new_n630), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT125), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1350gat));
  NAND3_X1  g732(.A1(new_n910), .A2(new_n277), .A3(new_n591), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n915), .A2(new_n591), .A3(new_n918), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  AND4_X1   g735(.A1(KEYINPUT126), .A2(new_n935), .A3(new_n936), .A4(G190gat), .ZN(new_n937));
  INV_X1    g736(.A(G190gat), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(KEYINPUT61), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n935), .A2(new_n940), .B1(KEYINPUT126), .B2(new_n936), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n934), .B1(new_n937), .B2(new_n941), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n669), .A2(new_n908), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n884), .A3(new_n744), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n540), .B1(new_n944), .B2(KEYINPUT127), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(KEYINPUT127), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n862), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n744), .A2(new_n540), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n947), .A2(G204gat), .A3(new_n657), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n943), .A2(new_n884), .A3(new_n656), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1353gat));
  OR3_X1    g753(.A1(new_n947), .A2(G211gat), .A3(new_n806), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n943), .A2(new_n884), .A3(new_n630), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n956), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT63), .B1(new_n956), .B2(G211gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(G1354gat));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n884), .A3(new_n591), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(G218gat), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n592), .A2(G218gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n947), .B2(new_n962), .ZN(G1355gat));
endmodule


