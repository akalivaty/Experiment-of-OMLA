//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n464), .B1(G2104), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR3_X1   g042(.A1(new_n467), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n462), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n459), .A2(new_n460), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n474), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n471), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n481), .A2(G124), .B1(G136), .B2(new_n461), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n482), .A2(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n471), .A2(G126), .A3(G2105), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n461), .A2(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n461), .A2(new_n494), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI211_X1 g073(.A(KEYINPUT69), .B(new_n497), .C1(new_n498), .C2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT5), .B1(new_n498), .B2(KEYINPUT69), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(G543), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n507), .A2(new_n516), .ZN(G166));
  NOR2_X1   g092(.A1(new_n508), .A2(new_n509), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n497), .B1(new_n500), .B2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT69), .B1(new_n498), .B2(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n521), .B2(new_n499), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n510), .A2(KEYINPUT71), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n529), .B(G543), .C1(new_n508), .C2(new_n509), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n527), .A2(new_n533), .ZN(G168));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  AOI22_X1  g110(.A1(G52), .A2(new_n531), .B1(new_n522), .B2(G90), .ZN(new_n536));
  AND2_X1   g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n504), .B2(G64), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  OAI21_X1  g114(.A(G651), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n521), .B2(new_n499), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n542), .A2(KEYINPUT72), .A3(new_n537), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n535), .B(new_n536), .C1(new_n540), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT72), .B1(new_n542), .B2(new_n537), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n504), .A2(G64), .ZN(new_n547));
  INV_X1    g122(.A(new_n537), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(new_n539), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(G651), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n535), .B1(new_n550), .B2(new_n536), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n545), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AND2_X1   g128(.A1(new_n504), .A2(G56), .ZN(new_n554));
  AND2_X1   g129(.A1(G68), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n531), .A2(G43), .ZN(new_n557));
  XOR2_X1   g132(.A(KEYINPUT74), .B(G81), .Z(new_n558));
  NAND2_X1  g133(.A1(new_n522), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  AOI22_X1  g141(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n567), .A2(new_n506), .B1(new_n568), .B2(new_n514), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n513), .A2(KEYINPUT75), .A3(G53), .A4(G543), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(G53), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n510), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n573), .A3(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n571), .B(new_n575), .C1(new_n510), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n569), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(KEYINPUT76), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n579), .B1(new_n527), .B2(new_n533), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n526), .A2(new_n525), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n581), .A2(KEYINPUT76), .A3(new_n532), .A4(new_n523), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G286));
  INV_X1    g159(.A(G166), .ZN(G303));
  AOI22_X1  g160(.A1(new_n522), .A2(G87), .B1(G49), .B2(new_n511), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n504), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n506), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n522), .A2(G86), .B1(G48), .B2(new_n511), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n531), .A2(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n514), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n506), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(new_n522), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n504), .A2(G66), .ZN(new_n603));
  INV_X1    g178(.A(G79), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n498), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n531), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g184(.A(new_n608), .B1(G171), .B2(G868), .ZN(G321));
  NOR2_X1   g185(.A1(G299), .A2(G868), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n583), .ZN(G297));
  AOI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n583), .ZN(G280));
  INV_X1    g188(.A(new_n607), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n469), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n471), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT78), .Z(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n481), .A2(G123), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT80), .Z(new_n635));
  AOI211_X1 g210(.A(new_n633), .B(new_n635), .C1(G135), .C2(new_n461), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n642), .A2(KEYINPUT81), .A3(KEYINPUT14), .ZN(new_n643));
  AOI21_X1  g218(.A(KEYINPUT81), .B1(new_n642), .B2(KEYINPUT14), .ZN(new_n644));
  OAI22_X1  g219(.A1(new_n643), .A2(new_n644), .B1(new_n640), .B2(new_n641), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n649), .A2(new_n651), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n628), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2096), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  MUX2_X1   g254(.A(new_n679), .B(new_n678), .S(new_n671), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT82), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n686), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  NOR2_X1   g269(.A1(G16), .A2(G22), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G166), .B2(G16), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT87), .B(G1971), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT88), .Z(new_n699));
  OR2_X1    g274(.A1(G6), .A2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(G305), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT32), .ZN(new_n703));
  INV_X1    g278(.A(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G23), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT85), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G288), .B2(new_n701), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT33), .B(G1976), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT86), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n699), .A2(new_n705), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n461), .A2(G131), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n465), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  INV_X1    g293(.A(G119), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n716), .B1(new_n717), .B2(new_n718), .C1(new_n719), .C2(new_n480), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G29), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT83), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT35), .B(G1991), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n701), .A2(G24), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT84), .Z(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G290), .B2(G16), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1986), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n714), .A2(new_n715), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT36), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n561), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G19), .ZN(new_n735));
  INV_X1    g310(.A(G1341), .ZN(new_n736));
  NAND2_X1  g311(.A1(G160), .A2(G29), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT24), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n722), .B1(new_n738), .B2(G34), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n738), .A2(G34), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2084), .ZN(new_n745));
  OAI22_X1  g320(.A1(new_n735), .A2(new_n736), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT30), .B(G28), .Z(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n636), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G35), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n751), .A2(KEYINPUT100), .A3(G29), .ZN(new_n752));
  OAI21_X1  g327(.A(KEYINPUT100), .B1(new_n751), .B2(G29), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(G162), .C2(new_n722), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT29), .B(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n750), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G1966), .ZN(new_n759));
  NOR2_X1   g334(.A1(G168), .A2(new_n701), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n701), .B2(G21), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n746), .B(new_n758), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n722), .A2(G33), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT25), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n461), .A2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n471), .A2(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n465), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n765), .B(new_n766), .C1(new_n769), .C2(KEYINPUT93), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n763), .B1(new_n772), .B2(new_n722), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G2072), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n761), .A2(new_n759), .B1(new_n773), .B2(G2072), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n774), .B(new_n775), .C1(new_n736), .C2(new_n735), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n701), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n614), .B2(new_n701), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n701), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT23), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n569), .A2(new_n577), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n701), .ZN(new_n784));
  INV_X1    g359(.A(G1956), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n762), .A2(new_n776), .A3(new_n780), .A4(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n722), .A2(G26), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G128), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT89), .Z(new_n793));
  NOR2_X1   g368(.A1(G104), .A2(G2105), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT90), .ZN(new_n795));
  INV_X1    g370(.A(G116), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n467), .B1(new_n796), .B2(G2105), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n795), .A2(new_n797), .B1(G140), .B2(new_n461), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n791), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT92), .B(G2067), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n722), .A2(G27), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT99), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n493), .A2(new_n495), .ZN(new_n805));
  INV_X1    g380(.A(new_n491), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(new_n807), .B2(G29), .ZN(new_n808));
  INV_X1    g383(.A(G2078), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n800), .A2(new_n801), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n802), .A2(new_n810), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n744), .A2(new_n745), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n722), .A2(G32), .ZN(new_n817));
  NAND3_X1  g392(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT26), .Z(new_n819));
  INV_X1    g394(.A(G129), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n480), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G105), .B2(new_n621), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n461), .A2(G141), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT95), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT96), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(KEYINPUT96), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n817), .B1(new_n828), .B2(new_n722), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT27), .B(G1996), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n816), .B1(new_n814), .B2(new_n815), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT97), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n701), .A2(G5), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G171), .B2(new_n701), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1961), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n787), .A2(new_n832), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n733), .A2(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  AND2_X1   g415(.A1(G80), .A2(G543), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n504), .B2(G67), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT101), .B1(new_n842), .B2(new_n506), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n521), .B2(new_n499), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n844), .B(G651), .C1(new_n846), .C2(new_n841), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(G55), .A2(new_n531), .B1(new_n522), .B2(G93), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n850), .A2(KEYINPUT102), .A3(new_n560), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n557), .A2(new_n559), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n555), .B1(new_n504), .B2(G56), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n853), .A2(new_n506), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT102), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n556), .A2(new_n856), .A3(new_n557), .A4(new_n559), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n855), .A2(new_n857), .A3(new_n848), .A4(new_n849), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT38), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n614), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n864));
  NOR3_X1   g439(.A1(new_n863), .A2(new_n864), .A3(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n850), .A2(G860), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT103), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  OR2_X1    g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  NAND2_X1  g444(.A1(new_n828), .A2(G164), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n826), .A2(new_n827), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n807), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n870), .A2(new_n799), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n799), .B1(new_n870), .B2(new_n872), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n873), .A2(new_n874), .B1(new_n771), .B2(new_n770), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n870), .A2(new_n872), .ZN(new_n876));
  INV_X1    g451(.A(new_n799), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n799), .A3(new_n872), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n772), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n625), .B(new_n720), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n461), .A2(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n465), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  INV_X1    g460(.A(G130), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n883), .B1(new_n884), .B2(new_n885), .C1(new_n886), .C2(new_n480), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n882), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT104), .B1(new_n881), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n875), .A3(new_n880), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n636), .B(G160), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(G162), .Z(new_n894));
  NAND4_X1  g469(.A1(new_n888), .A2(new_n875), .A3(new_n880), .A4(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n894), .B1(new_n881), .B2(new_n889), .ZN(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n897), .B2(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g475(.A(new_n617), .B(KEYINPUT105), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n859), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n614), .A2(G299), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n607), .A2(new_n783), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT106), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n607), .A2(KEYINPUT107), .A3(new_n783), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n903), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n614), .B2(G299), .ZN(new_n913));
  AOI22_X1  g488(.A1(new_n911), .A2(new_n912), .B1(new_n904), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n906), .B(KEYINPUT106), .C1(new_n902), .C2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n598), .A2(G305), .ZN(new_n916));
  NAND2_X1  g491(.A1(G166), .A2(G288), .ZN(new_n917));
  OR2_X1    g492(.A1(G166), .A2(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n598), .A2(G305), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(new_n917), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n916), .A2(new_n919), .B1(new_n918), .B2(new_n917), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n921), .A2(KEYINPUT42), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n916), .A2(new_n919), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n917), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n907), .A2(new_n915), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n907), .B2(new_n915), .ZN(new_n933));
  OAI21_X1  g508(.A(G868), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n850), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(G868), .B2(new_n935), .ZN(G295));
  OAI21_X1  g511(.A(new_n934), .B1(G868), .B2(new_n935), .ZN(G331));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n545), .A2(new_n551), .A3(G168), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n536), .B1(new_n540), .B2(new_n543), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT73), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n941), .A2(new_n544), .B1(new_n580), .B2(new_n582), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n859), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n583), .B1(new_n545), .B2(new_n551), .ZN(new_n944));
  INV_X1    g519(.A(G168), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n941), .A2(new_n945), .A3(new_n544), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n944), .A2(new_n946), .A3(new_n851), .A4(new_n858), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n905), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n946), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT109), .A3(new_n859), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(new_n930), .B(new_n948), .C1(new_n954), .C2(new_n914), .ZN(new_n955));
  INV_X1    g530(.A(G37), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n928), .A2(KEYINPUT108), .A3(new_n920), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n928), .B2(new_n920), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n947), .A2(new_n905), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n951), .B2(new_n953), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n905), .A2(new_n912), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n913), .A2(new_n909), .A3(new_n910), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n962), .A2(new_n963), .B1(new_n943), .B2(new_n947), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n959), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n955), .A2(new_n956), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n938), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n955), .A2(new_n956), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n952), .A2(KEYINPUT109), .A3(new_n859), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT109), .B1(new_n952), .B2(new_n859), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n947), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n914), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n930), .B1(new_n973), .B2(new_n948), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(new_n975), .B2(KEYINPUT43), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n968), .B2(new_n974), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n955), .A2(new_n965), .A3(new_n979), .A4(new_n956), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT110), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n968), .C2(new_n974), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n977), .B1(new_n984), .B2(new_n938), .ZN(new_n985));
  AOI211_X1 g560(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n982), .C2(new_n983), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n976), .B1(new_n985), .B2(new_n986), .ZN(G397));
  INV_X1    g562(.A(KEYINPUT126), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(G164), .B2(G1384), .ZN(new_n990));
  INV_X1    g565(.A(new_n470), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT66), .B1(new_n474), .B2(G2105), .ZN(new_n992));
  AOI211_X1 g567(.A(new_n476), .B(new_n465), .C1(new_n472), .C2(new_n473), .ZN(new_n993));
  OAI211_X1 g568(.A(G40), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1996), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n828), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n799), .B(G2067), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n871), .A2(G1996), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n726), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n720), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n720), .A2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n598), .B(G1986), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n995), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n783), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n807), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n994), .ZN(new_n1018));
  NOR2_X1   g593(.A1(G164), .A2(G1384), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n785), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n807), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT56), .B(G2072), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1018), .A2(new_n990), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1012), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT61), .B1(new_n1027), .B2(KEYINPUT122), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n783), .B(new_n1010), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n994), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1956), .B1(new_n1030), .B2(new_n1021), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1026), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1023), .A2(new_n1026), .A3(new_n1012), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1028), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(G160), .A2(G40), .A3(new_n1019), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT58), .B(G1341), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1018), .A2(new_n996), .A3(new_n990), .A4(new_n1024), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n560), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT59), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1044), .B(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1040), .A2(G2067), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1019), .A2(new_n1015), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1018), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1048), .B1(new_n779), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT60), .A3(new_n607), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1034), .A2(KEYINPUT61), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1029), .A2(KEYINPUT119), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1029), .A2(KEYINPUT119), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1056), .A2(new_n1057), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n607), .B1(new_n1052), .B2(KEYINPUT60), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1020), .B1(new_n807), .B2(new_n1013), .ZN(new_n1060));
  NOR3_X1   g635(.A1(G164), .A2(G1384), .A3(new_n1016), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n994), .ZN(new_n1062));
  OAI22_X1  g637(.A1(new_n1062), .A2(G1348), .B1(G2067), .B2(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n1055), .A2(new_n1058), .B1(new_n1059), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1028), .A2(KEYINPUT123), .A3(new_n1036), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1039), .A2(new_n1054), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1034), .A2(new_n614), .A3(new_n1063), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT120), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1024), .A2(new_n990), .A3(G160), .A4(G40), .ZN(new_n1073));
  INV_X1    g648(.A(G1971), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(KEYINPUT112), .A3(new_n1074), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(new_n1078), .C1(G2090), .C2(new_n1051), .ZN(new_n1079));
  NAND3_X1  g654(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(KEYINPUT114), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(KEYINPUT114), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(G166), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1079), .A2(G8), .A3(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT115), .B(G8), .Z(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n586), .A2(G1976), .A3(new_n587), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1089), .B(new_n1090), .C1(new_n1014), .C2(new_n994), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT116), .B(G1976), .Z(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n586), .B2(new_n587), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1040), .A2(new_n1089), .A3(new_n1090), .A4(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1092), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G305), .A2(G1981), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n590), .A2(new_n704), .A3(new_n591), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1098), .A2(KEYINPUT49), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT49), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1040), .A2(new_n1089), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NOR4_X1   g678(.A1(new_n1091), .A2(KEYINPUT117), .A3(KEYINPUT52), .A4(new_n1095), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1097), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1081), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1075), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1022), .A2(G2090), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1089), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  AND3_X1   g685(.A1(new_n1087), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1073), .A2(new_n759), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1049), .A2(new_n1050), .A3(new_n745), .A4(new_n1018), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1084), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G168), .A2(new_n1088), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1088), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT124), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1062), .A2(new_n745), .B1(new_n1073), .B2(new_n759), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1121), .B(new_n1118), .C1(new_n1122), .C2(new_n1088), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1116), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1122), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1115), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1073), .B2(G2078), .ZN(new_n1129));
  INV_X1    g704(.A(G1961), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1051), .A2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  OR3_X1    g707(.A1(new_n1073), .A2(new_n1128), .A3(G2078), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(G301), .A3(new_n1133), .ZN(new_n1134));
  AND4_X1   g709(.A1(KEYINPUT53), .A2(new_n991), .A3(G40), .A4(new_n809), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(new_n1024), .A3(new_n475), .A4(new_n990), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1129), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(new_n1138), .A3(G171), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1137), .B2(G171), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT54), .B(new_n1134), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  AOI21_X1  g717(.A(G301), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1137), .A2(G171), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AND4_X1   g720(.A1(new_n1111), .A2(new_n1127), .A3(new_n1141), .A4(new_n1145), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1127), .A2(KEYINPUT62), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1087), .A2(new_n1105), .A3(new_n1143), .A4(new_n1110), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(KEYINPUT62), .B2(new_n1127), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1072), .A2(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1103), .A2(G1976), .A3(G288), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1099), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1105), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1153), .A2(new_n1102), .B1(new_n1154), .B2(new_n1087), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1087), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1117), .A2(new_n583), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1079), .A2(G8), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1106), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1158), .A2(new_n1156), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1087), .A3(new_n1105), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1155), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1009), .B1(new_n1150), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1005), .A2(new_n995), .ZN(new_n1166));
  NOR4_X1   g741(.A1(G290), .A2(G1986), .A3(new_n990), .A4(new_n994), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  OAI22_X1  g743(.A1(new_n1000), .A2(new_n1004), .B1(G2067), .B2(new_n799), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1166), .A2(new_n1168), .B1(new_n995), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n998), .A2(new_n828), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n995), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n995), .A2(new_n996), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT46), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n988), .B1(new_n1165), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1072), .A2(new_n1146), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1149), .A2(new_n1147), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1164), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1008), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1177), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(KEYINPUT126), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1178), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g760(.A(KEYINPUT127), .ZN(new_n1187));
  NOR2_X1   g761(.A1(G227), .A2(new_n457), .ZN(new_n1188));
  OAI21_X1  g762(.A(new_n1188), .B1(new_n653), .B2(new_n654), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n1187), .B1(G229), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g764(.A(new_n691), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n688), .A2(new_n689), .ZN(new_n1192));
  NOR2_X1   g766(.A1(new_n684), .A2(new_n685), .ZN(new_n1193));
  OAI21_X1  g767(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g768(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g770(.A1(new_n1196), .A2(KEYINPUT127), .A3(new_n655), .A4(new_n1188), .ZN(new_n1197));
  AOI22_X1  g771(.A1(new_n896), .A2(new_n898), .B1(new_n1190), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g772(.A1(new_n1198), .A2(new_n984), .ZN(G225));
  INV_X1    g773(.A(G225), .ZN(G308));
endmodule


