

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  XNOR2_X1 U369 ( .A(n413), .B(n412), .ZN(n521) );
  XNOR2_X1 U370 ( .A(n448), .B(n447), .ZN(n499) );
  NAND2_X1 U371 ( .A1(n662), .A2(n453), .ZN(n659) );
  BUF_X1 U372 ( .A(G146), .Z(n347) );
  INV_X1 U373 ( .A(KEYINPUT64), .ZN(n397) );
  XNOR2_X2 U374 ( .A(n349), .B(n354), .ZN(n653) );
  NAND2_X1 U375 ( .A1(n348), .A2(n583), .ZN(n372) );
  NAND2_X1 U376 ( .A1(n370), .A2(n579), .ZN(n348) );
  XNOR2_X2 U377 ( .A(n368), .B(KEYINPUT32), .ZN(n739) );
  XNOR2_X1 U378 ( .A(n353), .B(G953), .ZN(n500) );
  INV_X1 U379 ( .A(n356), .ZN(n378) );
  NOR2_X1 U380 ( .A1(G237), .A2(G953), .ZN(n433) );
  NAND2_X1 U381 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U382 ( .A(n350), .B(n459), .ZN(n349) );
  XNOR2_X1 U383 ( .A(n351), .B(n635), .ZN(n350) );
  XNOR2_X1 U384 ( .A(n457), .B(G107), .ZN(n351) );
  XNOR2_X1 U385 ( .A(n390), .B(KEYINPUT48), .ZN(n569) );
  NAND2_X1 U386 ( .A1(n379), .A2(n376), .ZN(n587) );
  XNOR2_X1 U387 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U388 ( .A(n465), .B(n725), .ZN(n459) );
  XNOR2_X1 U389 ( .A(n458), .B(KEYINPUT96), .ZN(n635) );
  XNOR2_X1 U390 ( .A(n402), .B(G101), .ZN(n465) );
  XNOR2_X1 U391 ( .A(n455), .B(G137), .ZN(n352) );
  INV_X2 U392 ( .A(KEYINPUT64), .ZN(n353) );
  XNOR2_X2 U393 ( .A(n637), .B(n347), .ZN(n354) );
  XNOR2_X2 U394 ( .A(n456), .B(n352), .ZN(n637) );
  XNOR2_X2 U395 ( .A(n426), .B(n425), .ZN(n456) );
  XNOR2_X1 U396 ( .A(n395), .B(n354), .ZN(n628) );
  NOR2_X2 U397 ( .A1(n574), .A2(n573), .ZN(n368) );
  INV_X1 U398 ( .A(KEYINPUT89), .ZN(n360) );
  OR2_X1 U399 ( .A1(G237), .A2(G902), .ZN(n410) );
  XNOR2_X1 U400 ( .A(KEYINPUT84), .B(KEYINPUT46), .ZN(n392) );
  XNOR2_X1 U401 ( .A(G137), .B(G110), .ZN(n471) );
  XNOR2_X1 U402 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n473) );
  XNOR2_X1 U403 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n402) );
  XNOR2_X1 U404 ( .A(G104), .B(G110), .ZN(n725) );
  XNOR2_X1 U405 ( .A(n406), .B(n423), .ZN(n723) );
  XNOR2_X1 U406 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  XNOR2_X1 U407 ( .A(n387), .B(n386), .ZN(n537) );
  INV_X1 U408 ( .A(KEYINPUT108), .ZN(n386) );
  XNOR2_X1 U409 ( .A(n411), .B(KEYINPUT65), .ZN(n412) );
  NAND2_X1 U410 ( .A1(n512), .A2(n674), .ZN(n413) );
  OR2_X1 U411 ( .A1(n628), .A2(G902), .ZN(n468) );
  XNOR2_X1 U412 ( .A(KEYINPUT22), .B(KEYINPUT76), .ZN(n393) );
  AND2_X1 U413 ( .A1(n549), .A2(n453), .ZN(n454) );
  XNOR2_X1 U414 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U415 ( .A(n479), .B(KEYINPUT25), .ZN(n384) );
  OR2_X2 U416 ( .A1(n560), .A2(n391), .ZN(n390) );
  XNOR2_X1 U417 ( .A(G119), .B(KEYINPUT73), .ZN(n474) );
  INV_X1 U418 ( .A(KEYINPUT70), .ZN(n434) );
  NOR2_X1 U419 ( .A1(n659), .A2(n486), .ZN(n377) );
  NAND2_X1 U420 ( .A1(n659), .A2(n486), .ZN(n380) );
  NAND2_X1 U421 ( .A1(n478), .A2(G217), .ZN(n385) );
  XNOR2_X1 U422 ( .A(G119), .B(G113), .ZN(n405) );
  XNOR2_X1 U423 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U424 ( .A(G131), .B(G116), .ZN(n463) );
  INV_X1 U425 ( .A(G953), .ZN(n729) );
  AND2_X1 U426 ( .A1(n516), .A2(n674), .ZN(n510) );
  NAND2_X1 U427 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U428 ( .A(KEYINPUT0), .ZN(n422) );
  XNOR2_X1 U429 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U430 ( .A(n621), .B(n620), .ZN(n622) );
  XOR2_X1 U431 ( .A(G116), .B(G107), .Z(n355) );
  INV_X1 U432 ( .A(G902), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n559), .B(n392), .ZN(n391) );
  XNOR2_X1 U434 ( .A(n519), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U435 ( .A(n519), .B(KEYINPUT1), .ZN(n485) );
  NOR2_X2 U436 ( .A1(n658), .A2(n603), .ZN(n357) );
  NOR2_X1 U437 ( .A1(n658), .A2(n603), .ZN(n646) );
  XNOR2_X1 U438 ( .A(G128), .B(G140), .ZN(n472) );
  BUF_X1 U439 ( .A(n356), .Z(n660) );
  XNOR2_X2 U440 ( .A(n397), .B(G953), .ZN(n358) );
  NAND2_X1 U441 ( .A1(n683), .A2(n593), .ZN(n493) );
  XNOR2_X1 U442 ( .A(n491), .B(n490), .ZN(n683) );
  NAND2_X1 U443 ( .A1(n379), .A2(n376), .ZN(n359) );
  INV_X1 U444 ( .A(n532), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n382), .B(n600), .ZN(n730) );
  NAND2_X1 U446 ( .A1(n373), .A2(n372), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n374), .B(KEYINPUT87), .ZN(n373) );
  XNOR2_X1 U448 ( .A(n587), .B(n487), .ZN(n489) );
  NAND2_X1 U449 ( .A1(n521), .A2(n421), .ZN(n369) );
  XNOR2_X2 U450 ( .A(n361), .B(n360), .ZN(n580) );
  NOR2_X2 U451 ( .A1(n739), .A2(n575), .ZN(n361) );
  NAND2_X1 U452 ( .A1(n366), .A2(n365), .ZN(n367) );
  XNOR2_X1 U453 ( .A(n363), .B(n364), .ZN(n366) );
  XNOR2_X2 U454 ( .A(n362), .B(G469), .ZN(n519) );
  NOR2_X2 U455 ( .A1(n653), .A2(G902), .ZN(n362) );
  XNOR2_X1 U456 ( .A(n477), .B(n634), .ZN(n363) );
  INV_X1 U457 ( .A(n366), .ZN(n647) );
  NOR2_X1 U458 ( .A1(n470), .A2(n469), .ZN(n364) );
  XNOR2_X2 U459 ( .A(n367), .B(n383), .ZN(n662) );
  NAND2_X1 U460 ( .A1(n593), .A2(n454), .ZN(n394) );
  XNOR2_X2 U461 ( .A(n369), .B(n422), .ZN(n593) );
  XNOR2_X1 U462 ( .A(n578), .B(n577), .ZN(n370) );
  XNOR2_X1 U463 ( .A(n586), .B(KEYINPUT88), .ZN(n375) );
  NAND2_X1 U464 ( .A1(n375), .A2(n599), .ZN(n374) );
  AND2_X2 U465 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U466 ( .A1(n485), .A2(n486), .ZN(n381) );
  NAND2_X1 U467 ( .A1(n730), .A2(n639), .ZN(n602) );
  INV_X1 U468 ( .A(n603), .ZN(n449) );
  NAND2_X1 U469 ( .A1(n603), .A2(G234), .ZN(n450) );
  NOR2_X1 U470 ( .A1(n387), .A2(n591), .ZN(n592) );
  INV_X1 U471 ( .A(n659), .ZN(n388) );
  NAND2_X1 U472 ( .A1(n580), .A2(n576), .ZN(n578) );
  XNOR2_X2 U473 ( .A(n394), .B(n393), .ZN(n574) );
  BUF_X1 U474 ( .A(n646), .Z(n651) );
  BUF_X1 U475 ( .A(n617), .Z(n621) );
  XOR2_X1 U476 ( .A(n467), .B(n466), .Z(n395) );
  INV_X1 U477 ( .A(KEYINPUT104), .ZN(n487) );
  INV_X1 U478 ( .A(KEYINPUT75), .ZN(n577) );
  INV_X1 U479 ( .A(n570), .ZN(n488) );
  INV_X1 U480 ( .A(n506), .ZN(n453) );
  INV_X1 U481 ( .A(KEYINPUT34), .ZN(n492) );
  BUF_X1 U482 ( .A(n519), .Z(n532) );
  NOR2_X1 U483 ( .A1(n555), .A2(n554), .ZN(n556) );
  BUF_X1 U484 ( .A(n584), .Z(n576) );
  XNOR2_X2 U485 ( .A(G125), .B(G146), .ZN(n436) );
  XNOR2_X1 U486 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n436), .B(n396), .ZN(n399) );
  NAND2_X1 U488 ( .A1(n358), .A2(G224), .ZN(n398) );
  XNOR2_X1 U489 ( .A(n399), .B(n398), .ZN(n401) );
  XNOR2_X2 U490 ( .A(KEYINPUT69), .B(KEYINPUT4), .ZN(n455) );
  XNOR2_X2 U491 ( .A(G143), .B(G128), .ZN(n426) );
  XOR2_X1 U492 ( .A(n426), .B(n455), .Z(n400) );
  XNOR2_X1 U493 ( .A(n401), .B(n400), .ZN(n403) );
  XNOR2_X1 U494 ( .A(n403), .B(n459), .ZN(n407) );
  XNOR2_X1 U495 ( .A(n405), .B(n404), .ZN(n461) );
  XNOR2_X1 U496 ( .A(n461), .B(KEYINPUT16), .ZN(n406) );
  XNOR2_X1 U497 ( .A(G122), .B(n355), .ZN(n423) );
  XNOR2_X1 U498 ( .A(n407), .B(n723), .ZN(n617) );
  NOR2_X2 U499 ( .A1(n449), .A2(n617), .ZN(n409) );
  NAND2_X1 U500 ( .A1(G210), .A2(n410), .ZN(n408) );
  XNOR2_X2 U501 ( .A(n409), .B(n408), .ZN(n512) );
  NAND2_X1 U502 ( .A1(G214), .A2(n410), .ZN(n674) );
  INV_X1 U503 ( .A(KEYINPUT19), .ZN(n411) );
  NAND2_X1 U504 ( .A1(G234), .A2(G237), .ZN(n414) );
  XNOR2_X1 U505 ( .A(n414), .B(KEYINPUT92), .ZN(n415) );
  XNOR2_X1 U506 ( .A(KEYINPUT14), .B(n415), .ZN(n416) );
  NAND2_X1 U507 ( .A1(n416), .A2(G952), .ZN(n690) );
  NOR2_X1 U508 ( .A1(G953), .A2(n690), .ZN(n504) );
  NAND2_X1 U509 ( .A1(n416), .A2(G902), .ZN(n417) );
  XNOR2_X1 U510 ( .A(n417), .B(KEYINPUT94), .ZN(n501) );
  NOR2_X1 U511 ( .A1(n729), .A2(G898), .ZN(n418) );
  XNOR2_X1 U512 ( .A(n418), .B(KEYINPUT93), .ZN(n727) );
  NOR2_X1 U513 ( .A1(n501), .A2(n727), .ZN(n419) );
  NOR2_X1 U514 ( .A1(n504), .A2(n419), .ZN(n420) );
  XNOR2_X1 U515 ( .A(KEYINPUT95), .B(n420), .ZN(n421) );
  XOR2_X1 U516 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n424) );
  XNOR2_X1 U517 ( .A(n424), .B(n423), .ZN(n427) );
  INV_X1 U518 ( .A(G134), .ZN(n425) );
  XNOR2_X1 U519 ( .A(n456), .B(n427), .ZN(n431) );
  NAND2_X1 U520 ( .A1(n358), .A2(G234), .ZN(n428) );
  XNOR2_X1 U521 ( .A(n428), .B(KEYINPUT8), .ZN(n470) );
  INV_X1 U522 ( .A(G217), .ZN(n429) );
  OR2_X1 U523 ( .A1(n470), .A2(n429), .ZN(n430) );
  XNOR2_X1 U524 ( .A(n431), .B(n430), .ZN(n605) );
  NAND2_X1 U525 ( .A1(n605), .A2(n365), .ZN(n432) );
  XNOR2_X1 U526 ( .A(n432), .B(G478), .ZN(n498) );
  XNOR2_X1 U527 ( .A(n433), .B(KEYINPUT78), .ZN(n460) );
  NAND2_X1 U528 ( .A1(n460), .A2(G214), .ZN(n437) );
  XNOR2_X1 U529 ( .A(n434), .B(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U530 ( .A(n436), .B(n435), .ZN(n634) );
  XNOR2_X1 U531 ( .A(n437), .B(n634), .ZN(n446) );
  XOR2_X1 U532 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n439) );
  XNOR2_X1 U533 ( .A(KEYINPUT101), .B(KEYINPUT11), .ZN(n438) );
  XNOR2_X1 U534 ( .A(n439), .B(n438), .ZN(n444) );
  XNOR2_X2 U535 ( .A(G140), .B(G131), .ZN(n458) );
  XNOR2_X1 U536 ( .A(G113), .B(G104), .ZN(n441) );
  XNOR2_X1 U537 ( .A(G143), .B(G122), .ZN(n440) );
  XNOR2_X1 U538 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U539 ( .A(n458), .B(n442), .ZN(n443) );
  XNOR2_X1 U540 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U541 ( .A(n446), .B(n445), .ZN(n610) );
  OR2_X1 U542 ( .A1(n610), .A2(G902), .ZN(n448) );
  XOR2_X1 U543 ( .A(KEYINPUT13), .B(G475), .Z(n447) );
  NOR2_X1 U544 ( .A1(n498), .A2(n499), .ZN(n549) );
  XNOR2_X1 U545 ( .A(KEYINPUT20), .B(n450), .ZN(n478) );
  AND2_X1 U546 ( .A1(n478), .A2(G221), .ZN(n452) );
  INV_X1 U547 ( .A(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U548 ( .A(n452), .B(n451), .ZN(n506) );
  NAND2_X1 U549 ( .A1(n500), .A2(G227), .ZN(n457) );
  NAND2_X1 U550 ( .A1(n460), .A2(G210), .ZN(n462) );
  XNOR2_X1 U551 ( .A(n462), .B(n461), .ZN(n467) );
  XNOR2_X1 U552 ( .A(n463), .B(KEYINPUT5), .ZN(n464) );
  XNOR2_X1 U553 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X2 U554 ( .A(n468), .B(G472), .ZN(n591) );
  INV_X1 U555 ( .A(G221), .ZN(n469) );
  XNOR2_X1 U556 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U557 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U558 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT79), .Z(n479) );
  OR2_X1 U560 ( .A1(n591), .A2(n662), .ZN(n480) );
  OR2_X1 U561 ( .A1(n378), .A2(n480), .ZN(n481) );
  NOR2_X1 U562 ( .A1(n574), .A2(n481), .ZN(n575) );
  XOR2_X1 U563 ( .A(G110), .B(n575), .Z(G12) );
  XNOR2_X1 U564 ( .A(n591), .B(KEYINPUT6), .ZN(n570) );
  NOR2_X1 U565 ( .A1(n574), .A2(n488), .ZN(n482) );
  XOR2_X1 U566 ( .A(KEYINPUT86), .B(n482), .Z(n484) );
  NAND2_X1 U567 ( .A1(n660), .A2(n662), .ZN(n483) );
  NOR2_X1 U568 ( .A1(n484), .A2(n483), .ZN(n598) );
  XOR2_X1 U569 ( .A(G101), .B(n598), .Z(G3) );
  INV_X1 U570 ( .A(KEYINPUT77), .ZN(n486) );
  NAND2_X1 U571 ( .A1(n489), .A2(n488), .ZN(n491) );
  XNOR2_X1 U572 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n490) );
  XNOR2_X1 U573 ( .A(n493), .B(n492), .ZN(n495) );
  NAND2_X1 U574 ( .A1(n499), .A2(n498), .ZN(n538) );
  INV_X1 U575 ( .A(n538), .ZN(n494) );
  NAND2_X1 U576 ( .A1(n495), .A2(n494), .ZN(n497) );
  XNOR2_X1 U577 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U578 ( .A(n497), .B(n496), .ZN(n584) );
  XNOR2_X1 U579 ( .A(n576), .B(G122), .ZN(G24) );
  XOR2_X1 U580 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n514) );
  INV_X1 U581 ( .A(n498), .ZN(n524) );
  XNOR2_X1 U582 ( .A(KEYINPUT102), .B(n499), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n524), .A2(n525), .ZN(n557) );
  XNOR2_X1 U584 ( .A(KEYINPUT105), .B(n557), .ZN(n714) );
  NOR2_X1 U585 ( .A1(n501), .A2(n358), .ZN(n502) );
  XOR2_X1 U586 ( .A(KEYINPUT106), .B(n502), .Z(n503) );
  NOR2_X1 U587 ( .A1(G900), .A2(n503), .ZN(n505) );
  NOR2_X1 U588 ( .A1(n505), .A2(n504), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n535), .A2(n506), .ZN(n508) );
  INV_X1 U590 ( .A(n662), .ZN(n507) );
  NAND2_X1 U591 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U592 ( .A(n509), .B(KEYINPUT71), .ZN(n516) );
  NAND2_X1 U593 ( .A1(n714), .A2(n510), .ZN(n511) );
  NOR2_X1 U594 ( .A1(n511), .A2(n570), .ZN(n562) );
  BUF_X2 U595 ( .A(n512), .Z(n565) );
  NAND2_X1 U596 ( .A1(n562), .A2(n565), .ZN(n513) );
  XOR2_X1 U597 ( .A(n514), .B(n513), .Z(n515) );
  NOR2_X2 U598 ( .A1(n515), .A2(n660), .ZN(n719) );
  XNOR2_X1 U599 ( .A(n719), .B(KEYINPUT85), .ZN(n547) );
  INV_X1 U600 ( .A(KEYINPUT47), .ZN(n529) );
  XOR2_X1 U601 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n518) );
  NAND2_X1 U602 ( .A1(n516), .A2(n591), .ZN(n517) );
  XOR2_X1 U603 ( .A(n518), .B(n517), .Z(n520) );
  NOR2_X1 U604 ( .A1(n520), .A2(n532), .ZN(n551) );
  INV_X1 U605 ( .A(n551), .ZN(n523) );
  INV_X1 U606 ( .A(n521), .ZN(n522) );
  NOR2_X1 U607 ( .A1(n523), .A2(n522), .ZN(n712) );
  NOR2_X1 U608 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U609 ( .A(n526), .B(KEYINPUT103), .ZN(n704) );
  NAND2_X1 U610 ( .A1(n557), .A2(n704), .ZN(n594) );
  INV_X1 U611 ( .A(n594), .ZN(n680) );
  NOR2_X1 U612 ( .A1(n680), .A2(KEYINPUT81), .ZN(n527) );
  NAND2_X1 U613 ( .A1(n712), .A2(n527), .ZN(n528) );
  NAND2_X1 U614 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U615 ( .A1(n712), .A2(KEYINPUT47), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n531), .A2(n530), .ZN(n541) );
  NAND2_X1 U617 ( .A1(n591), .A2(n674), .ZN(n533) );
  XNOR2_X1 U618 ( .A(n533), .B(KEYINPUT30), .ZN(n534) );
  NOR2_X1 U619 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U620 ( .A1(n537), .A2(n536), .ZN(n555) );
  INV_X1 U621 ( .A(n565), .ZN(n548) );
  OR2_X1 U622 ( .A1(n548), .A2(n538), .ZN(n539) );
  NOR2_X1 U623 ( .A1(n555), .A2(n539), .ZN(n540) );
  XNOR2_X1 U624 ( .A(KEYINPUT109), .B(n540), .ZN(n738) );
  NAND2_X1 U625 ( .A1(n541), .A2(n738), .ZN(n545) );
  AND2_X1 U626 ( .A1(n712), .A2(KEYINPUT81), .ZN(n542) );
  NOR2_X1 U627 ( .A1(n542), .A2(KEYINPUT47), .ZN(n543) );
  NOR2_X1 U628 ( .A1(n594), .A2(n543), .ZN(n544) );
  NOR2_X1 U629 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n560) );
  XOR2_X1 U631 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n553) );
  XOR2_X1 U632 ( .A(KEYINPUT38), .B(n548), .Z(n554) );
  INV_X1 U633 ( .A(n554), .ZN(n675) );
  NAND2_X1 U634 ( .A1(n675), .A2(n674), .ZN(n679) );
  INV_X1 U635 ( .A(n549), .ZN(n678) );
  NOR2_X1 U636 ( .A1(n679), .A2(n678), .ZN(n550) );
  XNOR2_X1 U637 ( .A(KEYINPUT41), .B(n550), .ZN(n673) );
  INV_X1 U638 ( .A(n673), .ZN(n692) );
  NAND2_X1 U639 ( .A1(n692), .A2(n551), .ZN(n552) );
  XNOR2_X1 U640 ( .A(n553), .B(n552), .ZN(n741) );
  XNOR2_X1 U641 ( .A(n556), .B(KEYINPUT39), .ZN(n561) );
  OR2_X1 U642 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U643 ( .A(n558), .B(KEYINPUT40), .ZN(n742) );
  NAND2_X1 U644 ( .A1(n741), .A2(n742), .ZN(n559) );
  NOR2_X1 U645 ( .A1(n561), .A2(n704), .ZN(n721) );
  INV_X1 U646 ( .A(n721), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n562), .A2(n660), .ZN(n564) );
  XNOR2_X1 U648 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n563) );
  XNOR2_X1 U649 ( .A(n564), .B(n563), .ZN(n566) );
  OR2_X1 U650 ( .A1(n566), .A2(n565), .ZN(n722) );
  NAND2_X1 U651 ( .A1(n567), .A2(n722), .ZN(n568) );
  NOR2_X2 U652 ( .A1(n569), .A2(n568), .ZN(n639) );
  NOR2_X1 U653 ( .A1(n660), .A2(n662), .ZN(n571) );
  NAND2_X1 U654 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U655 ( .A(n572), .B(KEYINPUT80), .ZN(n573) );
  INV_X1 U656 ( .A(KEYINPUT44), .ZN(n579) );
  INV_X1 U657 ( .A(n580), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n577), .A2(KEYINPUT44), .ZN(n581) );
  OR2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n583) );
  INV_X1 U660 ( .A(n584), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n585), .A2(KEYINPUT44), .ZN(n586) );
  XOR2_X1 U662 ( .A(KEYINPUT31), .B(KEYINPUT99), .Z(n590) );
  INV_X1 U663 ( .A(n591), .ZN(n665) );
  NOR2_X1 U664 ( .A1(n359), .A2(n665), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n588), .B(KEYINPUT98), .ZN(n670) );
  NAND2_X1 U666 ( .A1(n670), .A2(n593), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n590), .B(n589), .ZN(n717) );
  AND2_X1 U668 ( .A1(n593), .A2(n592), .ZN(n705) );
  NOR2_X1 U669 ( .A1(n717), .A2(n705), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n594), .B(KEYINPUT81), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U673 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n600) );
  INV_X1 U674 ( .A(KEYINPUT2), .ZN(n601) );
  XNOR2_X2 U675 ( .A(n602), .B(n601), .ZN(n658) );
  NAND2_X1 U676 ( .A1(n357), .A2(G478), .ZN(n604) );
  XOR2_X1 U677 ( .A(n605), .B(n604), .Z(n608) );
  INV_X1 U678 ( .A(n358), .ZN(n607) );
  INV_X1 U679 ( .A(G952), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n631) );
  INV_X1 U681 ( .A(n631), .ZN(n656) );
  NOR2_X1 U682 ( .A1(n608), .A2(n656), .ZN(G63) );
  NAND2_X1 U683 ( .A1(n357), .A2(G475), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n609) );
  XNOR2_X1 U685 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n613), .A2(n631), .ZN(n616) );
  XOR2_X1 U687 ( .A(KEYINPUT122), .B(KEYINPUT60), .Z(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT66), .ZN(n615) );
  XNOR2_X1 U689 ( .A(n616), .B(n615), .ZN(G60) );
  NAND2_X1 U690 ( .A1(n357), .A2(G210), .ZN(n623) );
  XNOR2_X1 U691 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n619) );
  XNOR2_X1 U692 ( .A(KEYINPUT55), .B(KEYINPUT90), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n624), .A2(n631), .ZN(n626) );
  INV_X1 U696 ( .A(KEYINPUT56), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(G51) );
  NAND2_X1 U698 ( .A1(n646), .A2(G472), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT91), .B(KEYINPUT62), .ZN(n627) );
  XNOR2_X1 U700 ( .A(n630), .B(n629), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U702 ( .A(n633), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U703 ( .A(n635), .B(n634), .Z(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(n641) );
  XNOR2_X1 U705 ( .A(n641), .B(KEYINPUT126), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U707 ( .A1(n640), .A2(n500), .ZN(n645) );
  XOR2_X1 U708 ( .A(G227), .B(n641), .Z(n642) );
  NAND2_X1 U709 ( .A1(n642), .A2(G900), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n643), .A2(G953), .ZN(n644) );
  NAND2_X1 U711 ( .A1(n645), .A2(n644), .ZN(G72) );
  NAND2_X1 U712 ( .A1(n651), .A2(G217), .ZN(n649) );
  XOR2_X1 U713 ( .A(KEYINPUT123), .B(n647), .Z(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n650) );
  NOR2_X1 U715 ( .A1(n650), .A2(n656), .ZN(G66) );
  NAND2_X1 U716 ( .A1(n651), .A2(G469), .ZN(n655) );
  XOR2_X1 U717 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n652) );
  XNOR2_X1 U718 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U719 ( .A(n655), .B(n654), .ZN(n657) );
  NOR2_X1 U720 ( .A1(n657), .A2(n656), .ZN(G54) );
  BUF_X1 U721 ( .A(n658), .Z(n698) );
  NAND2_X1 U722 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U723 ( .A(KEYINPUT50), .B(n661), .Z(n668) );
  OR2_X1 U724 ( .A1(n662), .A2(n453), .ZN(n664) );
  XOR2_X1 U725 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n663) );
  XNOR2_X1 U726 ( .A(n664), .B(n663), .ZN(n666) );
  NAND2_X1 U727 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U728 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U729 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U730 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  NOR2_X1 U731 ( .A1(n673), .A2(n672), .ZN(n688) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U733 ( .A(KEYINPUT117), .B(n676), .Z(n677) );
  NOR2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U735 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U736 ( .A1(n682), .A2(n681), .ZN(n686) );
  BUF_X1 U737 ( .A(n683), .Z(n684) );
  INV_X1 U738 ( .A(n684), .ZN(n685) );
  NOR2_X1 U739 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U741 ( .A(n689), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U742 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U743 ( .A1(n692), .A2(n684), .ZN(n693) );
  XNOR2_X1 U744 ( .A(n693), .B(KEYINPUT118), .ZN(n694) );
  NAND2_X1 U745 ( .A1(n694), .A2(n729), .ZN(n695) );
  NOR2_X1 U746 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U747 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U748 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n699) );
  XNOR2_X1 U749 ( .A(n700), .B(n699), .ZN(G75) );
  XOR2_X1 U750 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n702) );
  NAND2_X1 U751 ( .A1(n705), .A2(n714), .ZN(n701) );
  XNOR2_X1 U752 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U753 ( .A(G104), .B(n703), .ZN(G6) );
  XOR2_X1 U754 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n707) );
  INV_X1 U755 ( .A(n704), .ZN(n716) );
  NAND2_X1 U756 ( .A1(n705), .A2(n716), .ZN(n706) );
  XNOR2_X1 U757 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U758 ( .A(G107), .B(n708), .ZN(G9) );
  XOR2_X1 U759 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n710) );
  NAND2_X1 U760 ( .A1(n712), .A2(n716), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n710), .B(n709), .ZN(n711) );
  XOR2_X1 U762 ( .A(G128), .B(n711), .Z(G30) );
  NAND2_X1 U763 ( .A1(n712), .A2(n714), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n713), .B(n347), .ZN(G48) );
  NAND2_X1 U765 ( .A1(n717), .A2(n714), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n715), .B(G113), .ZN(G15) );
  NAND2_X1 U767 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(G116), .ZN(G18) );
  XNOR2_X1 U769 ( .A(n719), .B(G125), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U771 ( .A(G134), .B(n721), .Z(G36) );
  XNOR2_X1 U772 ( .A(G140), .B(n722), .ZN(G42) );
  XOR2_X1 U773 ( .A(n723), .B(KEYINPUT125), .Z(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U775 ( .A(G101), .B(n726), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n737) );
  AND2_X1 U777 ( .A1(n730), .A2(n729), .ZN(n735) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n731) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n731), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G898), .ZN(n733) );
  XOR2_X1 U781 ( .A(KEYINPUT124), .B(n733), .Z(n734) );
  NOR2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U783 ( .A(n737), .B(n736), .ZN(G69) );
  XNOR2_X1 U784 ( .A(G143), .B(n738), .ZN(G45) );
  XNOR2_X1 U785 ( .A(G119), .B(KEYINPUT127), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(G21) );
  XNOR2_X1 U787 ( .A(G137), .B(n741), .ZN(G39) );
  XNOR2_X1 U788 ( .A(G131), .B(n742), .ZN(G33) );
endmodule

