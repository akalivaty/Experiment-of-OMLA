

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774;

  NAND2_X1 U385 ( .A1(n377), .A2(n376), .ZN(n665) );
  AND2_X1 U386 ( .A1(n365), .A2(n678), .ZN(n375) );
  AND2_X1 U387 ( .A1(n369), .A2(n378), .ZN(n365) );
  XNOR2_X1 U388 ( .A(n364), .B(n463), .ZN(n564) );
  NAND2_X1 U389 ( .A1(n460), .A2(n627), .ZN(n364) );
  NAND2_X2 U390 ( .A1(n363), .A2(n380), .ZN(n379) );
  NAND2_X1 U391 ( .A1(n384), .A2(n372), .ZN(n363) );
  XNOR2_X2 U392 ( .A(KEYINPUT93), .B(G110), .ZN(n406) );
  OR2_X1 U393 ( .A1(n637), .A2(G902), .ZN(n421) );
  XNOR2_X1 U394 ( .A(n449), .B(n448), .ZN(n758) );
  NOR2_X1 U395 ( .A1(n596), .A2(n695), .ZN(n576) );
  XNOR2_X2 U396 ( .A(n527), .B(n526), .ZN(n649) );
  NAND2_X2 U397 ( .A1(n401), .A2(n398), .ZN(n648) );
  AND2_X2 U398 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X2 U399 ( .A(G116), .B(G113), .ZN(n409) );
  XNOR2_X2 U400 ( .A(n412), .B(n411), .ZN(n479) );
  XNOR2_X2 U401 ( .A(G128), .B(KEYINPUT65), .ZN(n412) );
  INV_X2 U402 ( .A(G953), .ZN(n767) );
  XNOR2_X1 U403 ( .A(n386), .B(n541), .ZN(n740) );
  XNOR2_X1 U404 ( .A(n385), .B(KEYINPUT100), .ZN(n729) );
  NOR2_X1 U405 ( .A1(n705), .A2(n571), .ZN(n508) );
  XNOR2_X1 U406 ( .A(n518), .B(n517), .ZN(n553) );
  XNOR2_X1 U407 ( .A(n433), .B(n432), .ZN(n516) );
  XNOR2_X1 U408 ( .A(n421), .B(n420), .ZN(n538) );
  XNOR2_X1 U409 ( .A(n479), .B(n413), .ZN(n457) );
  XNOR2_X1 U410 ( .A(n407), .B(n406), .ZN(n756) );
  XNOR2_X1 U411 ( .A(G146), .B(G125), .ZN(n452) );
  XNOR2_X1 U412 ( .A(KEYINPUT69), .B(G101), .ZN(n441) );
  XNOR2_X1 U413 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n451) );
  XNOR2_X1 U414 ( .A(G107), .B(G104), .ZN(n407) );
  BUF_X1 U415 ( .A(n665), .Z(n366) );
  BUF_X1 U416 ( .A(n450), .Z(n367) );
  XNOR2_X1 U417 ( .A(n756), .B(n441), .ZN(n450) );
  XNOR2_X2 U418 ( .A(n393), .B(n520), .ZN(n719) );
  OR2_X2 U419 ( .A1(n564), .A2(n466), .ZN(n595) );
  XNOR2_X1 U420 ( .A(n457), .B(n414), .ZN(n436) );
  NAND2_X1 U421 ( .A1(n648), .A2(n644), .ZN(n515) );
  XNOR2_X1 U422 ( .A(n436), .B(KEYINPUT96), .ZN(n766) );
  XNOR2_X1 U423 ( .A(KEYINPUT15), .B(G902), .ZN(n627) );
  XNOR2_X1 U424 ( .A(n538), .B(KEYINPUT1), .ZN(n512) );
  INV_X1 U425 ( .A(G143), .ZN(n411) );
  INV_X1 U426 ( .A(n627), .ZN(n378) );
  XNOR2_X1 U427 ( .A(KEYINPUT72), .B(G131), .ZN(n495) );
  INV_X1 U428 ( .A(G902), .ZN(n484) );
  XNOR2_X1 U429 ( .A(G146), .B(G137), .ZN(n438) );
  XNOR2_X1 U430 ( .A(G140), .B(G137), .ZN(n423) );
  NAND2_X1 U431 ( .A1(n530), .A2(KEYINPUT44), .ZN(n382) );
  NAND2_X1 U432 ( .A1(n516), .A2(n688), .ZN(n518) );
  NOR2_X1 U433 ( .A1(n584), .A2(n472), .ZN(n473) );
  INV_X1 U434 ( .A(KEYINPUT4), .ZN(n413) );
  XNOR2_X1 U435 ( .A(KEYINPUT16), .B(G122), .ZN(n448) );
  XNOR2_X1 U436 ( .A(n447), .B(KEYINPUT83), .ZN(n404) );
  AND2_X1 U437 ( .A1(n446), .A2(n445), .ZN(n447) );
  NOR2_X1 U438 ( .A1(n534), .A2(KEYINPUT32), .ZN(n399) );
  INV_X1 U439 ( .A(G472), .ZN(n389) );
  NOR2_X1 U440 ( .A1(n629), .A2(G902), .ZN(n388) );
  AND2_X1 U441 ( .A1(n521), .A2(n553), .ZN(n387) );
  NOR2_X1 U442 ( .A1(n735), .A2(n707), .ZN(n589) );
  NOR2_X1 U443 ( .A1(G953), .A2(G237), .ZN(n487) );
  XOR2_X1 U444 ( .A(G140), .B(KEYINPUT12), .Z(n489) );
  XNOR2_X1 U445 ( .A(n452), .B(KEYINPUT10), .ZN(n497) );
  XNOR2_X1 U446 ( .A(G143), .B(G104), .ZN(n494) );
  XNOR2_X1 U447 ( .A(G113), .B(G122), .ZN(n490) );
  XOR2_X1 U448 ( .A(KEYINPUT101), .B(KEYINPUT11), .Z(n491) );
  AND2_X1 U449 ( .A1(n623), .A2(KEYINPUT2), .ZN(n397) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n468) );
  INV_X1 U451 ( .A(G237), .ZN(n461) );
  XNOR2_X1 U452 ( .A(n390), .B(n444), .ZN(n629) );
  INV_X1 U453 ( .A(n436), .ZN(n390) );
  XNOR2_X1 U454 ( .A(G119), .B(G128), .ZN(n425) );
  XNOR2_X1 U455 ( .A(n497), .B(n423), .ZN(n765) );
  XNOR2_X1 U456 ( .A(G116), .B(G134), .ZN(n474) );
  XNOR2_X1 U457 ( .A(G122), .B(KEYINPUT103), .ZN(n475) );
  XOR2_X1 U458 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n476) );
  XNOR2_X1 U459 ( .A(n766), .B(n419), .ZN(n637) );
  BUF_X1 U460 ( .A(n516), .Z(n689) );
  BUF_X2 U461 ( .A(n512), .Z(n696) );
  NAND2_X1 U462 ( .A1(n392), .A2(n368), .ZN(n376) );
  NAND2_X1 U463 ( .A1(n665), .A2(G475), .ZN(n661) );
  XNOR2_X1 U464 ( .A(n758), .B(n450), .ZN(n459) );
  NOR2_X1 U465 ( .A1(n767), .A2(G952), .ZN(n671) );
  XNOR2_X1 U466 ( .A(n395), .B(KEYINPUT40), .ZN(n581) );
  NAND2_X1 U467 ( .A1(n396), .A2(n569), .ZN(n395) );
  NAND2_X1 U468 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U469 ( .A1(n387), .A2(n539), .ZN(n385) );
  AND2_X1 U470 ( .A1(n378), .A2(KEYINPUT2), .ZN(n368) );
  AND2_X1 U471 ( .A1(n624), .A2(n623), .ZN(n369) );
  XOR2_X1 U472 ( .A(n426), .B(KEYINPUT23), .Z(n370) );
  AND2_X1 U473 ( .A1(n550), .A2(n528), .ZN(n372) );
  XNOR2_X1 U474 ( .A(n551), .B(KEYINPUT45), .ZN(n373) );
  OR2_X1 U475 ( .A1(n626), .A2(KEYINPUT78), .ZN(n374) );
  NAND2_X1 U476 ( .A1(n391), .A2(n375), .ZN(n377) );
  NOR2_X1 U477 ( .A1(n662), .A2(n671), .ZN(n664) );
  NOR2_X1 U478 ( .A1(n632), .A2(n671), .ZN(n634) );
  NOR2_X1 U479 ( .A1(n640), .A2(n671), .ZN(n642) );
  NOR2_X1 U480 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X2 U481 ( .A(n379), .B(n373), .ZN(n678) );
  NAND2_X1 U482 ( .A1(n382), .A2(n381), .ZN(n380) );
  AND2_X1 U483 ( .A1(n550), .A2(n531), .ZN(n381) );
  XNOR2_X1 U484 ( .A(n529), .B(KEYINPUT44), .ZN(n384) );
  NAND2_X1 U485 ( .A1(n740), .A2(n729), .ZN(n547) );
  NAND2_X1 U486 ( .A1(n387), .A2(n540), .ZN(n386) );
  XNOR2_X2 U487 ( .A(n388), .B(n389), .ZN(n691) );
  NAND2_X1 U488 ( .A1(n675), .A2(n374), .ZN(n391) );
  INV_X1 U489 ( .A(n675), .ZN(n392) );
  NAND2_X1 U490 ( .A1(n625), .A2(KEYINPUT78), .ZN(n675) );
  INV_X1 U491 ( .A(n696), .ZN(n686) );
  NAND2_X1 U492 ( .A1(n719), .A2(n521), .ZN(n523) );
  NAND2_X1 U493 ( .A1(n696), .A2(n394), .ZN(n393) );
  NOR2_X1 U494 ( .A1(n597), .A2(n685), .ZN(n394) );
  INV_X1 U495 ( .A(n581), .ZN(n647) );
  INV_X1 U496 ( .A(n618), .ZN(n396) );
  NAND2_X1 U497 ( .A1(n624), .A2(n397), .ZN(n676) );
  INV_X1 U498 ( .A(n404), .ZN(n400) );
  NAND2_X1 U499 ( .A1(n534), .A2(KEYINPUT32), .ZN(n402) );
  NAND2_X1 U500 ( .A1(n404), .A2(KEYINPUT32), .ZN(n403) );
  XNOR2_X2 U501 ( .A(n511), .B(n510), .ZN(n534) );
  INV_X1 U502 ( .A(n678), .ZN(n748) );
  NAND2_X1 U503 ( .A1(n678), .A2(n405), .ZN(n625) );
  INV_X1 U504 ( .A(n676), .ZN(n405) );
  XNOR2_X2 U505 ( .A(n409), .B(n408), .ZN(n449) );
  XNOR2_X2 U506 ( .A(KEYINPUT3), .B(G119), .ZN(n408) );
  XOR2_X1 U507 ( .A(KEYINPUT24), .B(G110), .Z(n410) );
  INV_X1 U508 ( .A(KEYINPUT108), .ZN(n598) );
  XNOR2_X1 U509 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U510 ( .A(n503), .B(n502), .ZN(n545) );
  INV_X1 U511 ( .A(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U512 ( .A(n495), .B(G134), .ZN(n414) );
  XNOR2_X1 U513 ( .A(G146), .B(KEYINPUT80), .ZN(n416) );
  NAND2_X1 U514 ( .A1(n767), .A2(G227), .ZN(n415) );
  XNOR2_X1 U515 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U516 ( .A(n417), .B(n423), .ZN(n418) );
  XNOR2_X1 U517 ( .A(n367), .B(n418), .ZN(n419) );
  XNOR2_X1 U518 ( .A(KEYINPUT74), .B(G469), .ZN(n420) );
  NAND2_X1 U519 ( .A1(G234), .A2(n767), .ZN(n422) );
  XOR2_X1 U520 ( .A(KEYINPUT8), .B(n422), .Z(n480) );
  NAND2_X1 U521 ( .A1(n480), .A2(G221), .ZN(n424) );
  XNOR2_X1 U522 ( .A(n424), .B(n765), .ZN(n428) );
  XNOR2_X1 U523 ( .A(n410), .B(n425), .ZN(n426) );
  XNOR2_X1 U524 ( .A(n370), .B(KEYINPUT97), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n428), .B(n427), .ZN(n650) );
  NAND2_X1 U526 ( .A1(n650), .A2(n484), .ZN(n433) );
  NAND2_X1 U527 ( .A1(G234), .A2(n627), .ZN(n429) );
  XNOR2_X1 U528 ( .A(KEYINPUT20), .B(n429), .ZN(n505) );
  NAND2_X1 U529 ( .A1(n505), .A2(G217), .ZN(n431) );
  XNOR2_X1 U530 ( .A(KEYINPUT79), .B(KEYINPUT25), .ZN(n430) );
  XNOR2_X1 U531 ( .A(n431), .B(n430), .ZN(n432) );
  INV_X1 U532 ( .A(n689), .ZN(n434) );
  NAND2_X1 U533 ( .A1(n512), .A2(n434), .ZN(n435) );
  XNOR2_X1 U534 ( .A(n435), .B(KEYINPUT107), .ZN(n446) );
  NAND2_X1 U535 ( .A1(G210), .A2(n487), .ZN(n437) );
  XNOR2_X1 U536 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U537 ( .A(n449), .B(n439), .ZN(n443) );
  XNOR2_X1 U538 ( .A(KEYINPUT99), .B(KEYINPUT5), .ZN(n440) );
  XNOR2_X1 U539 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U540 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U541 ( .A(n691), .B(KEYINPUT6), .ZN(n597) );
  XNOR2_X1 U542 ( .A(n597), .B(KEYINPUT84), .ZN(n445) );
  XNOR2_X1 U543 ( .A(n452), .B(n451), .ZN(n455) );
  NAND2_X1 U544 ( .A1(n767), .A2(G224), .ZN(n453) );
  XNOR2_X1 U545 ( .A(n453), .B(KEYINPUT81), .ZN(n454) );
  XNOR2_X1 U546 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U547 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U548 ( .A(n459), .B(n458), .ZN(n666) );
  INV_X1 U549 ( .A(n666), .ZN(n460) );
  NAND2_X1 U550 ( .A1(n484), .A2(n461), .ZN(n465) );
  NAND2_X1 U551 ( .A1(n465), .A2(G210), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n462), .B(KEYINPUT94), .ZN(n463) );
  NAND2_X1 U553 ( .A1(n465), .A2(G214), .ZN(n703) );
  INV_X1 U554 ( .A(n703), .ZN(n466) );
  XNOR2_X1 U555 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n467) );
  XNOR2_X1 U556 ( .A(n595), .B(n467), .ZN(n584) );
  XNOR2_X1 U557 ( .A(n468), .B(KEYINPUT14), .ZN(n469) );
  NAND2_X1 U558 ( .A1(G952), .A2(n469), .ZN(n716) );
  NOR2_X1 U559 ( .A1(n716), .A2(G953), .ZN(n560) );
  NAND2_X1 U560 ( .A1(G902), .A2(n469), .ZN(n557) );
  INV_X1 U561 ( .A(G898), .ZN(n751) );
  NAND2_X1 U562 ( .A1(G953), .A2(n751), .ZN(n760) );
  NOR2_X1 U563 ( .A1(n557), .A2(n760), .ZN(n470) );
  OR2_X1 U564 ( .A1(n560), .A2(n470), .ZN(n471) );
  XNOR2_X1 U565 ( .A(n471), .B(KEYINPUT95), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n473), .B(KEYINPUT0), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n474), .B(G107), .ZN(n478) );
  XNOR2_X1 U568 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U569 ( .A(n478), .B(n477), .Z(n483) );
  NAND2_X1 U570 ( .A1(G217), .A2(n480), .ZN(n481) );
  XNOR2_X1 U571 ( .A(n479), .B(n481), .ZN(n482) );
  XNOR2_X1 U572 ( .A(n483), .B(n482), .ZN(n655) );
  NAND2_X1 U573 ( .A1(n655), .A2(n484), .ZN(n486) );
  INV_X1 U574 ( .A(G478), .ZN(n485) );
  XNOR2_X1 U575 ( .A(n486), .B(n485), .ZN(n542) );
  NAND2_X1 U576 ( .A1(G214), .A2(n487), .ZN(n488) );
  XNOR2_X1 U577 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U579 ( .A(n493), .B(n492), .ZN(n499) );
  XNOR2_X1 U580 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U581 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U582 ( .A(n499), .B(n498), .ZN(n659) );
  NOR2_X1 U583 ( .A1(G902), .A2(n659), .ZN(n503) );
  XNOR2_X1 U584 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n501) );
  INV_X1 U585 ( .A(G475), .ZN(n500) );
  NAND2_X1 U586 ( .A1(n542), .A2(n545), .ZN(n504) );
  XOR2_X1 U587 ( .A(n504), .B(KEYINPUT105), .Z(n705) );
  XOR2_X1 U588 ( .A(KEYINPUT21), .B(KEYINPUT98), .Z(n507) );
  NAND2_X1 U589 ( .A1(n505), .A2(G221), .ZN(n506) );
  XOR2_X1 U590 ( .A(n507), .B(n506), .Z(n571) );
  XNOR2_X1 U591 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  NAND2_X1 U592 ( .A1(n521), .A2(n509), .ZN(n511) );
  XNOR2_X1 U593 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n510) );
  NOR2_X1 U594 ( .A1(n689), .A2(n691), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n686), .A2(n513), .ZN(n514) );
  OR2_X1 U596 ( .A1(n534), .A2(n514), .ZN(n644) );
  XNOR2_X2 U597 ( .A(n515), .B(KEYINPUT89), .ZN(n529) );
  INV_X1 U598 ( .A(n571), .ZN(n688) );
  INV_X1 U599 ( .A(KEYINPUT70), .ZN(n517) );
  INV_X1 U600 ( .A(n553), .ZN(n685) );
  INV_X1 U601 ( .A(KEYINPUT91), .ZN(n519) );
  XNOR2_X1 U602 ( .A(n519), .B(KEYINPUT33), .ZN(n520) );
  XNOR2_X1 U603 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n522) );
  XNOR2_X1 U604 ( .A(n523), .B(n522), .ZN(n524) );
  NOR2_X1 U605 ( .A1(n545), .A2(n542), .ZN(n607) );
  NAND2_X1 U606 ( .A1(n524), .A2(n607), .ZN(n527) );
  INV_X1 U607 ( .A(KEYINPUT82), .ZN(n525) );
  XNOR2_X1 U608 ( .A(n525), .B(KEYINPUT35), .ZN(n526) );
  AND2_X1 U609 ( .A1(n649), .A2(KEYINPUT88), .ZN(n528) );
  INV_X1 U610 ( .A(KEYINPUT88), .ZN(n535) );
  NAND2_X1 U611 ( .A1(n529), .A2(n535), .ZN(n530) );
  INV_X1 U612 ( .A(n649), .ZN(n531) );
  NAND2_X1 U613 ( .A1(n597), .A2(n689), .ZN(n532) );
  OR2_X1 U614 ( .A1(n696), .A2(n532), .ZN(n533) );
  OR2_X1 U615 ( .A1(n534), .A2(n533), .ZN(n645) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n536) );
  NAND2_X1 U617 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U618 ( .A1(n645), .A2(n537), .ZN(n549) );
  BUF_X1 U619 ( .A(n538), .Z(n552) );
  INV_X1 U620 ( .A(n691), .ZN(n695) );
  AND2_X1 U621 ( .A1(n552), .A2(n695), .ZN(n539) );
  AND2_X1 U622 ( .A1(n696), .A2(n691), .ZN(n540) );
  INV_X1 U623 ( .A(KEYINPUT31), .ZN(n541) );
  INV_X1 U624 ( .A(n542), .ZN(n544) );
  OR2_X1 U625 ( .A1(n545), .A2(n544), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT104), .ZN(n738) );
  NAND2_X1 U627 ( .A1(n545), .A2(n544), .ZN(n741) );
  AND2_X1 U628 ( .A1(n738), .A2(n741), .ZN(n707) );
  INV_X1 U629 ( .A(n707), .ZN(n546) );
  AND2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U631 ( .A1(n549), .A2(n548), .ZN(n550) );
  INV_X1 U632 ( .A(KEYINPUT64), .ZN(n551) );
  NAND2_X1 U633 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U634 ( .A(n554), .B(KEYINPUT109), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n691), .A2(n703), .ZN(n556) );
  XNOR2_X1 U636 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n555) );
  XNOR2_X1 U637 ( .A(n556), .B(n555), .ZN(n561) );
  OR2_X1 U638 ( .A1(n767), .A2(n557), .ZN(n558) );
  NOR2_X1 U639 ( .A1(n558), .A2(G900), .ZN(n559) );
  NOR2_X1 U640 ( .A1(n560), .A2(n559), .ZN(n572) );
  NOR2_X1 U641 ( .A1(n561), .A2(n572), .ZN(n562) );
  AND2_X1 U642 ( .A1(n563), .A2(n562), .ZN(n610) );
  INV_X1 U643 ( .A(KEYINPUT77), .ZN(n565) );
  XNOR2_X1 U644 ( .A(n565), .B(KEYINPUT38), .ZN(n566) );
  XNOR2_X1 U645 ( .A(n564), .B(n566), .ZN(n702) );
  NAND2_X1 U646 ( .A1(n610), .A2(n702), .ZN(n568) );
  INV_X1 U647 ( .A(KEYINPUT39), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n568), .B(n567), .ZN(n618) );
  INV_X1 U649 ( .A(n738), .ZN(n569) );
  NAND2_X1 U650 ( .A1(n703), .A2(n702), .ZN(n706) );
  NOR2_X1 U651 ( .A1(n705), .A2(n706), .ZN(n570) );
  XNOR2_X1 U652 ( .A(KEYINPUT41), .B(n570), .ZN(n718) );
  NOR2_X1 U653 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U654 ( .A(KEYINPUT73), .B(n573), .ZN(n574) );
  OR2_X1 U655 ( .A1(n574), .A2(n516), .ZN(n596) );
  XOR2_X1 U656 ( .A(KEYINPUT111), .B(KEYINPUT28), .Z(n575) );
  XNOR2_X1 U657 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U658 ( .A1(n577), .A2(n552), .ZN(n585) );
  NOR2_X1 U659 ( .A1(n718), .A2(n585), .ZN(n579) );
  XNOR2_X1 U660 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n578) );
  XNOR2_X1 U661 ( .A(n579), .B(n578), .ZN(n774) );
  INV_X1 U662 ( .A(n774), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n583) );
  INV_X1 U664 ( .A(KEYINPUT46), .ZN(n582) );
  XNOR2_X1 U665 ( .A(n583), .B(n582), .ZN(n615) );
  OR2_X1 U666 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U667 ( .A(KEYINPUT85), .ZN(n586) );
  XNOR2_X1 U668 ( .A(n587), .B(n586), .ZN(n735) );
  XNOR2_X1 U669 ( .A(KEYINPUT47), .B(KEYINPUT71), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n605), .A2(KEYINPUT76), .ZN(n588) );
  NAND2_X1 U671 ( .A1(n589), .A2(n588), .ZN(n594) );
  INV_X1 U672 ( .A(n589), .ZN(n592) );
  INV_X1 U673 ( .A(KEYINPUT76), .ZN(n590) );
  NOR2_X1 U674 ( .A1(n590), .A2(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U675 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U676 ( .A1(n594), .A2(n593), .ZN(n613) );
  INV_X1 U677 ( .A(n595), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n599), .B(n598), .ZN(n600) );
  NOR2_X1 U680 ( .A1(n738), .A2(n600), .ZN(n619) );
  NAND2_X1 U681 ( .A1(n601), .A2(n619), .ZN(n603) );
  XNOR2_X1 U682 ( .A(KEYINPUT36), .B(KEYINPUT113), .ZN(n602) );
  XNOR2_X1 U683 ( .A(n603), .B(n602), .ZN(n604) );
  AND2_X1 U684 ( .A1(n696), .A2(n604), .ZN(n744) );
  NOR2_X1 U685 ( .A1(n605), .A2(KEYINPUT76), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n744), .A2(n606), .ZN(n611) );
  INV_X1 U687 ( .A(n607), .ZN(n608) );
  NOR2_X1 U688 ( .A1(n608), .A2(n564), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n643) );
  AND2_X1 U690 ( .A1(n611), .A2(n643), .ZN(n612) );
  AND2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U693 ( .A(KEYINPUT48), .ZN(n616) );
  XNOR2_X1 U694 ( .A(n617), .B(n616), .ZN(n624) );
  OR2_X1 U695 ( .A1(n618), .A2(n741), .ZN(n746) );
  NAND2_X1 U696 ( .A1(n703), .A2(n619), .ZN(n620) );
  OR2_X1 U697 ( .A1(n696), .A2(n620), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT43), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n622), .A2(n564), .ZN(n646) );
  AND2_X1 U700 ( .A1(n746), .A2(n646), .ZN(n623) );
  INV_X1 U701 ( .A(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n665), .A2(G472), .ZN(n631) );
  XNOR2_X1 U703 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(G57) );
  NAND2_X1 U707 ( .A1(n665), .A2(G469), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n635) );
  XNOR2_X1 U709 ( .A(n635), .B(KEYINPUT58), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U711 ( .A(n639), .B(n638), .ZN(n640) );
  INV_X1 U712 ( .A(KEYINPUT121), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(G54) );
  XNOR2_X1 U714 ( .A(n643), .B(G143), .ZN(G45) );
  XNOR2_X1 U715 ( .A(n644), .B(G110), .ZN(G12) );
  XNOR2_X1 U716 ( .A(n645), .B(G101), .ZN(G3) );
  XNOR2_X1 U717 ( .A(n646), .B(G140), .ZN(G42) );
  XOR2_X1 U718 ( .A(G131), .B(n647), .Z(G33) );
  XNOR2_X1 U719 ( .A(n648), .B(G119), .ZN(G21) );
  XNOR2_X1 U720 ( .A(n649), .B(G122), .ZN(G24) );
  NAND2_X1 U721 ( .A1(n366), .A2(G217), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n650), .B(KEYINPUT123), .ZN(n651) );
  XNOR2_X1 U723 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n653), .A2(n671), .ZN(G66) );
  NAND2_X1 U725 ( .A1(n366), .A2(G478), .ZN(n654) );
  XOR2_X1 U726 ( .A(n655), .B(n654), .Z(n656) );
  NOR2_X1 U727 ( .A1(n656), .A2(n671), .ZN(G63) );
  XOR2_X1 U728 ( .A(KEYINPUT92), .B(KEYINPUT122), .Z(n657) );
  XNOR2_X1 U729 ( .A(n657), .B(KEYINPUT59), .ZN(n658) );
  XNOR2_X1 U730 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(G60) );
  NAND2_X1 U734 ( .A1(n665), .A2(G210), .ZN(n670) );
  XOR2_X1 U735 ( .A(KEYINPUT90), .B(KEYINPUT54), .Z(n667) );
  XNOR2_X1 U736 ( .A(n667), .B(KEYINPUT55), .ZN(n668) );
  XNOR2_X1 U737 ( .A(n666), .B(n668), .ZN(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(n669), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X1 U740 ( .A1(n678), .A2(KEYINPUT2), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(KEYINPUT86), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n676), .A2(KEYINPUT78), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n675), .A2(n679), .ZN(n681) );
  OR2_X1 U745 ( .A1(n369), .A2(KEYINPUT2), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT87), .ZN(n725) );
  NAND2_X1 U749 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n687), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U752 ( .A(KEYINPUT49), .B(n690), .Z(n692) );
  NOR2_X1 U753 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U754 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n685), .A2(n695), .ZN(n697) );
  NAND2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U758 ( .A(KEYINPUT51), .B(n700), .ZN(n701) );
  NOR2_X1 U759 ( .A1(n701), .A2(n718), .ZN(n714) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U763 ( .A(KEYINPUT119), .B(n708), .Z(n709) );
  NOR2_X1 U764 ( .A1(n710), .A2(n709), .ZN(n712) );
  INV_X1 U765 ( .A(n719), .ZN(n711) );
  NOR2_X1 U766 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U767 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n715), .B(KEYINPUT52), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n717), .A2(n716), .ZN(n723) );
  INV_X1 U770 ( .A(n718), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n721), .A2(n767), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U775 ( .A(KEYINPUT53), .B(n726), .Z(G75) );
  XNOR2_X1 U776 ( .A(G104), .B(KEYINPUT115), .ZN(n728) );
  NOR2_X1 U777 ( .A1(n738), .A2(n729), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(G6) );
  NOR2_X1 U779 ( .A1(n729), .A2(n741), .ZN(n731) );
  XNOR2_X1 U780 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U782 ( .A(G107), .B(n732), .ZN(G9) );
  NOR2_X1 U783 ( .A1(n741), .A2(n735), .ZN(n734) );
  XNOR2_X1 U784 ( .A(G128), .B(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U785 ( .A(n734), .B(n733), .ZN(G30) );
  NOR2_X1 U786 ( .A1(n738), .A2(n735), .ZN(n736) );
  XOR2_X1 U787 ( .A(KEYINPUT116), .B(n736), .Z(n737) );
  XNOR2_X1 U788 ( .A(G146), .B(n737), .ZN(G48) );
  NOR2_X1 U789 ( .A1(n738), .A2(n740), .ZN(n739) );
  XOR2_X1 U790 ( .A(G113), .B(n739), .Z(G15) );
  NOR2_X1 U791 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U792 ( .A(G116), .B(KEYINPUT117), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G18) );
  XNOR2_X1 U794 ( .A(n744), .B(G125), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n745), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U796 ( .A(n746), .B(G134), .ZN(n747) );
  XNOR2_X1 U797 ( .A(KEYINPUT118), .B(n747), .ZN(G36) );
  NOR2_X1 U798 ( .A1(n748), .A2(G953), .ZN(n754) );
  XOR2_X1 U799 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n750) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n752) );
  NOR2_X1 U802 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U803 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U804 ( .A(n755), .B(KEYINPUT125), .ZN(n764) );
  XNOR2_X1 U805 ( .A(n756), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U806 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U807 ( .A(G101), .B(n759), .ZN(n761) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U809 ( .A(n762), .B(KEYINPUT127), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(G69) );
  XOR2_X1 U811 ( .A(n766), .B(n765), .Z(n769) );
  XNOR2_X1 U812 ( .A(n369), .B(n769), .ZN(n768) );
  NAND2_X1 U813 ( .A1(n768), .A2(n767), .ZN(n773) );
  XOR2_X1 U814 ( .A(G227), .B(n769), .Z(n770) );
  NAND2_X1 U815 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U816 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U817 ( .A1(n773), .A2(n772), .ZN(G72) );
  XOR2_X1 U818 ( .A(G137), .B(n774), .Z(G39) );
endmodule

