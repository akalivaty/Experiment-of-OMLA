//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G119), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n187), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AND3_X1   g008(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n196));
  OAI22_X1  g010(.A1(new_n195), .A2(new_n196), .B1(KEYINPUT2), .B2(G113), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n194), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G143), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(new_n203), .B2(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n204), .A2(new_n207), .B1(new_n210), .B2(new_n205), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  OR2_X1    g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT11), .B1(new_n214), .B2(G134), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(G137), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G137), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT11), .A4(G134), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n213), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n217), .A2(new_n213), .A3(new_n221), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n211), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n210), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT64), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n232), .A3(G143), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n232), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n201), .B1(new_n235), .B2(new_n200), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n203), .B2(G143), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT68), .B(new_n204), .C1(new_n239), .C2(new_n229), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n227), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(G134), .B1(new_n218), .B2(new_n220), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n216), .A2(G137), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n217), .A2(new_n221), .A3(new_n212), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n199), .B(new_n224), .C1(new_n241), .C2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(G237), .A2(G953), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G210), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n249), .B(KEYINPUT27), .Z(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n237), .A2(new_n240), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n210), .A2(new_n226), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n246), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n223), .A2(new_n222), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n204), .A2(new_n207), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n210), .A2(new_n205), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT30), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n224), .C1(new_n241), .C2(new_n246), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT71), .B1(new_n266), .B2(new_n198), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n268));
  AOI211_X1 g082(.A(new_n268), .B(new_n199), .C1(new_n263), .C2(new_n265), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n254), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT31), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n198), .B1(new_n257), .B2(new_n262), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(new_n247), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n247), .A2(new_n272), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n252), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n278), .B(new_n254), .C1(new_n267), .C2(new_n269), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT72), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n280), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n280), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT74), .B1(new_n274), .B2(new_n276), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n276), .A2(KEYINPUT74), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT29), .A4(new_n253), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n283), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n247), .B1(new_n267), .B2(new_n269), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT29), .B1(new_n292), .B2(new_n252), .ZN(new_n293));
  INV_X1    g107(.A(new_n274), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(new_n275), .A3(new_n253), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n294), .A2(new_n297), .A3(new_n275), .A4(new_n253), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n291), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  OAI22_X1  g114(.A1(new_n286), .A2(new_n287), .B1(new_n282), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G104), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(new_n302), .B2(G107), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n304));
  INV_X1    g118(.A(G107), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G104), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(G107), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT78), .A4(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(G101), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n303), .A2(new_n306), .A3(new_n313), .A4(new_n307), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n314), .A2(KEYINPUT4), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n310), .A2(G101), .A3(new_n311), .A4(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n198), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n194), .A2(new_n197), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n191), .A2(KEYINPUT5), .A3(new_n193), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n322), .B(G113), .C1(KEYINPUT5), .C2(new_n193), .ZN(new_n323));
  XNOR2_X1  g137(.A(G104), .B(G107), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT81), .B1(new_n324), .B2(new_n313), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n305), .A2(G104), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n307), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G101), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n321), .A2(new_n323), .A3(new_n314), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G110), .B(G122), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n319), .A2(new_n335), .A3(new_n331), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G224), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(G953), .ZN(new_n341));
  AOI211_X1 g155(.A(G125), .B(new_n227), .C1(new_n237), .C2(new_n240), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n259), .B2(new_n260), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n255), .A2(new_n343), .A3(new_n256), .ZN(new_n346));
  INV_X1    g160(.A(new_n341), .ZN(new_n347));
  INV_X1    g161(.A(new_n344), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n351), .A3(new_n336), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n339), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT86), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n339), .A2(new_n350), .A3(new_n355), .A4(new_n352), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n335), .B(KEYINPUT8), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n358), .A2(new_n322), .A3(G113), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n325), .A2(new_n329), .A3(new_n314), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n359), .A2(new_n360), .A3(new_n320), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n321), .A2(new_n323), .B1(new_n330), .B2(new_n314), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n338), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n341), .A2(KEYINPUT7), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n346), .B2(new_n348), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n341), .B(new_n344), .C1(new_n241), .C2(new_n343), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(new_n356), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(G210), .B1(G237), .B2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT87), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n354), .A2(new_n373), .A3(new_n371), .A4(new_n356), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G214), .B1(G237), .B2(G902), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n372), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT91), .ZN(new_n382));
  NOR2_X1   g196(.A1(G475), .A2(G902), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT19), .ZN(new_n386));
  INV_X1    g200(.A(G140), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G125), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n343), .A2(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(KEYINPUT88), .ZN(new_n391));
  XNOR2_X1  g205(.A(G125), .B(G140), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT19), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n235), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n387), .A3(G125), .ZN(new_n397));
  OAI211_X1 g211(.A(G146), .B(new_n397), .C1(new_n390), .C2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n385), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT19), .B1(new_n392), .B2(new_n393), .ZN(new_n401));
  AND4_X1   g215(.A1(new_n393), .A2(new_n388), .A3(new_n389), .A4(KEYINPUT19), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n203), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT89), .A3(new_n398), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n248), .A2(G143), .A3(G214), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(G143), .B1(new_n248), .B2(G214), .ZN(new_n407));
  OAI21_X1  g221(.A(G131), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n212), .A3(new_n405), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n404), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n392), .A2(new_n203), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n208), .B2(new_n392), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT18), .B(G131), .C1(new_n406), .C2(new_n407), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n409), .A2(new_n405), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n302), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT17), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n410), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT90), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n397), .B1(new_n390), .B2(new_n396), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n208), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n398), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n408), .A2(new_n410), .A3(new_n431), .A4(new_n424), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n408), .A2(new_n424), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n426), .A2(new_n430), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n421), .A3(new_n418), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n384), .B1(new_n423), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n382), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n434), .A2(new_n421), .A3(new_n418), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n421), .B1(new_n412), .B2(new_n418), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n383), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n437), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n421), .B1(new_n434), .B2(new_n418), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n283), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G475), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT92), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(KEYINPUT92), .A3(new_n447), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT70), .B(G116), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT14), .A3(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(G122), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n187), .A2(G122), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(G107), .B(new_n452), .C1(new_n455), .C2(KEYINPUT14), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n229), .A2(G143), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n225), .A2(G143), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n216), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n216), .B1(new_n457), .B2(new_n459), .ZN(new_n462));
  OAI221_X1 g276(.A(new_n456), .B1(G107), .B2(new_n455), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n200), .A2(KEYINPUT13), .A3(G128), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n464), .B(KEYINPUT93), .Z(new_n465));
  OAI21_X1  g279(.A(new_n457), .B1(KEYINPUT13), .B2(new_n458), .ZN(new_n466));
  OAI21_X1  g280(.A(G134), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n305), .B1(new_n453), .B2(new_n454), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n455), .A2(G107), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n467), .B(new_n460), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT9), .B(G234), .ZN(new_n472));
  INV_X1    g286(.A(G217), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n472), .A2(new_n473), .A3(G953), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n470), .A3(new_n474), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n283), .ZN(new_n479));
  INV_X1    g293(.A(G478), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(G902), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  INV_X1    g297(.A(new_n481), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G953), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G952), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n488), .B1(G234), .B2(G237), .ZN(new_n489));
  AOI211_X1 g303(.A(new_n283), .B(new_n487), .C1(G234), .C2(G237), .ZN(new_n490));
  XNOR2_X1  g304(.A(KEYINPUT21), .B(G898), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n486), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n449), .A2(new_n450), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n381), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G221), .ZN(new_n496));
  INV_X1    g310(.A(new_n472), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n283), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT10), .B1(new_n241), .B2(new_n360), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n225), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n210), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n360), .B1(new_n501), .B2(new_n256), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT10), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n316), .A2(new_n211), .A3(new_n318), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n316), .A2(KEYINPUT80), .A3(new_n211), .A4(new_n318), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n505), .A2(new_n510), .A3(new_n258), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT82), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n499), .A2(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n258), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G110), .B(G140), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n487), .A2(G227), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n505), .A2(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(new_n258), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n516), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n255), .A2(new_n256), .A3(new_n360), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT83), .ZN(new_n527));
  INV_X1    g341(.A(new_n502), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT83), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n241), .A2(new_n529), .A3(new_n360), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n531), .A2(new_n532), .A3(new_n522), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n532), .B1(new_n531), .B2(new_n522), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n520), .B1(new_n535), .B2(new_n516), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G469), .B1(new_n537), .B2(G902), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n514), .B1(new_n513), .B2(new_n258), .ZN(new_n539));
  AND4_X1   g353(.A1(new_n514), .A2(new_n505), .A3(new_n510), .A4(new_n258), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n523), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n519), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n516), .A3(new_n520), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(KEYINPUT84), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT84), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n541), .A2(new_n546), .A3(new_n519), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n544), .A2(new_n545), .A3(new_n283), .A4(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n498), .B1(new_n538), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  INV_X1    g366(.A(G119), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(G128), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(G128), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n229), .A2(G119), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n555), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT24), .B(G110), .ZN(new_n561));
  OAI221_X1 g375(.A(new_n429), .B1(new_n557), .B2(new_n558), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n551), .A2(new_n556), .A3(new_n558), .ZN(new_n563));
  INV_X1    g377(.A(new_n561), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n559), .B2(new_n555), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT75), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n560), .A2(new_n561), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n551), .A2(new_n558), .A3(new_n556), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n398), .A2(new_n413), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT76), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT76), .ZN(new_n575));
  AOI211_X1 g389(.A(new_n575), .B(new_n572), .C1(new_n566), .C2(new_n570), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n562), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n487), .A2(G221), .A3(G234), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n578), .B(new_n579), .Z(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n562), .B(new_n580), .C1(new_n574), .C2(new_n576), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n550), .B1(new_n584), .B2(G902), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n582), .A2(KEYINPUT25), .A3(new_n283), .A4(new_n583), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n473), .B1(G234), .B2(new_n283), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n584), .ZN(new_n590));
  INV_X1    g404(.A(new_n588), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n283), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT77), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n301), .A2(new_n495), .A3(new_n549), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n280), .A2(new_n285), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n282), .B1(new_n280), .B2(new_n283), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n600), .A2(new_n601), .A3(new_n595), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n602), .A2(new_n549), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n375), .A2(KEYINPUT94), .A3(new_n377), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n371), .A2(new_n356), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n373), .A4(new_n354), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n379), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(G478), .A2(G902), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n479), .B2(G478), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n478), .B(KEYINPUT33), .Z(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(new_n611), .B2(G478), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n444), .A2(KEYINPUT92), .A3(new_n447), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n448), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n608), .A2(new_n614), .A3(new_n492), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n603), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n379), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n606), .B1(new_n372), .B2(new_n374), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n377), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n438), .A2(new_n442), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n622), .A2(new_n623), .B1(new_n437), .B2(new_n436), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n438), .A2(new_n442), .A3(KEYINPUT95), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n624), .A2(new_n625), .B1(G475), .B2(new_n446), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n621), .A2(new_n626), .A3(new_n486), .A4(new_n607), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n492), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n603), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT35), .B(G107), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  OR2_X1    g445(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n577), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n577), .A2(new_n632), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n633), .A2(new_n593), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT96), .B1(new_n589), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n591), .B1(new_n585), .B2(new_n586), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n639), .A3(new_n635), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n600), .A2(new_n601), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n495), .A2(new_n549), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n622), .A2(new_n623), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n443), .A3(new_n625), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n447), .A3(new_n486), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n608), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n301), .A2(new_n649), .A3(new_n641), .ZN(new_n650));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n490), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n489), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n549), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n225), .ZN(G30));
  XNOR2_X1  g471(.A(new_n654), .B(KEYINPUT39), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n549), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT97), .Z(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(KEYINPUT40), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n378), .A2(new_n380), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT38), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n589), .A2(new_n636), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n619), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n613), .A2(new_n448), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n668), .A3(new_n486), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n599), .A2(KEYINPUT32), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n280), .A2(new_n281), .A3(new_n285), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n292), .A2(new_n253), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n273), .A2(new_n247), .A3(new_n252), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n283), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n664), .B(new_n669), .C1(new_n672), .C2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n661), .A2(new_n662), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  OAI211_X1 g494(.A(new_n612), .B(new_n654), .C1(new_n613), .C2(new_n448), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n608), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n301), .A2(new_n682), .A3(new_n549), .A4(new_n641), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT98), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n589), .A2(KEYINPUT96), .A3(new_n636), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n639), .B1(new_n638), .B2(new_n635), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n293), .A2(new_n299), .ZN(new_n688));
  INV_X1    g502(.A(new_n291), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n282), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n687), .B1(new_n672), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n693), .A3(new_n549), .A4(new_n682), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n684), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT99), .B(G146), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G48));
  NAND2_X1  g511(.A1(new_n301), .A2(new_n596), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n544), .A2(new_n283), .A3(new_n547), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  INV_X1    g514(.A(new_n498), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n548), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n615), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n628), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  INV_X1    g522(.A(new_n608), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n701), .A3(new_n548), .A4(new_n700), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n667), .A3(new_n493), .A4(new_n692), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND4_X1  g527(.A1(new_n668), .A2(new_n486), .A3(new_n607), .A4(new_n621), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n702), .A3(new_n492), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT100), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n288), .A2(new_n716), .A3(new_n289), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n288), .B2(new_n289), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n717), .A2(new_n718), .A3(new_n253), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n271), .A2(new_n279), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n285), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n280), .A2(new_n283), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G472), .ZN(new_n725));
  OAI211_X1 g539(.A(KEYINPUT101), .B(new_n285), .C1(new_n719), .C2(new_n720), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n715), .A2(new_n596), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  AOI21_X1  g543(.A(new_n601), .B1(new_n721), .B2(new_n722), .ZN(new_n730));
  INV_X1    g544(.A(new_n681), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n665), .A3(new_n731), .A4(new_n726), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n710), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n343), .ZN(G27));
  NAND2_X1  g548(.A1(G469), .A2(G902), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n524), .A2(KEYINPUT102), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n535), .A2(new_n516), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n519), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n516), .A2(new_n739), .A3(new_n520), .A4(new_n523), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n738), .A3(G469), .A4(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n548), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n619), .B1(new_n378), .B2(new_n380), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n701), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n690), .B1(new_n670), .B2(new_n671), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(new_n595), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n301), .A2(KEYINPUT103), .A3(new_n596), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(new_n749), .A3(KEYINPUT104), .A4(new_n750), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n698), .A2(new_n744), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n731), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n753), .A2(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n212), .ZN(G33));
  INV_X1    g573(.A(new_n744), .ZN(new_n760));
  INV_X1    g574(.A(new_n654), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n648), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(new_n596), .A3(new_n301), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  AOI21_X1  g578(.A(new_n642), .B1(new_n589), .B2(new_n636), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n667), .A2(new_n612), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT43), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n765), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n765), .A2(new_n770), .A3(KEYINPUT44), .A4(new_n771), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n743), .A3(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n736), .A2(new_n738), .A3(KEYINPUT45), .A4(new_n740), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(G469), .C1(KEYINPUT45), .C2(new_n537), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n735), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n548), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n701), .B(new_n658), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(KEYINPUT106), .B(G137), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G39));
  OAI21_X1  g601(.A(new_n701), .B1(new_n782), .B2(new_n783), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT47), .Z(new_n789));
  INV_X1    g603(.A(new_n743), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n301), .A2(new_n790), .A3(new_n596), .A4(new_n681), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR2_X1   g607(.A1(G952), .A2(G953), .ZN(new_n794));
  INV_X1    g608(.A(new_n732), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n748), .A2(new_n627), .A3(new_n687), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n549), .A2(new_n654), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n795), .A2(new_n711), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n638), .A2(new_n635), .A3(new_n761), .ZN(new_n799));
  INV_X1    g613(.A(new_n548), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n741), .A2(new_n735), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n701), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT108), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n742), .A2(new_n804), .A3(new_n701), .A4(new_n799), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n714), .B1(new_n672), .B2(new_n677), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n798), .A2(new_n695), .A3(new_n808), .ZN(new_n809));
  XOR2_X1   g623(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n710), .A2(new_n732), .B1(new_n650), .B2(new_n655), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n694), .B2(new_n684), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n806), .B2(new_n807), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n812), .A2(new_n816), .A3(new_n798), .A4(new_n695), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n811), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n723), .A2(new_n725), .A3(new_n665), .A4(new_n726), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n731), .A3(new_n760), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT107), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n486), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT107), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n647), .A2(new_n827), .A3(new_n447), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n743), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n797), .A2(new_n692), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n763), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n449), .A2(new_n450), .A3(new_n826), .A4(new_n825), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n492), .B1(new_n833), .B2(new_n614), .ZN(new_n834));
  INV_X1    g648(.A(new_n381), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n602), .A2(new_n834), .A3(new_n549), .A4(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n597), .A3(new_n643), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n820), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n748), .A2(new_n829), .A3(new_n687), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n755), .A2(new_n762), .B1(new_n839), .B2(new_n797), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n836), .A2(new_n597), .A3(new_n643), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT112), .A4(new_n823), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n838), .A2(new_n842), .A3(KEYINPUT53), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n703), .B1(new_n615), .B2(new_n628), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n712), .A3(new_n728), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT113), .B1(new_n758), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n753), .A2(new_n754), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n756), .A2(new_n757), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  INV_X1    g664(.A(new_n845), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n819), .A2(new_n843), .A3(new_n846), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT53), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n809), .B(KEYINPUT52), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n840), .A2(new_n841), .A3(new_n823), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n849), .A2(new_n858), .A3(new_n851), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n855), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n758), .A2(new_n857), .A3(new_n845), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n814), .A2(KEYINPUT52), .A3(new_n808), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n809), .A2(new_n815), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT111), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n816), .A2(new_n798), .A3(new_n695), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(KEYINPUT109), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n814), .A2(new_n812), .A3(new_n816), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(new_n809), .B2(new_n810), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n855), .B1(new_n871), .B2(new_n859), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT111), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n862), .A2(new_n865), .A3(new_n873), .A4(KEYINPUT53), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n867), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n861), .B1(KEYINPUT54), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n702), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n489), .A3(new_n743), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n770), .A2(new_n771), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n749), .A2(new_n750), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n672), .A2(new_n677), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n878), .A2(new_n595), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n668), .A3(new_n612), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n770), .A2(new_n489), .A3(new_n771), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n727), .A2(new_n596), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n488), .B1(new_n889), .B2(new_n711), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n880), .A2(new_n821), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n668), .A2(new_n612), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n885), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n664), .A2(new_n877), .A3(new_n619), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT114), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n889), .A2(new_n743), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n788), .B(KEYINPUT47), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n700), .A2(new_n548), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n701), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n899), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n894), .A2(new_n908), .A3(new_n898), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n910), .B2(new_n905), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n891), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n794), .B1(new_n876), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n902), .B(KEYINPUT49), .Z(new_n914));
  NAND3_X1  g728(.A1(new_n596), .A2(new_n701), .A3(new_n379), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n884), .A2(new_n766), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n916), .A3(new_n664), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT115), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n862), .B2(new_n865), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n843), .A2(new_n852), .A3(new_n846), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n819), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n854), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n924), .A3(new_n912), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(G952), .B2(G953), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n927), .A3(new_n917), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n919), .A2(new_n928), .ZN(G75));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n853), .A2(new_n860), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(G210), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n339), .A2(new_n352), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT116), .Z(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT55), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT117), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n350), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n934), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n934), .A2(new_n940), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n487), .A2(G952), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G51));
  NAND2_X1  g758(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n924), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n735), .B(KEYINPUT118), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT57), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n544), .A3(new_n547), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n932), .A2(new_n778), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n943), .B1(new_n950), .B2(new_n951), .ZN(G54));
  NAND4_X1  g766(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n439), .A2(new_n440), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n943), .ZN(G60));
  XOR2_X1   g771(.A(new_n609), .B(KEYINPUT59), .Z(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n920), .B2(new_n924), .ZN(new_n959));
  INV_X1    g773(.A(new_n611), .ZN(new_n960));
  OAI21_X1  g774(.A(KEYINPUT119), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n611), .C1(new_n876), .C2(new_n958), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n611), .A2(new_n958), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n943), .B1(new_n946), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(G63));
  INV_X1    g780(.A(KEYINPUT120), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n923), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n931), .A2(KEYINPUT120), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n584), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n633), .A2(new_n634), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT120), .B1(new_n931), .B2(new_n971), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n967), .B(new_n969), .C1(new_n853), .C2(new_n860), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n943), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n973), .A2(new_n977), .A3(KEYINPUT61), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  INV_X1    g797(.A(new_n491), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n487), .B1(new_n984), .B2(G224), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n845), .A2(new_n837), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT121), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(new_n487), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n936), .B1(G898), .B2(new_n487), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT122), .Z(new_n990));
  XNOR2_X1  g804(.A(new_n988), .B(new_n990), .ZN(G69));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n814), .B(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n679), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n833), .A2(new_n614), .ZN(new_n997));
  OR4_X1    g811(.A1(new_n698), .A2(new_n660), .A3(new_n790), .A4(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n792), .A2(new_n785), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n995), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n487), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n391), .A2(new_n394), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n266), .B(new_n1002), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n763), .B1(new_n776), .B2(new_n784), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n784), .A2(new_n714), .A3(new_n881), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n792), .A2(new_n1006), .A3(new_n993), .A4(new_n849), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(G953), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1009));
  AOI22_X1  g823(.A1(new_n1001), .A2(new_n1003), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n487), .B1(G227), .B2(G900), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1010), .B(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n1007), .B2(new_n987), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n292), .A2(new_n253), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(KEYINPUT124), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n943), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT125), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1015), .B1(new_n1000), .B2(new_n987), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1021), .A2(new_n674), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1017), .A2(new_n673), .A3(new_n1015), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT126), .Z(new_n1024));
  NAND2_X1  g838(.A1(new_n875), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT127), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1020), .A2(new_n1022), .A3(new_n1027), .ZN(G57));
endmodule


