

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U560 ( .A(n621), .B(KEYINPUT26), .ZN(n632) );
  NOR2_X1 U561 ( .A1(G164), .A2(G1384), .ZN(n732) );
  INV_X1 U562 ( .A(KEYINPUT66), .ZN(n526) );
  OR2_X1 U563 ( .A1(n714), .A2(n713), .ZN(n748) );
  NAND2_X1 U564 ( .A1(n870), .A2(G114), .ZN(n528) );
  NOR2_X1 U565 ( .A1(n536), .A2(n535), .ZN(G164) );
  NAND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X2 U567 ( .A(n527), .B(n526), .ZN(n870) );
  XNOR2_X1 U568 ( .A(n528), .B(KEYINPUT97), .ZN(n536) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n529), .Z(n874) );
  NAND2_X1 U571 ( .A1(n874), .A2(G138), .ZN(n534) );
  INV_X1 U572 ( .A(G2105), .ZN(n530) );
  AND2_X1 U573 ( .A1(n530), .A2(G2104), .ZN(n873) );
  NAND2_X1 U574 ( .A1(G102), .A2(n873), .ZN(n532) );
  NOR2_X1 U575 ( .A1(G2104), .A2(n530), .ZN(n869) );
  NAND2_X1 U576 ( .A1(G126), .A2(n869), .ZN(n531) );
  AND2_X1 U577 ( .A1(n532), .A2(n531), .ZN(n533) );
  NAND2_X1 U578 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U579 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n538) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n593) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(G651), .ZN(n539) );
  NOR2_X1 U582 ( .A1(n593), .A2(n539), .ZN(n805) );
  NAND2_X1 U583 ( .A1(G73), .A2(n805), .ZN(n537) );
  XNOR2_X1 U584 ( .A(n538), .B(n537), .ZN(n549) );
  XNOR2_X1 U585 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n542) );
  NOR2_X1 U586 ( .A1(G543), .A2(n539), .ZN(n540) );
  XNOR2_X1 U587 ( .A(n540), .B(KEYINPUT1), .ZN(n541) );
  XNOR2_X1 U588 ( .A(n542), .B(n541), .ZN(n800) );
  NAND2_X1 U589 ( .A1(G61), .A2(n800), .ZN(n544) );
  NOR2_X1 U590 ( .A1(n593), .A2(G651), .ZN(n801) );
  NAND2_X1 U591 ( .A1(G48), .A2(n801), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n544), .A2(n543), .ZN(n547) );
  NOR2_X1 U593 ( .A1(G543), .A2(G651), .ZN(n804) );
  NAND2_X1 U594 ( .A1(n804), .A2(G86), .ZN(n545) );
  XOR2_X1 U595 ( .A(KEYINPUT86), .B(n545), .Z(n546) );
  NOR2_X1 U596 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n549), .A2(n548), .ZN(G305) );
  NAND2_X1 U598 ( .A1(n804), .A2(G89), .ZN(n550) );
  XNOR2_X1 U599 ( .A(KEYINPUT4), .B(n550), .ZN(n553) );
  NAND2_X1 U600 ( .A1(G76), .A2(n805), .ZN(n551) );
  XOR2_X1 U601 ( .A(KEYINPUT79), .B(n551), .Z(n552) );
  NAND2_X1 U602 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U603 ( .A(n554), .B(KEYINPUT5), .ZN(n559) );
  NAND2_X1 U604 ( .A1(G63), .A2(n800), .ZN(n556) );
  NAND2_X1 U605 ( .A1(G51), .A2(n801), .ZN(n555) );
  NAND2_X1 U606 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n557), .Z(n558) );
  NAND2_X1 U608 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U609 ( .A(n560), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U610 ( .A1(n874), .A2(G137), .ZN(n563) );
  NAND2_X1 U611 ( .A1(G101), .A2(n873), .ZN(n561) );
  XOR2_X1 U612 ( .A(KEYINPUT23), .B(n561), .Z(n562) );
  NAND2_X1 U613 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U614 ( .A1(n869), .A2(G125), .ZN(n565) );
  NAND2_X1 U615 ( .A1(G113), .A2(n870), .ZN(n564) );
  NAND2_X1 U616 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U617 ( .A1(n567), .A2(n566), .ZN(G160) );
  NAND2_X1 U618 ( .A1(G64), .A2(n800), .ZN(n569) );
  NAND2_X1 U619 ( .A1(G52), .A2(n801), .ZN(n568) );
  NAND2_X1 U620 ( .A1(n569), .A2(n568), .ZN(n575) );
  NAND2_X1 U621 ( .A1(G90), .A2(n804), .ZN(n571) );
  NAND2_X1 U622 ( .A1(G77), .A2(n805), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U624 ( .A(KEYINPUT70), .B(n572), .Z(n573) );
  XNOR2_X1 U625 ( .A(KEYINPUT9), .B(n573), .ZN(n574) );
  NOR2_X1 U626 ( .A1(n575), .A2(n574), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G53), .A2(n801), .ZN(n576) );
  XNOR2_X1 U628 ( .A(n576), .B(KEYINPUT72), .ZN(n583) );
  NAND2_X1 U629 ( .A1(G65), .A2(n800), .ZN(n578) );
  NAND2_X1 U630 ( .A1(G91), .A2(n804), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U632 ( .A1(G78), .A2(n805), .ZN(n579) );
  XNOR2_X1 U633 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U635 ( .A1(n583), .A2(n582), .ZN(G299) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G75), .A2(n805), .ZN(n590) );
  NAND2_X1 U638 ( .A1(G62), .A2(n800), .ZN(n585) );
  NAND2_X1 U639 ( .A1(G50), .A2(n801), .ZN(n584) );
  NAND2_X1 U640 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U641 ( .A1(n804), .A2(G88), .ZN(n586) );
  XOR2_X1 U642 ( .A(KEYINPUT88), .B(n586), .Z(n587) );
  NOR2_X1 U643 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U644 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U645 ( .A(KEYINPUT89), .B(n591), .ZN(G166) );
  INV_X1 U646 ( .A(G166), .ZN(G303) );
  NAND2_X1 U647 ( .A1(G49), .A2(n801), .ZN(n592) );
  XNOR2_X1 U648 ( .A(n592), .B(KEYINPUT84), .ZN(n596) );
  NAND2_X1 U649 ( .A1(G87), .A2(n593), .ZN(n594) );
  XOR2_X1 U650 ( .A(KEYINPUT85), .B(n594), .Z(n595) );
  NAND2_X1 U651 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U652 ( .A1(n800), .A2(n597), .ZN(n599) );
  NAND2_X1 U653 ( .A1(G651), .A2(G74), .ZN(n598) );
  NAND2_X1 U654 ( .A1(n599), .A2(n598), .ZN(G288) );
  NAND2_X1 U655 ( .A1(G60), .A2(n800), .ZN(n601) );
  NAND2_X1 U656 ( .A1(G47), .A2(n801), .ZN(n600) );
  NAND2_X1 U657 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U658 ( .A1(G85), .A2(n804), .ZN(n603) );
  NAND2_X1 U659 ( .A1(G72), .A2(n805), .ZN(n602) );
  NAND2_X1 U660 ( .A1(n603), .A2(n602), .ZN(n604) );
  OR2_X1 U661 ( .A1(n605), .A2(n604), .ZN(G290) );
  XOR2_X1 U662 ( .A(G1981), .B(G305), .Z(n978) );
  NAND2_X1 U663 ( .A1(G160), .A2(G40), .ZN(n731) );
  INV_X1 U664 ( .A(n731), .ZN(n606) );
  NAND2_X1 U665 ( .A1(n606), .A2(n732), .ZN(n608) );
  INV_X1 U666 ( .A(KEYINPUT64), .ZN(n607) );
  XNOR2_X1 U667 ( .A(n608), .B(n607), .ZN(n620) );
  INV_X1 U668 ( .A(n620), .ZN(n618) );
  INV_X1 U669 ( .A(n618), .ZN(n655) );
  INV_X1 U670 ( .A(n655), .ZN(n672) );
  NAND2_X1 U671 ( .A1(n672), .A2(G8), .ZN(n712) );
  NOR2_X1 U672 ( .A1(G1966), .A2(n712), .ZN(n684) );
  NOR2_X1 U673 ( .A1(n618), .A2(G2084), .ZN(n609) );
  XNOR2_X1 U674 ( .A(KEYINPUT103), .B(n609), .ZN(n681) );
  NAND2_X1 U675 ( .A1(G8), .A2(n681), .ZN(n610) );
  NOR2_X1 U676 ( .A1(n684), .A2(n610), .ZN(n611) );
  XOR2_X1 U677 ( .A(KEYINPUT30), .B(n611), .Z(n612) );
  NOR2_X1 U678 ( .A1(G168), .A2(n612), .ZN(n616) );
  XNOR2_X1 U679 ( .A(G2078), .B(KEYINPUT25), .ZN(n960) );
  NAND2_X1 U680 ( .A1(n655), .A2(n960), .ZN(n614) );
  INV_X1 U681 ( .A(G1961), .ZN(n981) );
  NAND2_X1 U682 ( .A1(n672), .A2(n981), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n666) );
  NOR2_X1 U684 ( .A1(G171), .A2(n666), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(KEYINPUT31), .B(n617), .ZN(n670) );
  NAND2_X1 U687 ( .A1(n618), .A2(G1341), .ZN(n619) );
  XNOR2_X1 U688 ( .A(KEYINPUT105), .B(n619), .ZN(n634) );
  NAND2_X1 U689 ( .A1(n620), .A2(G1996), .ZN(n621) );
  NAND2_X1 U690 ( .A1(G43), .A2(n801), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT74), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G56), .A2(n800), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(KEYINPUT14), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n631) );
  NAND2_X1 U695 ( .A1(n804), .A2(G81), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n626), .B(KEYINPUT12), .ZN(n628) );
  NAND2_X1 U697 ( .A1(G68), .A2(n805), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U699 ( .A(KEYINPUT13), .B(n629), .Z(n630) );
  NOR2_X1 U700 ( .A1(n631), .A2(n630), .ZN(n778) );
  NAND2_X1 U701 ( .A1(n632), .A2(n778), .ZN(n633) );
  OR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U703 ( .A(n635), .B(KEYINPUT65), .ZN(n649) );
  NAND2_X1 U704 ( .A1(n805), .A2(G79), .ZN(n642) );
  NAND2_X1 U705 ( .A1(G66), .A2(n800), .ZN(n637) );
  NAND2_X1 U706 ( .A1(G92), .A2(n804), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U708 ( .A1(G54), .A2(n801), .ZN(n638) );
  XNOR2_X1 U709 ( .A(KEYINPUT77), .B(n638), .ZN(n639) );
  NOR2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n643), .B(KEYINPUT15), .ZN(n989) );
  NAND2_X1 U713 ( .A1(n649), .A2(n989), .ZN(n647) );
  NOR2_X1 U714 ( .A1(n672), .A2(G2067), .ZN(n645) );
  NOR2_X1 U715 ( .A1(G1348), .A2(n655), .ZN(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n648), .B(KEYINPUT106), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n989), .A2(n649), .ZN(n650) );
  XNOR2_X1 U720 ( .A(KEYINPUT107), .B(n650), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n652), .A2(n651), .ZN(n659) );
  INV_X1 U722 ( .A(G299), .ZN(n818) );
  NAND2_X1 U723 ( .A1(n655), .A2(G2072), .ZN(n654) );
  XNOR2_X1 U724 ( .A(KEYINPUT27), .B(KEYINPUT104), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n657) );
  INV_X1 U726 ( .A(G1956), .ZN(n910) );
  NOR2_X1 U727 ( .A1(n655), .A2(n910), .ZN(n656) );
  NOR2_X1 U728 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n818), .A2(n660), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n818), .A2(n660), .ZN(n661) );
  XOR2_X1 U732 ( .A(n661), .B(KEYINPUT28), .Z(n662) );
  NAND2_X1 U733 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U734 ( .A(KEYINPUT29), .B(KEYINPUT108), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n665), .B(n664), .ZN(n668) );
  AND2_X1 U736 ( .A1(n666), .A2(G171), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n683) );
  INV_X1 U739 ( .A(n683), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(G286), .ZN(n677) );
  NOR2_X1 U741 ( .A1(n672), .A2(G2090), .ZN(n674) );
  NOR2_X1 U742 ( .A1(G1971), .A2(n712), .ZN(n673) );
  NOR2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U744 ( .A1(G303), .A2(n675), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n678), .A2(G8), .ZN(n680) );
  XNOR2_X1 U747 ( .A(KEYINPUT110), .B(KEYINPUT32), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(n679), .ZN(n690) );
  INV_X1 U749 ( .A(n681), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n682), .A2(G8), .ZN(n688) );
  INV_X1 U751 ( .A(KEYINPUT109), .ZN(n686) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U753 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n705) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n985) );
  XOR2_X1 U758 ( .A(n985), .B(KEYINPUT111), .Z(n691) );
  NOR2_X1 U759 ( .A1(n986), .A2(n691), .ZN(n693) );
  INV_X1 U760 ( .A(KEYINPUT33), .ZN(n692) );
  AND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U762 ( .A1(n705), .A2(n694), .ZN(n698) );
  NAND2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U764 ( .A(n987), .ZN(n695) );
  NOR2_X1 U765 ( .A1(n712), .A2(n695), .ZN(n696) );
  OR2_X1 U766 ( .A1(KEYINPUT33), .A2(n696), .ZN(n697) );
  NAND2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n986), .A2(KEYINPUT33), .ZN(n699) );
  NOR2_X1 U769 ( .A1(n699), .A2(n712), .ZN(n700) );
  NOR2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n978), .A2(n702), .ZN(n709) );
  NOR2_X1 U772 ( .A1(G2090), .A2(G303), .ZN(n703) );
  NAND2_X1 U773 ( .A1(G8), .A2(n703), .ZN(n704) );
  NAND2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n706), .B(KEYINPUT112), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n707), .A2(n712), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n714) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n710) );
  XOR2_X1 U779 ( .A(n710), .B(KEYINPUT24), .Z(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U781 ( .A1(n873), .A2(G105), .ZN(n716) );
  XNOR2_X1 U782 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n715) );
  XNOR2_X1 U783 ( .A(n716), .B(n715), .ZN(n723) );
  NAND2_X1 U784 ( .A1(G141), .A2(n874), .ZN(n718) );
  NAND2_X1 U785 ( .A1(G117), .A2(n870), .ZN(n717) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U787 ( .A1(G129), .A2(n869), .ZN(n719) );
  XNOR2_X1 U788 ( .A(KEYINPUT101), .B(n719), .ZN(n720) );
  NOR2_X1 U789 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n882) );
  AND2_X1 U791 ( .A1(n882), .A2(G1996), .ZN(n935) );
  NAND2_X1 U792 ( .A1(G119), .A2(n869), .ZN(n724) );
  XNOR2_X1 U793 ( .A(n724), .B(KEYINPUT100), .ZN(n726) );
  NAND2_X1 U794 ( .A1(n874), .A2(G131), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U796 ( .A1(G95), .A2(n873), .ZN(n728) );
  NAND2_X1 U797 ( .A1(G107), .A2(n870), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n881) );
  INV_X1 U800 ( .A(G1991), .ZN(n914) );
  NOR2_X1 U801 ( .A1(n881), .A2(n914), .ZN(n937) );
  OR2_X1 U802 ( .A1(n935), .A2(n937), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n732), .A2(n731), .ZN(n760) );
  AND2_X1 U804 ( .A1(n733), .A2(n760), .ZN(n752) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n995) );
  NAND2_X1 U806 ( .A1(n995), .A2(n760), .ZN(n734) );
  XNOR2_X1 U807 ( .A(n734), .B(KEYINPUT98), .ZN(n745) );
  XNOR2_X1 U808 ( .A(G2067), .B(KEYINPUT37), .ZN(n757) );
  NAND2_X1 U809 ( .A1(G104), .A2(n873), .ZN(n736) );
  NAND2_X1 U810 ( .A1(G140), .A2(n874), .ZN(n735) );
  NAND2_X1 U811 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U812 ( .A(KEYINPUT34), .B(n737), .ZN(n743) );
  NAND2_X1 U813 ( .A1(G116), .A2(n870), .ZN(n738) );
  XOR2_X1 U814 ( .A(KEYINPUT99), .B(n738), .Z(n740) );
  NAND2_X1 U815 ( .A1(n869), .A2(G128), .ZN(n739) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U817 ( .A(KEYINPUT35), .B(n741), .Z(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U819 ( .A(KEYINPUT36), .B(n744), .ZN(n890) );
  NOR2_X1 U820 ( .A1(n757), .A2(n890), .ZN(n953) );
  NAND2_X1 U821 ( .A1(n760), .A2(n953), .ZN(n755) );
  NAND2_X1 U822 ( .A1(n745), .A2(n755), .ZN(n746) );
  NOR2_X1 U823 ( .A1(n752), .A2(n746), .ZN(n747) );
  NAND2_X1 U824 ( .A1(n748), .A2(n747), .ZN(n763) );
  NOR2_X1 U825 ( .A1(G1996), .A2(n882), .ZN(n932) );
  AND2_X1 U826 ( .A1(n914), .A2(n881), .ZN(n936) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n749) );
  XOR2_X1 U828 ( .A(n749), .B(KEYINPUT113), .Z(n750) );
  NOR2_X1 U829 ( .A1(n936), .A2(n750), .ZN(n751) );
  NOR2_X1 U830 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U831 ( .A1(n932), .A2(n753), .ZN(n754) );
  XNOR2_X1 U832 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U833 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U834 ( .A1(n757), .A2(n890), .ZN(n950) );
  NAND2_X1 U835 ( .A1(n758), .A2(n950), .ZN(n759) );
  NAND2_X1 U836 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U837 ( .A(n761), .B(KEYINPUT114), .ZN(n762) );
  NAND2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U839 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U840 ( .A(G2435), .B(G2454), .Z(n766) );
  XNOR2_X1 U841 ( .A(KEYINPUT115), .B(G2438), .ZN(n765) );
  XNOR2_X1 U842 ( .A(n766), .B(n765), .ZN(n773) );
  XOR2_X1 U843 ( .A(G2446), .B(G2430), .Z(n768) );
  XNOR2_X1 U844 ( .A(G2451), .B(G2443), .ZN(n767) );
  XNOR2_X1 U845 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U846 ( .A(n769), .B(G2427), .Z(n771) );
  XNOR2_X1 U847 ( .A(G1341), .B(G1348), .ZN(n770) );
  XNOR2_X1 U848 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U849 ( .A(n773), .B(n772), .ZN(n774) );
  AND2_X1 U850 ( .A1(n774), .A2(G14), .ZN(G401) );
  AND2_X1 U851 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U852 ( .A(G108), .ZN(G238) );
  INV_X1 U853 ( .A(G120), .ZN(G236) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  INV_X1 U856 ( .A(G82), .ZN(G220) );
  XOR2_X1 U857 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n776) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n775) );
  XOR2_X1 U859 ( .A(n776), .B(n775), .Z(n846) );
  INV_X1 U860 ( .A(n846), .ZN(G223) );
  INV_X1 U861 ( .A(G567), .ZN(n841) );
  NOR2_X1 U862 ( .A1(n841), .A2(G223), .ZN(n777) );
  XNOR2_X1 U863 ( .A(n777), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U864 ( .A(n778), .ZN(n998) );
  XNOR2_X1 U865 ( .A(G860), .B(KEYINPUT75), .ZN(n786) );
  OR2_X1 U866 ( .A1(n998), .A2(n786), .ZN(G153) );
  XOR2_X1 U867 ( .A(KEYINPUT76), .B(G171), .Z(G301) );
  INV_X1 U868 ( .A(G868), .ZN(n824) );
  NOR2_X1 U869 ( .A1(G301), .A2(n824), .ZN(n780) );
  AND2_X1 U870 ( .A1(n824), .A2(n989), .ZN(n779) );
  NOR2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U872 ( .A(KEYINPUT78), .B(n781), .ZN(G284) );
  NOR2_X1 U873 ( .A1(G286), .A2(n824), .ZN(n782) );
  XNOR2_X1 U874 ( .A(n782), .B(KEYINPUT80), .ZN(n784) );
  NOR2_X1 U875 ( .A1(G299), .A2(G868), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U877 ( .A(KEYINPUT81), .B(n785), .Z(G297) );
  NAND2_X1 U878 ( .A1(n786), .A2(G559), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n787), .A2(n989), .ZN(n788) );
  XNOR2_X1 U880 ( .A(n788), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U881 ( .A1(n989), .A2(G868), .ZN(n789) );
  NOR2_X1 U882 ( .A1(G559), .A2(n789), .ZN(n791) );
  NOR2_X1 U883 ( .A1(G868), .A2(n998), .ZN(n790) );
  NOR2_X1 U884 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U885 ( .A1(G123), .A2(n869), .ZN(n792) );
  XNOR2_X1 U886 ( .A(n792), .B(KEYINPUT18), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n873), .A2(G99), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G135), .A2(n874), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G111), .A2(n870), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n934) );
  XNOR2_X1 U893 ( .A(G2096), .B(n934), .ZN(n799) );
  INV_X1 U894 ( .A(G2100), .ZN(n905) );
  NAND2_X1 U895 ( .A1(n799), .A2(n905), .ZN(G156) );
  NAND2_X1 U896 ( .A1(G67), .A2(n800), .ZN(n803) );
  NAND2_X1 U897 ( .A1(G55), .A2(n801), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G93), .A2(n804), .ZN(n807) );
  NAND2_X1 U900 ( .A1(G80), .A2(n805), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  OR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n823) );
  XNOR2_X1 U903 ( .A(n998), .B(KEYINPUT82), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G559), .A2(n989), .ZN(n810) );
  XNOR2_X1 U905 ( .A(n811), .B(n810), .ZN(n821) );
  XOR2_X1 U906 ( .A(n821), .B(KEYINPUT83), .Z(n812) );
  NOR2_X1 U907 ( .A1(G860), .A2(n812), .ZN(n813) );
  XOR2_X1 U908 ( .A(n823), .B(n813), .Z(G145) );
  XOR2_X1 U909 ( .A(n823), .B(G290), .Z(n816) );
  XNOR2_X1 U910 ( .A(KEYINPUT90), .B(KEYINPUT19), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n814), .B(G288), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U913 ( .A(G305), .B(n817), .ZN(n820) );
  XOR2_X1 U914 ( .A(G303), .B(n818), .Z(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n896) );
  XNOR2_X1 U916 ( .A(n821), .B(n896), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n822), .A2(G868), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n826), .A2(n825), .ZN(G295) );
  NAND2_X1 U920 ( .A1(G2078), .A2(G2084), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT91), .B(KEYINPUT20), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT92), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(G2090), .ZN(n832) );
  XOR2_X1 U925 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n831) );
  XNOR2_X1 U926 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U927 ( .A1(n833), .A2(G2072), .ZN(n834) );
  XNOR2_X1 U928 ( .A(n834), .B(KEYINPUT94), .ZN(G158) );
  XNOR2_X1 U929 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U930 ( .A1(G220), .A2(G219), .ZN(n835) );
  XOR2_X1 U931 ( .A(KEYINPUT22), .B(n835), .Z(n836) );
  NOR2_X1 U932 ( .A1(G218), .A2(n836), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G96), .A2(n837), .ZN(n852) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n852), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n838), .B(KEYINPUT95), .ZN(n843) );
  NOR2_X1 U936 ( .A1(G236), .A2(G238), .ZN(n839) );
  NAND2_X1 U937 ( .A1(G69), .A2(n839), .ZN(n840) );
  NOR2_X1 U938 ( .A1(G237), .A2(n840), .ZN(n851) );
  NOR2_X1 U939 ( .A1(n841), .A2(n851), .ZN(n842) );
  NOR2_X1 U940 ( .A1(n843), .A2(n842), .ZN(G319) );
  INV_X1 U941 ( .A(G319), .ZN(n925) );
  NAND2_X1 U942 ( .A1(G483), .A2(G661), .ZN(n844) );
  NOR2_X1 U943 ( .A1(n925), .A2(n844), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G36), .A2(n848), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n845), .B(KEYINPUT96), .ZN(G176) );
  NAND2_X1 U946 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U947 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U950 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n850), .B(KEYINPUT116), .ZN(G188) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(n851), .ZN(n853) );
  NOR2_X1 U955 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  NAND2_X1 U957 ( .A1(G124), .A2(n869), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n873), .A2(G100), .ZN(n855) );
  NAND2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G136), .A2(n874), .ZN(n858) );
  NAND2_X1 U962 ( .A1(G112), .A2(n870), .ZN(n857) );
  NAND2_X1 U963 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U964 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U965 ( .A1(n869), .A2(G127), .ZN(n862) );
  NAND2_X1 U966 ( .A1(G115), .A2(n870), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U968 ( .A(n863), .B(KEYINPUT47), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G139), .A2(n874), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n873), .A2(G103), .ZN(n866) );
  XOR2_X1 U972 ( .A(KEYINPUT120), .B(n866), .Z(n867) );
  NOR2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n944) );
  NAND2_X1 U974 ( .A1(n869), .A2(G130), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G118), .A2(n870), .ZN(n871) );
  NAND2_X1 U976 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT45), .B(n877), .Z(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n944), .B(n880), .ZN(n886) );
  XOR2_X1 U983 ( .A(G162), .B(n881), .Z(n884) );
  XOR2_X1 U984 ( .A(G160), .B(n882), .Z(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n886), .B(n885), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n888) );
  XNOR2_X1 U988 ( .A(G164), .B(n934), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U992 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U993 ( .A(KEYINPUT121), .B(n998), .ZN(n895) );
  XNOR2_X1 U994 ( .A(G171), .B(n989), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n898) );
  XNOR2_X1 U996 ( .A(G286), .B(n896), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U998 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U999 ( .A(KEYINPUT42), .B(G2084), .Z(n901) );
  XNOR2_X1 U1000 ( .A(G2090), .B(G2078), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1002 ( .A(n902), .B(G2096), .Z(n904) );
  XNOR2_X1 U1003 ( .A(G2067), .B(G2072), .ZN(n903) );
  XNOR2_X1 U1004 ( .A(n904), .B(n903), .ZN(n909) );
  XOR2_X1 U1005 ( .A(KEYINPUT43), .B(G2678), .Z(n907) );
  XOR2_X1 U1006 ( .A(KEYINPUT117), .B(n905), .Z(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1008 ( .A(n909), .B(n908), .Z(G227) );
  XOR2_X1 U1009 ( .A(KEYINPUT118), .B(G1986), .Z(n912) );
  XOR2_X1 U1010 ( .A(G1971), .B(n910), .Z(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n913), .B(KEYINPUT41), .Z(n916) );
  XOR2_X1 U1013 ( .A(G1996), .B(n914), .Z(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n920) );
  XOR2_X1 U1015 ( .A(G1976), .B(G1981), .Z(n918) );
  XOR2_X1 U1016 ( .A(n981), .B(G1966), .Z(n917) );
  XNOR2_X1 U1017 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(n920), .B(n919), .Z(n922) );
  XNOR2_X1 U1019 ( .A(KEYINPUT119), .B(G2474), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(G229) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(G397), .A2(n924), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(G401), .A2(n925), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT122), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(G395), .A2(n929), .ZN(n930) );
  XOR2_X1 U1028 ( .A(KEYINPUT123), .B(n930), .Z(G308) );
  INV_X1 U1029 ( .A(G308), .ZN(G225) );
  INV_X1 U1030 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n933), .Z(n943) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n941) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1040 ( .A(G2072), .B(n944), .Z(n946) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1043 ( .A(KEYINPUT50), .B(n947), .Z(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n951) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n974), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n966) );
  XOR2_X1 U1054 ( .A(G25), .B(G1991), .Z(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(G28), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G1996), .B(G32), .Z(n962) );
  XNOR2_X1 U1057 ( .A(n960), .B(G27), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(KEYINPUT53), .ZN(n970) );
  XOR2_X1 U1062 ( .A(G2084), .B(KEYINPUT54), .Z(n968) );
  XNOR2_X1 U1063 ( .A(G34), .B(n968), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G35), .B(G2090), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n974), .B(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(G29), .A2(n975), .ZN(n976) );
  XOR2_X1 U1069 ( .A(KEYINPUT124), .B(n976), .Z(n977) );
  NAND2_X1 U1070 ( .A1(G11), .A2(n977), .ZN(n1033) );
  INV_X1 U1071 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1072 ( .A(n1029), .B(KEYINPUT56), .Z(n1004) );
  XNOR2_X1 U1073 ( .A(G168), .B(G1966), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT57), .ZN(n1002) );
  XOR2_X1 U1076 ( .A(G299), .B(G1956), .Z(n983) );
  XOR2_X1 U1077 ( .A(G171), .B(n981), .Z(n982) );
  NAND2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n997) );
  INV_X1 U1080 ( .A(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1082 ( .A(n989), .B(G1348), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n998), .B(G1341), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  XOR2_X1 U1092 ( .A(G5), .B(G1961), .Z(n1016) );
  XOR2_X1 U1093 ( .A(G20), .B(G1956), .Z(n1008) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT59), .B(G1348), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT60), .B(n1012), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1026) );
  XNOR2_X1 U1105 ( .A(KEYINPUT125), .B(G1971), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G1976), .B(KEYINPUT126), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(G23), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G24), .B(G1986), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1023), .Z(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .ZN(G150) );
  INV_X1 U1121 ( .A(G150), .ZN(G311) );
endmodule

