//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G131), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G137), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n192), .A4(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G134), .ZN(new_n196));
  OAI21_X1  g010(.A(G131), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  OAI211_X1 g017(.A(G128), .B(new_n200), .C1(new_n201), .C2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n206), .C1(KEYINPUT1), .C2(new_n207), .ZN(new_n208));
  AND3_X1   g022(.A1(new_n204), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(KEYINPUT67), .B1(new_n204), .B2(new_n208), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n198), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n194), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n206), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  XNOR2_X1  g031(.A(G143), .B(G146), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT0), .B(G128), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n222), .B(new_n223), .C1(new_n201), .C2(new_n203), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n217), .B1(new_n224), .B2(new_n216), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n214), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n227));
  INV_X1    g041(.A(G113), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT65), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n230), .B1(KEYINPUT2), .B2(G113), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n231), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  XNOR2_X1  g046(.A(G116), .B(G119), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n231), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n235), .A2(new_n236), .A3(new_n233), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n211), .A2(new_n226), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT28), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n239), .A2(KEYINPUT72), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT72), .B1(new_n239), .B2(new_n240), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n204), .A2(new_n208), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n204), .A2(KEYINPUT67), .A3(new_n208), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n220), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n248), .A2(new_n198), .B1(new_n251), .B2(new_n214), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(new_n238), .ZN(new_n253));
  INV_X1    g067(.A(new_n239), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n243), .B1(new_n240), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n257));
  XOR2_X1   g071(.A(KEYINPUT26), .B(G101), .Z(new_n258));
  NOR2_X1   g072(.A1(G237), .A2(G953), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G210), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NOR3_X1   g077(.A1(new_n256), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G902), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n266));
  INV_X1    g080(.A(new_n249), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n214), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n204), .A2(new_n208), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n198), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n238), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n252), .B2(new_n238), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n266), .B1(new_n272), .B2(new_n240), .ZN(new_n273));
  INV_X1    g087(.A(new_n238), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n249), .B1(new_n194), .B2(new_n213), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n194), .A2(new_n204), .A3(new_n197), .A4(new_n208), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n240), .B1(new_n239), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT71), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n243), .A2(new_n273), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n280), .B2(new_n263), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n275), .B2(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT64), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT64), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n285), .B(new_n282), .C1(new_n275), .C2(new_n276), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n252), .B2(KEYINPUT30), .ZN(new_n289));
  AND4_X1   g103(.A1(new_n288), .A2(new_n211), .A3(new_n226), .A4(KEYINPUT30), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n274), .B(new_n287), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n239), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n263), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n281), .A2(new_n257), .A3(new_n293), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n280), .A2(KEYINPUT74), .A3(new_n263), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n265), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n239), .A2(new_n240), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n239), .A2(KEYINPUT72), .A3(new_n240), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n302), .B(new_n303), .C1(KEYINPUT71), .C2(new_n278), .ZN(new_n304));
  INV_X1    g118(.A(new_n279), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n263), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI211_X1 g122(.A(KEYINPUT73), .B(new_n263), .C1(new_n304), .C2(new_n305), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n263), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n291), .A2(new_n239), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT31), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n291), .A2(new_n239), .A3(new_n311), .A4(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT32), .B(new_n299), .C1(new_n310), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT32), .ZN(new_n318));
  INV_X1    g132(.A(new_n309), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT73), .B1(new_n280), .B2(new_n263), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n313), .B(new_n315), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n321), .B2(new_n298), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n297), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(KEYINPUT78), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n327), .A2(KEYINPUT78), .A3(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n326), .B1(new_n331), .B2(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT16), .ZN(new_n333));
  AOI211_X1 g147(.A(KEYINPUT79), .B(new_n333), .C1(new_n329), .C2(new_n330), .ZN(new_n334));
  OAI21_X1  g148(.A(G146), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n326), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n327), .A2(KEYINPUT78), .A3(G140), .ZN(new_n337));
  XNOR2_X1  g151(.A(G125), .B(G140), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT78), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n339), .B2(new_n333), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n331), .A2(new_n341), .A3(KEYINPUT16), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n202), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT24), .B(G110), .Z(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(KEYINPUT75), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n207), .A2(G119), .ZN(new_n347));
  INV_X1    g161(.A(G119), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G110), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT77), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g175(.A1(KEYINPUT76), .A2(new_n355), .B1(new_n348), .B2(G128), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n359), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n354), .B1(new_n365), .B2(new_n347), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n344), .B(new_n351), .C1(new_n352), .C2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n366), .B2(new_n352), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n363), .B1(new_n362), .B2(new_n359), .ZN(new_n369));
  AND4_X1   g183(.A1(new_n363), .A2(new_n349), .A3(new_n359), .A4(new_n356), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n347), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(KEYINPUT80), .A3(new_n352), .A4(new_n353), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n346), .A2(new_n350), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n335), .A2(KEYINPUT81), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n340), .A2(new_n342), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT81), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n338), .A2(new_n202), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n367), .B1(new_n375), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G137), .ZN(new_n383));
  INV_X1    g197(.A(G953), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n384), .A2(G221), .A3(G234), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n383), .B(new_n385), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n367), .B(new_n386), .C1(new_n375), .C2(new_n381), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(KEYINPUT25), .A3(new_n389), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G217), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(G234), .B2(new_n389), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n388), .A2(new_n390), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(G902), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n233), .A2(KEYINPUT5), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n348), .A2(G116), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n404), .B(G113), .C1(KEYINPUT5), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(G104), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT83), .B1(new_n410), .B2(G107), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT83), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n408), .A3(G104), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(KEYINPUT84), .A3(G107), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n409), .A2(new_n411), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n232), .A2(new_n233), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n408), .A2(G104), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT3), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n410), .B2(G107), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(KEYINPUT3), .A3(G104), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G101), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n406), .A2(new_n416), .A3(new_n417), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n418), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n408), .A2(KEYINPUT3), .A3(G104), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT3), .B1(new_n408), .B2(G104), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT82), .A3(G101), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n422), .B2(new_n423), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n422), .B2(new_n423), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n433), .A3(G101), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n436), .B1(new_n234), .B2(new_n237), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n425), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G110), .B(G122), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n425), .B(new_n439), .C1(new_n435), .C2(new_n437), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(KEYINPUT6), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n267), .A2(G125), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(G125), .B2(new_n244), .ZN(new_n445));
  INV_X1    g259(.A(G224), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(G953), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT85), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n445), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n438), .A2(new_n450), .A3(new_n440), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n443), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n443), .A2(KEYINPUT86), .A3(new_n449), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(new_n446), .B2(G953), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n445), .B(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n406), .A2(new_n417), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n416), .A2(new_n424), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n425), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n439), .B(KEYINPUT8), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n442), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(new_n389), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n456), .A2(new_n457), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n457), .B1(new_n456), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G140), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n384), .A2(G227), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n214), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n430), .A2(new_n432), .A3(new_n434), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n251), .A3(new_n436), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT10), .ZN(new_n477));
  INV_X1    g291(.A(new_n461), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n248), .B2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n461), .A2(KEYINPUT10), .A3(new_n244), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n474), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n477), .A3(new_n269), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n461), .B1(new_n247), .B2(new_n246), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n474), .B1(new_n485), .B2(new_n476), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n473), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n473), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n269), .B1(new_n424), .B2(new_n416), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n461), .A2(new_n244), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n214), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT12), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n493), .B(new_n214), .C1(new_n489), .C2(new_n490), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n481), .A2(new_n488), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n389), .ZN(new_n498));
  NAND2_X1  g312(.A1(G469), .A2(G902), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n481), .A2(new_n492), .A3(new_n494), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n473), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n214), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n481), .A3(new_n488), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(G469), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n498), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G221), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT9), .B(G234), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n507), .B1(new_n509), .B2(new_n389), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(G214), .B1(G237), .B2(G902), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n470), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n517));
  INV_X1    g331(.A(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n384), .A3(G214), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n199), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n517), .B1(new_n522), .B2(G131), .ZN(new_n523));
  AOI211_X1 g337(.A(KEYINPUT89), .B(new_n192), .C1(new_n520), .C2(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT17), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n259), .A2(G143), .A3(G214), .ZN(new_n526));
  AOI21_X1  g340(.A(G143), .B1(new_n259), .B2(G214), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT89), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n517), .A3(G131), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n520), .A2(new_n192), .A3(new_n521), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n335), .A2(new_n525), .A3(new_n533), .A4(new_n343), .ZN(new_n534));
  NAND2_X1  g348(.A1(KEYINPUT18), .A2(G131), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n522), .B(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n338), .B2(new_n202), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n331), .B2(new_n202), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n329), .A2(new_n330), .A3(new_n537), .A4(G146), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT88), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT90), .B(G104), .Z(new_n545));
  XNOR2_X1  g359(.A(G113), .B(G122), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n534), .A2(new_n543), .A3(new_n547), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n516), .B1(new_n551), .B2(new_n389), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT20), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n378), .B1(new_n377), .B2(G146), .ZN(new_n555));
  AOI211_X1 g369(.A(KEYINPUT81), .B(new_n202), .C1(new_n340), .C2(new_n342), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n523), .A2(new_n524), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n331), .A2(KEYINPUT19), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n338), .A2(KEYINPUT19), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n558), .A2(new_n532), .B1(new_n202), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n542), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n539), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n557), .A2(new_n562), .B1(new_n536), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n550), .B1(new_n566), .B2(new_n547), .ZN(new_n567));
  NOR2_X1   g381(.A1(G475), .A2(G902), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n554), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n376), .A3(new_n379), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n547), .B1(new_n570), .B2(new_n543), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n534), .A2(new_n543), .A3(new_n547), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n554), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n553), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G478), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n576), .A2(KEYINPUT15), .ZN(new_n577));
  INV_X1    g391(.A(G122), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(G116), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n408), .B1(new_n579), .B2(KEYINPUT14), .ZN(new_n580));
  XNOR2_X1  g394(.A(G116), .B(G122), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n582), .B2(KEYINPUT14), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n408), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n207), .A2(G143), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n199), .A2(G128), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n188), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n585), .A2(new_n586), .A3(G134), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n583), .B(new_n584), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n585), .B2(KEYINPUT13), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT13), .B1(new_n199), .B2(G128), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n199), .A2(G128), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n593), .A2(new_n591), .A3(new_n594), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(KEYINPUT92), .A3(G134), .A4(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n578), .A2(G116), .ZN(new_n599));
  OAI21_X1  g413(.A(G107), .B1(new_n599), .B2(new_n579), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n589), .B1(new_n600), .B2(new_n584), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n597), .A2(G134), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT92), .B1(new_n603), .B2(new_n596), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n590), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n384), .A2(G217), .ZN(new_n607));
  OR3_X1    g421(.A1(new_n508), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n508), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT94), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n610), .B(new_n590), .C1(new_n602), .C2(new_n604), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(KEYINPUT94), .A3(new_n611), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n577), .B1(new_n616), .B2(new_n389), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n615), .A2(new_n614), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n389), .B(new_n577), .C1(new_n618), .C2(new_n612), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n575), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(G952), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(G953), .ZN(new_n625));
  NAND2_X1  g439(.A1(G234), .A2(G237), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT21), .B(G898), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT96), .Z(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(G902), .A3(G953), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n323), .A2(new_n403), .A3(new_n515), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n321), .B2(new_n389), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n299), .B1(new_n310), .B2(new_n316), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n402), .A2(new_n512), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n513), .B(new_n631), .C1(new_n468), .C2(new_n469), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n614), .A2(KEYINPUT33), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n608), .A2(new_n609), .A3(KEYINPUT98), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT98), .B1(new_n608), .B2(new_n609), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n605), .A2(KEYINPUT99), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT99), .B1(new_n605), .B2(new_n644), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT100), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n641), .B(KEYINPUT100), .C1(new_n645), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n576), .A2(G902), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n616), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT97), .B(new_n653), .C1(new_n618), .C2(new_n612), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n651), .B(new_n652), .C1(new_n654), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n616), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n576), .B1(new_n658), .B2(G902), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n575), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n640), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n638), .A2(new_n639), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  OAI21_X1  g479(.A(new_n568), .B1(new_n571), .B2(new_n572), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT20), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n552), .B1(new_n667), .B2(new_n573), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n622), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n640), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n638), .A2(new_n639), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT101), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  OAI21_X1  g488(.A(new_n382), .B1(KEYINPUT36), .B2(new_n387), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n367), .B(new_n676), .C1(new_n375), .C2(new_n381), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n675), .A2(new_n400), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n675), .A2(KEYINPUT102), .A3(new_n400), .A4(new_n677), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n398), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n683), .A2(new_n631), .A3(new_n623), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n638), .A3(new_n515), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT37), .B(G110), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT103), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G12));
  XOR2_X1   g502(.A(new_n627), .B(KEYINPUT104), .Z(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(G900), .B2(new_n630), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n669), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n456), .A2(new_n467), .ZN(new_n693));
  INV_X1    g507(.A(new_n457), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n456), .A2(new_n457), .A3(new_n467), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n514), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n506), .A2(new_n511), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n697), .A2(new_n698), .A3(new_n683), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n323), .A2(new_n692), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n323), .A2(new_n699), .A3(KEYINPUT105), .A4(new_n692), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  MUX2_X1   g519(.A(new_n255), .B(new_n292), .S(new_n311), .Z(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n706), .B2(G902), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n317), .B2(new_n322), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n690), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n698), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n680), .A2(new_n681), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n397), .B2(new_n395), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n668), .A2(new_n514), .A3(new_n621), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n470), .B(KEYINPUT38), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n719));
  OR4_X1    g533(.A1(new_n709), .A2(new_n717), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  NOR2_X1   g535(.A1(new_n661), .A2(new_n691), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n323), .A2(new_n699), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n488), .B1(new_n503), .B2(new_n481), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n481), .A2(new_n488), .A3(new_n492), .A4(new_n494), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n389), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n498), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n725), .B1(new_n730), .B2(new_n510), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n498), .A3(KEYINPUT107), .A4(new_n511), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n323), .A2(new_n403), .A3(new_n662), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  NAND4_X1  g550(.A1(new_n323), .A2(new_n403), .A3(new_n670), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G116), .ZN(G18));
  AND3_X1   g552(.A1(new_n697), .A2(new_n731), .A3(new_n732), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n323), .A2(new_n684), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND3_X1  g555(.A1(new_n697), .A2(new_n731), .A3(new_n732), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n575), .A2(new_n743), .A3(new_n622), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT108), .B1(new_n668), .B2(new_n621), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n631), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n256), .A2(new_n263), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n299), .B1(new_n316), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n636), .A2(new_n402), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  NOR3_X1   g567(.A1(new_n636), .A2(new_n715), .A3(new_n750), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n739), .A3(new_n722), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  AND2_X1   g570(.A1(new_n323), .A2(new_n403), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n695), .A2(new_n513), .A3(new_n696), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n504), .A2(KEYINPUT110), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n503), .A2(new_n761), .A3(new_n481), .A4(new_n488), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n760), .A2(G469), .A3(new_n501), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n499), .B(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n498), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n511), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n758), .B1(new_n759), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n764), .ZN(new_n768));
  AOI21_X1  g582(.A(G902), .B1(new_n487), .B2(new_n495), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n768), .B1(new_n769), .B2(new_n497), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n510), .B1(new_n770), .B2(new_n763), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n470), .A2(new_n771), .A3(KEYINPUT111), .A4(new_n513), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n757), .A2(KEYINPUT42), .A3(new_n722), .A4(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n323), .A3(new_n403), .A4(new_n722), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G131), .ZN(G33));
  NAND4_X1  g593(.A1(new_n773), .A2(new_n323), .A3(new_n403), .A4(new_n692), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G134), .ZN(G36));
  AND2_X1   g595(.A1(new_n657), .A2(new_n659), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(KEYINPUT43), .A3(new_n575), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n575), .B(KEYINPUT114), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n660), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n783), .B1(new_n785), .B2(KEYINPUT43), .ZN(new_n786));
  INV_X1    g600(.A(new_n638), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n787), .A3(new_n683), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n759), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n787), .A4(new_n683), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT115), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT45), .B1(new_n501), .B2(new_n504), .ZN(new_n795));
  OR3_X1    g609(.A1(new_n795), .A2(KEYINPUT112), .A3(new_n497), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT112), .B1(new_n795), .B2(new_n497), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n760), .A2(KEYINPUT45), .A3(new_n501), .A4(new_n762), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n768), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT46), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n498), .B1(new_n802), .B2(KEYINPUT46), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n511), .B(new_n711), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n790), .A2(new_n807), .A3(new_n791), .A4(new_n792), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n794), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G137), .ZN(G39));
  OAI21_X1  g624(.A(new_n511), .B1(new_n803), .B2(new_n804), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(KEYINPUT47), .B(new_n511), .C1(new_n803), .C2(new_n804), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n722), .A2(new_n791), .A3(new_n402), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n323), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NOR3_X1   g633(.A1(new_n402), .A2(new_n514), .A3(new_n510), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT116), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n730), .B(KEYINPUT49), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n785), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n709), .A3(new_n718), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n746), .A2(new_n697), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n683), .A2(new_n766), .A3(new_n691), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n708), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n723), .A2(new_n828), .A3(new_n755), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n704), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n704), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n512), .A2(new_n622), .A3(new_n575), .A4(new_n691), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n323), .A2(new_n683), .A3(new_n791), .A4(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n773), .A2(new_n722), .A3(new_n754), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n780), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n777), .B2(new_n774), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n752), .A2(new_n734), .A3(new_n737), .A4(new_n740), .ZN(new_n838));
  INV_X1    g652(.A(new_n661), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n697), .A3(new_n840), .A4(new_n631), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT117), .B1(new_n640), .B2(new_n661), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n638), .A4(new_n639), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n633), .A2(new_n843), .A3(new_n671), .A4(new_n685), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n837), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n825), .B1(new_n832), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n704), .A2(new_n829), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n704), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n837), .A2(new_n845), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n844), .A2(new_n825), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n632), .A2(new_n683), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n742), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n860), .A2(new_n323), .B1(new_n748), .B2(new_n751), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n862), .A3(new_n734), .A4(new_n737), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n857), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n852), .A2(new_n864), .A3(new_n837), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n847), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n856), .B1(KEYINPUT54), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n733), .A2(new_n791), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT119), .Z(new_n869));
  AOI211_X1 g683(.A(new_n689), .B(new_n783), .C1(new_n785), .C2(KEYINPUT43), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n869), .A2(new_n754), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n708), .A2(new_n402), .A3(new_n627), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n782), .A2(new_n668), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n751), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n718), .A2(new_n514), .A3(new_n733), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n876), .A2(new_n759), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n730), .A2(new_n511), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n815), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT51), .ZN(new_n886));
  OAI221_X1 g700(.A(new_n625), .B1(new_n742), .B2(new_n876), .C1(new_n873), .C2(new_n661), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n869), .A2(new_n757), .A3(new_n870), .ZN(new_n888));
  XNOR2_X1  g702(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n888), .A2(new_n890), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n867), .A2(new_n885), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n824), .B1(new_n895), .B2(new_n896), .ZN(G75));
  NOR2_X1   g711(.A1(new_n384), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n866), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(G210), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n443), .A2(new_n451), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n449), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT55), .Z(new_n906));
  OAI21_X1  g720(.A(new_n899), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n906), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n903), .A2(KEYINPUT121), .A3(new_n906), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n800), .A2(new_n801), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT123), .Z(new_n914));
  NOR2_X1   g728(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n764), .B(KEYINPUT57), .Z(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n852), .B2(new_n853), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n837), .A2(new_n863), .A3(new_n858), .A4(new_n857), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n832), .A2(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n919), .A3(KEYINPUT54), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n847), .B2(new_n865), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n916), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n496), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n923), .A2(KEYINPUT122), .A3(new_n496), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n898), .B1(new_n926), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n567), .ZN(new_n929));
  NAND2_X1  g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n901), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n899), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n901), .A2(new_n929), .A3(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G60));
  NOR2_X1   g748(.A1(new_n654), .A2(new_n656), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n649), .B2(new_n650), .ZN(new_n936));
  NAND2_X1  g750(.A1(G478), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT59), .Z(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n867), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n936), .B(new_n939), .C1(new_n920), .C2(new_n922), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n899), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT124), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT60), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n946), .B1(new_n847), .B2(new_n865), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(new_n399), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n677), .A3(new_n675), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n899), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G66));
  INV_X1    g766(.A(new_n629), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n953), .B2(new_n446), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n845), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n904), .B1(G898), .B2(new_n384), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND3_X1  g771(.A1(new_n806), .A2(new_n757), .A3(new_n826), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n818), .A2(new_n778), .A3(new_n780), .A4(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n704), .A2(new_n723), .A3(new_n755), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n809), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n809), .A2(KEYINPUT126), .A3(new_n960), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n384), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT125), .Z(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(new_n561), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n384), .B1(G227), .B2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n661), .A2(new_n669), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n712), .A2(new_n759), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n757), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n809), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n960), .A2(new_n720), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n815), .A2(new_n817), .B1(new_n979), .B2(KEYINPUT62), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n982), .A2(new_n384), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n972), .B(new_n974), .C1(new_n983), .C2(new_n969), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n969), .ZN(new_n985));
  INV_X1    g799(.A(new_n971), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n965), .B2(new_n384), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n973), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n984), .A2(new_n988), .ZN(G72));
  XNOR2_X1  g803(.A(new_n292), .B(KEYINPUT127), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n263), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n965), .A2(new_n845), .ZN(new_n992));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n978), .A2(new_n981), .A3(new_n845), .A4(new_n980), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n263), .B(new_n990), .C1(new_n996), .C2(new_n994), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n293), .A2(new_n312), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n855), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n995), .A2(new_n997), .A3(new_n898), .A4(new_n999), .ZN(G57));
endmodule


