

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781;

  OR2_X1 U378 ( .A1(n738), .A2(n419), .ZN(n418) );
  XNOR2_X2 U379 ( .A(n390), .B(n389), .ZN(n388) );
  XNOR2_X2 U380 ( .A(n770), .B(n440), .ZN(n489) );
  XNOR2_X2 U381 ( .A(n506), .B(n439), .ZN(n770) );
  XNOR2_X2 U382 ( .A(n595), .B(KEYINPUT35), .ZN(n779) );
  AND2_X1 U383 ( .A1(n675), .A2(n576), .ZN(n559) );
  INV_X1 U384 ( .A(KEYINPUT48), .ZN(n389) );
  INV_X4 U385 ( .A(G953), .ZN(n771) );
  AND2_X1 U386 ( .A1(n414), .A2(n423), .ZN(n413) );
  NAND2_X1 U387 ( .A1(n399), .A2(n617), .ZN(n398) );
  XNOR2_X1 U388 ( .A(n416), .B(KEYINPUT32), .ZN(n647) );
  XNOR2_X1 U389 ( .A(n559), .B(n558), .ZN(n778) );
  XNOR2_X1 U390 ( .A(n394), .B(n393), .ZN(n671) );
  XNOR2_X1 U391 ( .A(n606), .B(n405), .ZN(n604) );
  XNOR2_X1 U392 ( .A(n466), .B(n387), .ZN(n702) );
  AND2_X2 U393 ( .A1(n418), .A2(n358), .ZN(n417) );
  XNOR2_X1 U394 ( .A(n537), .B(KEYINPUT4), .ZN(n506) );
  XNOR2_X1 U395 ( .A(KEYINPUT70), .B(KEYINPUT3), .ZN(n441) );
  NAND2_X2 U396 ( .A1(n413), .A2(n411), .ZN(n642) );
  NAND2_X1 U397 ( .A1(n370), .A2(n623), .ZN(n380) );
  NOR2_X1 U398 ( .A1(n604), .A2(n359), .ZN(n370) );
  NAND2_X1 U399 ( .A1(n604), .A2(n359), .ZN(n382) );
  XNOR2_X1 U400 ( .A(n438), .B(G125), .ZN(n500) );
  XNOR2_X1 U401 ( .A(n408), .B(G140), .ZN(n484) );
  INV_X1 U402 ( .A(G137), .ZN(n408) );
  INV_X1 U403 ( .A(n381), .ZN(n374) );
  AND2_X1 U404 ( .A1(n380), .A2(n373), .ZN(n372) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n443) );
  NOR2_X1 U406 ( .A1(n675), .A2(n671), .ZN(n566) );
  NAND2_X1 U407 ( .A1(n400), .A2(n620), .ZN(n399) );
  XNOR2_X1 U408 ( .A(KEYINPUT10), .B(KEYINPUT69), .ZN(n452) );
  XNOR2_X1 U409 ( .A(G122), .B(G113), .ZN(n516) );
  XNOR2_X1 U410 ( .A(n525), .B(n518), .ZN(n397) );
  INV_X1 U411 ( .A(KEYINPUT12), .ZN(n518) );
  INV_X1 U412 ( .A(n723), .ZN(n433) );
  NAND2_X1 U413 ( .A1(n634), .A2(n420), .ZN(n419) );
  INV_X1 U414 ( .A(n509), .ZN(n420) );
  XNOR2_X1 U415 ( .A(n464), .B(KEYINPUT77), .ZN(n465) );
  NAND2_X1 U416 ( .A1(n367), .A2(n364), .ZN(n552) );
  AND2_X1 U417 ( .A1(n369), .A2(n368), .ZN(n367) );
  NAND2_X1 U418 ( .A1(n491), .A2(n366), .ZN(n365) );
  NOR2_X1 U419 ( .A1(n703), .A2(n702), .ZN(n706) );
  INV_X1 U420 ( .A(G122), .ZN(n495) );
  XNOR2_X1 U421 ( .A(n363), .B(G143), .ZN(n537) );
  XNOR2_X1 U422 ( .A(G128), .B(KEYINPUT81), .ZN(n363) );
  INV_X1 U423 ( .A(G107), .ZN(n533) );
  INV_X1 U424 ( .A(KEYINPUT64), .ZN(n641) );
  XNOR2_X1 U425 ( .A(n485), .B(n410), .ZN(n409) );
  INV_X1 U426 ( .A(KEYINPUT78), .ZN(n410) );
  AND2_X1 U427 ( .A1(n378), .A2(n376), .ZN(n375) );
  INV_X1 U428 ( .A(n553), .ZN(n606) );
  XNOR2_X1 U429 ( .A(n541), .B(n540), .ZN(n564) );
  XNOR2_X1 U430 ( .A(n528), .B(n527), .ZN(n565) );
  XNOR2_X1 U431 ( .A(n526), .B(n648), .ZN(n527) );
  NAND2_X1 U432 ( .A1(n589), .A2(n588), .ZN(n591) );
  INV_X1 U433 ( .A(n606), .ZN(n406) );
  XNOR2_X1 U434 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U435 ( .A(KEYINPUT92), .B(n646), .Z(n756) );
  NAND2_X1 U436 ( .A1(n647), .A2(n610), .ZN(n415) );
  NAND2_X1 U437 ( .A1(G469), .A2(G902), .ZN(n368) );
  NAND2_X1 U438 ( .A1(n392), .A2(n391), .ZN(n390) );
  AND2_X1 U439 ( .A1(n575), .A2(n356), .ZN(n391) );
  INV_X1 U440 ( .A(n415), .ZN(n617) );
  AND2_X1 U441 ( .A1(n638), .A2(n427), .ZN(n424) );
  NAND2_X1 U442 ( .A1(n691), .A2(n425), .ZN(n423) );
  NOR2_X1 U443 ( .A1(n636), .A2(n640), .ZN(n425) );
  XNOR2_X1 U444 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n502) );
  NAND2_X1 U445 ( .A1(G237), .A2(G234), .ZN(n468) );
  NOR2_X1 U446 ( .A1(n709), .A2(n406), .ZN(n710) );
  INV_X1 U447 ( .A(G237), .ZN(n508) );
  NAND2_X1 U448 ( .A1(n380), .A2(n627), .ZN(n377) );
  NAND2_X1 U449 ( .A1(n639), .A2(n509), .ZN(n421) );
  XNOR2_X1 U450 ( .A(n552), .B(KEYINPUT1), .ZN(n583) );
  INV_X1 U451 ( .A(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U452 ( .A(n489), .B(n449), .ZN(n657) );
  XNOR2_X1 U453 ( .A(n453), .B(n484), .ZN(n769) );
  XNOR2_X1 U454 ( .A(G128), .B(G119), .ZN(n454) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n650) );
  XNOR2_X1 U456 ( .A(n521), .B(n519), .ZN(n395) );
  XNOR2_X1 U457 ( .A(n523), .B(n397), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n432), .B(n431), .ZN(n717) );
  XNOR2_X1 U459 ( .A(n549), .B(KEYINPUT112), .ZN(n431) );
  NAND2_X1 U460 ( .A1(n623), .A2(n406), .ZN(n713) );
  XNOR2_X1 U461 ( .A(n554), .B(n386), .ZN(n385) );
  INV_X1 U462 ( .A(KEYINPUT30), .ZN(n386) );
  AND2_X1 U463 ( .A1(n542), .A2(n406), .ZN(n483) );
  XNOR2_X1 U464 ( .A(n465), .B(n467), .ZN(n387) );
  BUF_X1 U465 ( .A(n583), .Z(n705) );
  XNOR2_X1 U466 ( .A(n498), .B(n497), .ZN(n764) );
  XOR2_X1 U467 ( .A(KEYINPUT16), .B(KEYINPUT73), .Z(n496) );
  XNOR2_X1 U468 ( .A(n539), .B(n538), .ZN(n754) );
  XNOR2_X1 U469 ( .A(n536), .B(n535), .ZN(n539) );
  XNOR2_X1 U470 ( .A(n489), .B(n490), .ZN(n747) );
  XNOR2_X1 U471 ( .A(n409), .B(n484), .ZN(n487) );
  NAND2_X1 U472 ( .A1(n375), .A2(n371), .ZN(n594) );
  INV_X1 U473 ( .A(KEYINPUT104), .ZN(n393) );
  NAND2_X1 U474 ( .A1(n565), .A2(n564), .ZN(n394) );
  NOR2_X1 U475 ( .A1(n626), .A2(n406), .ZN(n628) );
  INV_X1 U476 ( .A(KEYINPUT126), .ZN(n428) );
  INV_X1 U477 ( .A(G902), .ZN(n366) );
  OR2_X1 U478 ( .A1(n381), .A2(n379), .ZN(n699) );
  INV_X1 U479 ( .A(G146), .ZN(n438) );
  AND2_X1 U480 ( .A1(n547), .A2(n686), .ZN(n356) );
  INV_X1 U481 ( .A(n691), .ZN(n638) );
  AND2_X1 U482 ( .A1(n418), .A2(n421), .ZN(n357) );
  AND2_X1 U483 ( .A1(n421), .A2(n719), .ZN(n358) );
  XOR2_X1 U484 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n359) );
  AND2_X1 U485 ( .A1(n426), .A2(n427), .ZN(n360) );
  INV_X1 U486 ( .A(KEYINPUT34), .ZN(n384) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(KEYINPUT45), .Z(n361) );
  NAND2_X1 U488 ( .A1(n639), .A2(n637), .ZN(n362) );
  NAND2_X1 U489 ( .A1(n747), .A2(G469), .ZN(n369) );
  OR2_X1 U490 ( .A1(n747), .A2(n365), .ZN(n364) );
  NAND2_X1 U491 ( .A1(n374), .A2(n372), .ZN(n371) );
  AND2_X1 U492 ( .A1(n627), .A2(KEYINPUT34), .ZN(n373) );
  NAND2_X1 U493 ( .A1(n377), .A2(n384), .ZN(n376) );
  NAND2_X1 U494 ( .A1(n381), .A2(n384), .ZN(n378) );
  INV_X1 U495 ( .A(n380), .ZN(n379) );
  NAND2_X1 U496 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U497 ( .A1(n622), .A2(n359), .ZN(n383) );
  NOR2_X1 U498 ( .A1(n695), .A2(n362), .ZN(n412) );
  NOR2_X1 U499 ( .A1(n691), .A2(n695), .ZN(n690) );
  OR2_X1 U500 ( .A1(n695), .A2(G953), .ZN(n759) );
  XNOR2_X2 U501 ( .A(n407), .B(n361), .ZN(n695) );
  NAND2_X1 U502 ( .A1(n583), .A2(n706), .ZN(n622) );
  NAND2_X1 U503 ( .A1(n412), .A2(n424), .ZN(n411) );
  NAND2_X2 U504 ( .A1(n388), .A2(n582), .ZN(n691) );
  AND2_X2 U505 ( .A1(n608), .A2(n604), .ZN(n611) );
  AND2_X2 U506 ( .A1(n781), .A2(n632), .ZN(n402) );
  XNOR2_X2 U507 ( .A(n544), .B(n512), .ZN(n589) );
  NAND2_X2 U508 ( .A1(n417), .A2(n422), .ZN(n544) );
  OR2_X2 U509 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U510 ( .A1(n385), .A2(n555), .ZN(n556) );
  NAND2_X1 U511 ( .A1(n600), .A2(n433), .ZN(n432) );
  NAND2_X1 U512 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U513 ( .A1(n779), .A2(n596), .ZN(n618) );
  XNOR2_X1 U514 ( .A(n560), .B(KEYINPUT46), .ZN(n392) );
  NAND2_X1 U515 ( .A1(n401), .A2(n398), .ZN(n407) );
  NAND2_X1 U516 ( .A1(n597), .A2(n596), .ZN(n400) );
  AND2_X2 U517 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X2 U518 ( .A(n616), .B(KEYINPUT106), .ZN(n781) );
  NAND2_X1 U519 ( .A1(n404), .A2(n621), .ZN(n403) );
  NAND2_X1 U520 ( .A1(n618), .A2(n619), .ZN(n404) );
  XNOR2_X1 U521 ( .A(n488), .B(KEYINPUT79), .ZN(n490) );
  NAND2_X1 U522 ( .A1(n695), .A2(n360), .ZN(n414) );
  NAND2_X1 U523 ( .A1(n415), .A2(n620), .ZN(n619) );
  NAND2_X1 U524 ( .A1(n611), .A2(n605), .ZN(n416) );
  NAND2_X1 U525 ( .A1(n422), .A2(n357), .ZN(n581) );
  NAND2_X1 U526 ( .A1(n738), .A2(n509), .ZN(n422) );
  INV_X1 U527 ( .A(n636), .ZN(n426) );
  INV_X1 U528 ( .A(n640), .ZN(n427) );
  XNOR2_X1 U529 ( .A(n429), .B(n428), .ZN(G66) );
  NAND2_X1 U530 ( .A1(n430), .A2(n756), .ZN(n429) );
  XNOR2_X1 U531 ( .A(n645), .B(n644), .ZN(n430) );
  XNOR2_X1 U532 ( .A(n500), .B(n452), .ZN(n522) );
  NOR2_X1 U533 ( .A1(n656), .A2(n643), .ZN(n645) );
  XNOR2_X1 U534 ( .A(n494), .B(n493), .ZN(n498) );
  XOR2_X1 U535 ( .A(n447), .B(n446), .Z(n434) );
  XOR2_X1 U536 ( .A(n580), .B(KEYINPUT43), .Z(n435) );
  AND2_X1 U537 ( .A1(n676), .A2(n573), .ZN(n436) );
  INV_X1 U538 ( .A(n555), .ZN(n481) );
  INV_X1 U539 ( .A(n494), .ZN(n445) );
  NOR2_X1 U540 ( .A1(n481), .A2(n703), .ZN(n482) );
  AND2_X1 U541 ( .A1(n702), .A2(n482), .ZN(n542) );
  XNOR2_X1 U542 ( .A(n448), .B(n434), .ZN(n449) );
  XNOR2_X1 U543 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U544 ( .A(KEYINPUT47), .B(KEYINPUT84), .ZN(n515) );
  INV_X1 U545 ( .A(KEYINPUT67), .ZN(n437) );
  XNOR2_X1 U546 ( .A(n437), .B(G101), .ZN(n499) );
  XNOR2_X1 U547 ( .A(n499), .B(G146), .ZN(n440) );
  XOR2_X1 U548 ( .A(G134), .B(G131), .Z(n439) );
  XOR2_X2 U549 ( .A(G113), .B(G119), .Z(n442) );
  XNOR2_X2 U550 ( .A(n442), .B(n441), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT75), .B(n443), .Z(n520) );
  NAND2_X1 U552 ( .A1(n520), .A2(G210), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n445), .B(n444), .ZN(n448) );
  XOR2_X1 U554 ( .A(G137), .B(KEYINPUT98), .Z(n447) );
  XNOR2_X1 U555 ( .A(G116), .B(KEYINPUT5), .ZN(n446) );
  NOR2_X1 U556 ( .A1(G902), .A2(n657), .ZN(n451) );
  XNOR2_X1 U557 ( .A(KEYINPUT99), .B(G472), .ZN(n450) );
  XNOR2_X1 U558 ( .A(n451), .B(n450), .ZN(n553) );
  INV_X1 U559 ( .A(n522), .ZN(n453) );
  XNOR2_X1 U560 ( .A(n769), .B(KEYINPUT23), .ZN(n461) );
  XOR2_X1 U561 ( .A(KEYINPUT71), .B(G110), .Z(n455) );
  XNOR2_X1 U562 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U563 ( .A(n456), .B(KEYINPUT24), .Z(n459) );
  NAND2_X1 U564 ( .A1(G234), .A2(n771), .ZN(n457) );
  XOR2_X1 U565 ( .A(KEYINPUT8), .B(n457), .Z(n529) );
  AND2_X1 U566 ( .A1(n529), .A2(G221), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n644) );
  NOR2_X1 U568 ( .A1(n644), .A2(G902), .ZN(n466) );
  XNOR2_X1 U569 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n462) );
  XNOR2_X1 U570 ( .A(n462), .B(n366), .ZN(n634) );
  NAND2_X1 U571 ( .A1(n634), .A2(G234), .ZN(n463) );
  XNOR2_X1 U572 ( .A(n463), .B(KEYINPUT20), .ZN(n478) );
  NAND2_X1 U573 ( .A1(G217), .A2(n478), .ZN(n464) );
  XOR2_X1 U574 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n467) );
  XNOR2_X1 U575 ( .A(n468), .B(KEYINPUT14), .ZN(n472) );
  NAND2_X1 U576 ( .A1(G902), .A2(n472), .ZN(n585) );
  OR2_X1 U577 ( .A1(n771), .A2(n585), .ZN(n469) );
  XNOR2_X1 U578 ( .A(KEYINPUT108), .B(n469), .ZN(n470) );
  NOR2_X1 U579 ( .A1(G900), .A2(n470), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n471), .B(KEYINPUT109), .ZN(n477) );
  NAND2_X1 U581 ( .A1(n472), .A2(G952), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n473), .B(KEYINPUT94), .ZN(n732) );
  NOR2_X1 U583 ( .A1(G953), .A2(n732), .ZN(n475) );
  INV_X1 U584 ( .A(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U585 ( .A(n475), .B(n474), .ZN(n586) );
  INV_X1 U586 ( .A(n586), .ZN(n476) );
  NAND2_X1 U587 ( .A1(n477), .A2(n476), .ZN(n555) );
  AND2_X1 U588 ( .A1(n478), .A2(G221), .ZN(n480) );
  INV_X1 U589 ( .A(KEYINPUT21), .ZN(n479) );
  XNOR2_X1 U590 ( .A(n480), .B(n479), .ZN(n703) );
  XNOR2_X1 U591 ( .A(n483), .B(KEYINPUT28), .ZN(n492) );
  NAND2_X1 U592 ( .A1(n771), .A2(G227), .ZN(n485) );
  XNOR2_X1 U593 ( .A(G107), .B(G104), .ZN(n486) );
  XNOR2_X1 U594 ( .A(n486), .B(G110), .ZN(n493) );
  XNOR2_X1 U595 ( .A(n487), .B(n493), .ZN(n488) );
  INV_X1 U596 ( .A(G469), .ZN(n491) );
  NAND2_X1 U597 ( .A1(n492), .A2(n552), .ZN(n550) );
  XNOR2_X1 U598 ( .A(n495), .B(G116), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n496), .B(n532), .ZN(n497) );
  XNOR2_X1 U600 ( .A(n500), .B(n499), .ZN(n504) );
  NAND2_X1 U601 ( .A1(n771), .A2(G224), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U603 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U604 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U605 ( .A(n764), .B(n507), .ZN(n738) );
  INV_X1 U606 ( .A(n634), .ZN(n639) );
  NAND2_X1 U607 ( .A1(n366), .A2(n508), .ZN(n510) );
  NAND2_X1 U608 ( .A1(n510), .A2(G210), .ZN(n509) );
  NAND2_X1 U609 ( .A1(n510), .A2(G214), .ZN(n719) );
  XNOR2_X1 U610 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n511), .B(KEYINPUT66), .ZN(n512) );
  INV_X1 U612 ( .A(n589), .ZN(n513) );
  NOR2_X1 U613 ( .A1(n550), .A2(n513), .ZN(n676) );
  INV_X1 U614 ( .A(n676), .ZN(n514) );
  NAND2_X1 U615 ( .A1(n515), .A2(n514), .ZN(n547) );
  XOR2_X1 U616 ( .A(KEYINPUT101), .B(G104), .Z(n517) );
  XNOR2_X1 U617 ( .A(n517), .B(n516), .ZN(n519) );
  NAND2_X1 U618 ( .A1(G214), .A2(n520), .ZN(n521) );
  XNOR2_X1 U619 ( .A(n522), .B(G140), .ZN(n523) );
  XNOR2_X1 U620 ( .A(G143), .B(G131), .ZN(n524) );
  XNOR2_X1 U621 ( .A(n524), .B(KEYINPUT11), .ZN(n525) );
  NOR2_X1 U622 ( .A1(G902), .A2(n650), .ZN(n528) );
  XNOR2_X1 U623 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n526) );
  INV_X1 U624 ( .A(G475), .ZN(n648) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n531) );
  NAND2_X1 U626 ( .A1(G217), .A2(n529), .ZN(n530) );
  XNOR2_X1 U627 ( .A(n531), .B(n530), .ZN(n536) );
  XNOR2_X1 U628 ( .A(G134), .B(n532), .ZN(n534) );
  INV_X1 U629 ( .A(n537), .ZN(n538) );
  NAND2_X1 U630 ( .A1(n754), .A2(n366), .ZN(n541) );
  XOR2_X1 U631 ( .A(G478), .B(KEYINPUT103), .Z(n540) );
  OR2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n678) );
  INV_X1 U633 ( .A(n678), .ZN(n675) );
  NAND2_X1 U634 ( .A1(n542), .A2(n675), .ZN(n543) );
  OR2_X1 U635 ( .A1(n543), .A2(n604), .ZN(n577) );
  NOR2_X1 U636 ( .A1(n577), .A2(n544), .ZN(n545) );
  XNOR2_X1 U637 ( .A(n545), .B(KEYINPUT36), .ZN(n546) );
  NAND2_X1 U638 ( .A1(n546), .A2(n705), .ZN(n686) );
  INV_X1 U639 ( .A(n564), .ZN(n548) );
  AND2_X1 U640 ( .A1(n565), .A2(n548), .ZN(n600) );
  INV_X1 U641 ( .A(n600), .ZN(n722) );
  XNOR2_X1 U642 ( .A(n581), .B(KEYINPUT38), .ZN(n720) );
  XNOR2_X1 U643 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n549) );
  NOR2_X1 U644 ( .A1(n550), .A2(n717), .ZN(n551) );
  XNOR2_X1 U645 ( .A(n551), .B(KEYINPUT42), .ZN(n780) );
  NAND2_X1 U646 ( .A1(n552), .A2(n706), .ZN(n626) );
  NAND2_X1 U647 ( .A1(n553), .A2(n719), .ZN(n554) );
  NOR2_X2 U648 ( .A1(n626), .A2(n556), .ZN(n563) );
  NAND2_X1 U649 ( .A1(n563), .A2(n720), .ZN(n557) );
  XNOR2_X1 U650 ( .A(n557), .B(KEYINPUT39), .ZN(n576) );
  XNOR2_X1 U651 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n558) );
  NOR2_X1 U652 ( .A1(n780), .A2(n778), .ZN(n560) );
  INV_X1 U653 ( .A(n565), .ZN(n561) );
  NAND2_X1 U654 ( .A1(n561), .A2(n564), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n592), .A2(n581), .ZN(n562) );
  AND2_X1 U656 ( .A1(n563), .A2(n562), .ZN(n674) );
  XNOR2_X1 U657 ( .A(n674), .B(KEYINPUT85), .ZN(n568) );
  XNOR2_X1 U658 ( .A(n566), .B(KEYINPUT105), .ZN(n630) );
  INV_X1 U659 ( .A(n630), .ZN(n724) );
  NAND2_X1 U660 ( .A1(KEYINPUT47), .A2(n724), .ZN(n567) );
  NAND2_X1 U661 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U662 ( .A(KEYINPUT82), .B(n569), .ZN(n574) );
  XOR2_X1 U663 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n570) );
  NAND2_X1 U664 ( .A1(n570), .A2(n630), .ZN(n571) );
  XNOR2_X1 U665 ( .A(KEYINPUT74), .B(n571), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n572), .A2(KEYINPUT84), .ZN(n573) );
  NOR2_X1 U667 ( .A1(n574), .A2(n436), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n576), .A2(n671), .ZN(n687) );
  INV_X1 U669 ( .A(n577), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n578), .A2(n719), .ZN(n579) );
  NOR2_X1 U671 ( .A1(n705), .A2(n579), .ZN(n580) );
  NAND2_X1 U672 ( .A1(n435), .A2(n581), .ZN(n688) );
  AND2_X1 U673 ( .A1(n687), .A2(n688), .ZN(n582) );
  NOR2_X1 U674 ( .A1(G898), .A2(n771), .ZN(n584) );
  XOR2_X1 U675 ( .A(KEYINPUT96), .B(n584), .Z(n765) );
  NOR2_X1 U676 ( .A1(n765), .A2(n585), .ZN(n587) );
  OR2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U678 ( .A(KEYINPUT0), .ZN(n590) );
  XNOR2_X2 U679 ( .A(n591), .B(n590), .ZN(n627) );
  INV_X1 U680 ( .A(n627), .ZN(n624) );
  XOR2_X1 U681 ( .A(n592), .B(KEYINPUT80), .Z(n593) );
  NAND2_X1 U682 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U683 ( .A(n779), .ZN(n597) );
  INV_X1 U684 ( .A(KEYINPUT44), .ZN(n596) );
  INV_X1 U685 ( .A(KEYINPUT65), .ZN(n620) );
  NAND2_X1 U686 ( .A1(n705), .A2(n702), .ZN(n598) );
  XNOR2_X1 U687 ( .A(n598), .B(KEYINPUT107), .ZN(n605) );
  INV_X1 U688 ( .A(n703), .ZN(n599) );
  AND2_X1 U689 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U690 ( .A1(n627), .A2(n601), .ZN(n603) );
  INV_X1 U691 ( .A(KEYINPUT22), .ZN(n602) );
  XNOR2_X1 U692 ( .A(n603), .B(n602), .ZN(n608) );
  NAND2_X1 U693 ( .A1(n702), .A2(n606), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n705), .A2(n607), .ZN(n609) );
  AND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n670) );
  INV_X1 U696 ( .A(n670), .ZN(n610) );
  XNOR2_X1 U697 ( .A(n611), .B(KEYINPUT89), .ZN(n615) );
  INV_X1 U698 ( .A(n702), .ZN(n613) );
  INV_X1 U699 ( .A(n705), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n620), .A2(n596), .ZN(n621) );
  INV_X1 U702 ( .A(n622), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n713), .A2(n624), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT31), .ZN(n682) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n667) );
  NAND2_X1 U706 ( .A1(n682), .A2(n667), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n629), .B(KEYINPUT100), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n632) );
  INV_X1 U709 ( .A(KEYINPUT87), .ZN(n633) );
  OR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n635), .A2(KEYINPUT2), .ZN(n636) );
  INV_X1 U712 ( .A(KEYINPUT2), .ZN(n637) );
  NOR2_X1 U713 ( .A1(n639), .A2(KEYINPUT87), .ZN(n640) );
  XNOR2_X2 U714 ( .A(n642), .B(n641), .ZN(n656) );
  INV_X1 U715 ( .A(G217), .ZN(n643) );
  NOR2_X1 U716 ( .A1(n771), .A2(G952), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(G119), .ZN(G21) );
  INV_X1 U718 ( .A(KEYINPUT60), .ZN(n655) );
  NOR2_X1 U719 ( .A1(n656), .A2(n648), .ZN(n652) );
  XOR2_X1 U720 ( .A(KEYINPUT90), .B(KEYINPUT59), .Z(n649) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n653), .A2(n756), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G60) );
  INV_X1 U725 ( .A(n656), .ZN(n753) );
  NAND2_X1 U726 ( .A1(n753), .A2(G472), .ZN(n659) );
  XOR2_X1 U727 ( .A(n657), .B(KEYINPUT62), .Z(n658) );
  XNOR2_X1 U728 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n660), .A2(n756), .ZN(n663) );
  XNOR2_X1 U730 ( .A(KEYINPUT63), .B(KEYINPUT113), .ZN(n661) );
  XNOR2_X1 U731 ( .A(n661), .B(KEYINPUT91), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n663), .B(n662), .ZN(G57) );
  NOR2_X1 U733 ( .A1(n667), .A2(n678), .ZN(n664) );
  XOR2_X1 U734 ( .A(G104), .B(n664), .Z(G6) );
  XOR2_X1 U735 ( .A(KEYINPUT26), .B(KEYINPUT114), .Z(n666) );
  XNOR2_X1 U736 ( .A(G107), .B(KEYINPUT27), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n669) );
  INV_X1 U738 ( .A(n671), .ZN(n683) );
  NOR2_X1 U739 ( .A1(n667), .A2(n683), .ZN(n668) );
  XOR2_X1 U740 ( .A(n669), .B(n668), .Z(G9) );
  XOR2_X1 U741 ( .A(G110), .B(n670), .Z(G12) );
  XOR2_X1 U742 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U743 ( .A1(n676), .A2(n671), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n673), .B(n672), .ZN(G30) );
  XOR2_X1 U745 ( .A(G143), .B(n674), .Z(G45) );
  NAND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(G146), .ZN(G48) );
  NOR2_X1 U748 ( .A1(n678), .A2(n682), .ZN(n680) );
  XNOR2_X1 U749 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U751 ( .A(G113), .B(n681), .ZN(G15) );
  NOR2_X1 U752 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U753 ( .A(G116), .B(n684), .Z(G18) );
  XOR2_X1 U754 ( .A(G125), .B(KEYINPUT37), .Z(n685) );
  XNOR2_X1 U755 ( .A(n686), .B(n685), .ZN(G27) );
  XNOR2_X1 U756 ( .A(G134), .B(n687), .ZN(G36) );
  XOR2_X1 U757 ( .A(G140), .B(n688), .Z(n689) );
  XNOR2_X1 U758 ( .A(n689), .B(KEYINPUT117), .ZN(G42) );
  NAND2_X1 U759 ( .A1(n690), .A2(KEYINPUT2), .ZN(n693) );
  XNOR2_X1 U760 ( .A(KEYINPUT2), .B(KEYINPUT83), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n691), .A2(n694), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U764 ( .A(KEYINPUT86), .B(n696), .Z(n697) );
  NOR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U766 ( .A1(n717), .A2(n699), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n735) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U769 ( .A(KEYINPUT49), .B(n704), .Z(n711) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n708) );
  XNOR2_X1 U771 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U775 ( .A(n714), .B(KEYINPUT119), .Z(n715) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n715), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(KEYINPUT120), .ZN(n729) );
  NOR2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n699), .A2(n727), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U785 ( .A(n730), .B(KEYINPUT52), .ZN(n731) );
  NOR2_X1 U786 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U787 ( .A1(G953), .A2(n733), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT121), .B(n736), .ZN(n737) );
  XNOR2_X1 U790 ( .A(KEYINPUT53), .B(n737), .ZN(G75) );
  NAND2_X1 U791 ( .A1(n753), .A2(G210), .ZN(n741) );
  XOR2_X1 U792 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n739) );
  XOR2_X1 U793 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U794 ( .A(n741), .B(n740), .ZN(n742) );
  NAND2_X1 U795 ( .A1(n742), .A2(n756), .ZN(n744) );
  XOR2_X1 U796 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n743) );
  XNOR2_X1 U797 ( .A(n744), .B(n743), .ZN(G51) );
  INV_X1 U798 ( .A(n756), .ZN(n752) );
  XOR2_X1 U799 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n746) );
  XNOR2_X1 U800 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n745) );
  XNOR2_X1 U801 ( .A(n746), .B(n745), .ZN(n748) );
  XNOR2_X1 U802 ( .A(n748), .B(n747), .ZN(n750) );
  NAND2_X1 U803 ( .A1(n753), .A2(G469), .ZN(n749) );
  XOR2_X1 U804 ( .A(n750), .B(n749), .Z(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(G54) );
  NAND2_X1 U806 ( .A1(n753), .A2(G478), .ZN(n755) );
  XNOR2_X1 U807 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U809 ( .A(n758), .B(KEYINPUT125), .ZN(G63) );
  XOR2_X1 U810 ( .A(KEYINPUT127), .B(n759), .Z(n763) );
  NAND2_X1 U811 ( .A1(G953), .A2(G224), .ZN(n760) );
  XNOR2_X1 U812 ( .A(KEYINPUT61), .B(n760), .ZN(n761) );
  NAND2_X1 U813 ( .A1(n761), .A2(G898), .ZN(n762) );
  NAND2_X1 U814 ( .A1(n763), .A2(n762), .ZN(n768) );
  XOR2_X1 U815 ( .A(n764), .B(G101), .Z(n766) );
  NAND2_X1 U816 ( .A1(n766), .A2(n765), .ZN(n767) );
  XOR2_X1 U817 ( .A(n768), .B(n767), .Z(G69) );
  XOR2_X1 U818 ( .A(n770), .B(n769), .Z(n773) );
  XNOR2_X1 U819 ( .A(n691), .B(n773), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n772), .A2(n771), .ZN(n777) );
  XNOR2_X1 U821 ( .A(G227), .B(n773), .ZN(n774) );
  NAND2_X1 U822 ( .A1(n774), .A2(G900), .ZN(n775) );
  NAND2_X1 U823 ( .A1(n775), .A2(G953), .ZN(n776) );
  NAND2_X1 U824 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U825 ( .A(n778), .B(G131), .Z(G33) );
  XOR2_X1 U826 ( .A(n779), .B(G122), .Z(G24) );
  XOR2_X1 U827 ( .A(n780), .B(G137), .Z(G39) );
  XNOR2_X1 U828 ( .A(G101), .B(n781), .ZN(G3) );
endmodule

