//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G140), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n187), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(KEYINPUT78), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n193), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G953), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G953), .ZN(new_n204));
  INV_X1    g018(.A(G237), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n202), .A2(new_n204), .A3(G214), .A4(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(G953), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n209), .A2(G143), .A3(G214), .A4(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT18), .A2(G131), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n200), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n211), .B1(new_n208), .B2(new_n210), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT90), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n217), .A3(new_n200), .A4(new_n212), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G113), .B(G122), .ZN(new_n220));
  INV_X1    g034(.A(G104), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n189), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n198), .B2(new_n223), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n193), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n224), .B(G146), .C1(new_n198), .C2(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n210), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT17), .A3(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(G131), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n208), .A2(new_n210), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n229), .B(new_n231), .C1(new_n235), .C2(KEYINPUT17), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n219), .A2(new_n222), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT19), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n192), .A2(new_n238), .A3(new_n196), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n198), .A2(KEYINPUT19), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n193), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n241), .A2(new_n227), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n215), .A2(new_n218), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n237), .B1(new_n222), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G475), .A2(G902), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT91), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n247));
  INV_X1    g061(.A(G902), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n219), .A2(new_n222), .A3(new_n236), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n222), .B1(new_n219), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n246), .A2(new_n247), .B1(G475), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n242), .A2(new_n235), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n222), .B1(new_n219), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n245), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n244), .A2(KEYINPUT91), .A3(new_n245), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(KEYINPUT20), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G478), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(KEYINPUT15), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n207), .A2(G128), .ZN(new_n262));
  INV_X1    g076(.A(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n265), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G116), .B(G122), .ZN(new_n268));
  INV_X1    g082(.A(G107), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G116), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT14), .A3(G122), .ZN(new_n272));
  INV_X1    g086(.A(new_n268), .ZN(new_n273));
  OAI211_X1 g087(.A(G107), .B(new_n272), .C1(new_n273), .C2(KEYINPUT14), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n267), .A2(new_n270), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n262), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n264), .B1(new_n276), .B2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n262), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G134), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n268), .B(new_n269), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n265), .A2(new_n266), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT9), .B(G234), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(G953), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n275), .B2(new_n283), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n248), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n275), .A2(new_n283), .ZN(new_n292));
  INV_X1    g106(.A(new_n286), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT92), .A3(new_n248), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n261), .B1(new_n291), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n261), .ZN(new_n299));
  INV_X1    g113(.A(new_n289), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(KEYINPUT92), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT93), .B(G952), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(G234), .A2(G237), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n209), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n307), .A2(G902), .A3(new_n304), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT21), .B(G898), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n298), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n252), .A2(new_n259), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G469), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(new_n221), .B2(G107), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n269), .A3(G104), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n221), .A2(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G101), .ZN(new_n319));
  AOI21_X1  g133(.A(G101), .B1(new_n221), .B2(G107), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n314), .A2(new_n320), .A3(new_n316), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G143), .B(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT0), .A2(G128), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT64), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(KEYINPUT0), .B2(G128), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n193), .A2(G143), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n207), .A2(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT0), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT64), .B1(new_n332), .B2(new_n263), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n324), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n318), .A2(new_n336), .A3(G101), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n322), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n266), .B2(G137), .ZN(new_n340));
  INV_X1    g154(.A(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT11), .A3(G134), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n266), .A2(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G131), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n340), .A2(new_n342), .A3(new_n233), .A4(new_n343), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT1), .B1(new_n207), .B2(G146), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n207), .A2(G146), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n193), .A2(G143), .ZN(new_n351));
  OAI211_X1 g165(.A(G128), .B(new_n349), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n221), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n269), .A2(G104), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n329), .B(new_n330), .C1(KEYINPUT1), .C2(new_n263), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n352), .A2(new_n355), .A3(new_n321), .A4(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n357), .A2(KEYINPUT10), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(KEYINPUT10), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n338), .B(new_n348), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n357), .B(KEYINPUT10), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n363), .A2(KEYINPUT83), .A3(new_n348), .A4(new_n338), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n209), .A2(G227), .ZN(new_n366));
  XOR2_X1   g180(.A(G110), .B(G140), .Z(new_n367));
  XNOR2_X1  g181(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n357), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n356), .A2(new_n352), .B1(new_n355), .B2(new_n321), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n347), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT12), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n365), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n338), .B1(new_n358), .B2(new_n359), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT84), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n363), .A2(new_n378), .A3(new_n338), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n347), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n369), .B1(new_n365), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n313), .B(new_n248), .C1(new_n375), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(G469), .A2(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n365), .A2(new_n374), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n368), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n365), .A2(new_n380), .A3(new_n369), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G469), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G221), .B1(new_n284), .B2(G902), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G214), .B1(G237), .B2(G902), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n325), .B1(new_n323), .B2(new_n327), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n331), .A2(new_n324), .A3(new_n333), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n188), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G125), .B1(new_n352), .B2(new_n356), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT87), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n201), .A2(G224), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n400), .B(KEYINPUT88), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n397), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n352), .A2(new_n356), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n188), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(KEYINPUT87), .C1(new_n335), .C2(new_n188), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n401), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT2), .A2(G113), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT67), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT67), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT2), .A3(G113), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT2), .ZN(new_n413));
  INV_X1    g227(.A(G113), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G116), .B(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT68), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n271), .A2(G119), .ZN(new_n419));
  INV_X1    g233(.A(G119), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(G116), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n271), .A2(G119), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT68), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n417), .B1(new_n426), .B2(new_n415), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n322), .A3(new_n337), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n355), .A2(new_n321), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(new_n422), .B2(new_n425), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n414), .B1(new_n419), .B2(new_n431), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n430), .B(new_n417), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n436), .A2(new_n438), .B1(new_n439), .B2(KEYINPUT6), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(KEYINPUT6), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n437), .B(new_n441), .C1(new_n428), .C2(new_n435), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n428), .A2(new_n435), .A3(new_n437), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT86), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT86), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n428), .A2(new_n435), .A3(new_n446), .A4(new_n437), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n408), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n447), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n429), .B(new_n417), .C1(new_n432), .C2(new_n434), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n433), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n417), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n430), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n437), .B(KEYINPUT8), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n400), .A2(KEYINPUT7), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n397), .B2(new_n399), .ZN(new_n459));
  INV_X1    g273(.A(new_n458), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n406), .A2(new_n398), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n450), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n248), .ZN(new_n464));
  OAI21_X1  g278(.A(G210), .B1(G237), .B2(G902), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n449), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n408), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n445), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n318), .A2(new_n336), .A3(G101), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n410), .A2(new_n412), .ZN(new_n471));
  NOR2_X1   g285(.A1(KEYINPUT2), .A2(G113), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n422), .B(new_n425), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n417), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT68), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT68), .B1(new_n423), .B2(new_n424), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT5), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n477), .A2(new_n433), .B1(new_n415), .B2(new_n416), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n474), .A2(new_n322), .B1(new_n478), .B2(new_n430), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n441), .B1(new_n479), .B2(new_n437), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT6), .A4(new_n438), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n468), .B1(new_n469), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n450), .B2(new_n462), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n465), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n391), .B1(new_n467), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n466), .B1(new_n449), .B2(new_n464), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n465), .A3(new_n484), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n391), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n312), .B(new_n390), .C1(new_n487), .C2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(G472), .A2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT32), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(KEYINPUT71), .A2(KEYINPUT31), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT31), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n502));
  XNOR2_X1  g316(.A(G134), .B(G137), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(new_n233), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n341), .A2(G134), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n343), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT65), .A3(G131), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n504), .A2(new_n507), .B1(new_n508), .B2(new_n233), .ZN(new_n509));
  INV_X1    g323(.A(new_n404), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n427), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n335), .A2(new_n347), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n510), .B1(new_n509), .B2(KEYINPUT66), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT65), .B1(new_n506), .B2(G131), .ZN(new_n518));
  AOI211_X1 g332(.A(new_n502), .B(new_n233), .C1(new_n505), .C2(new_n343), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT66), .B(new_n346), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n516), .B(new_n513), .C1(new_n517), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n513), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT30), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n515), .B1(new_n525), .B2(new_n427), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n209), .A2(G210), .A3(new_n205), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT26), .B(G101), .Z(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(new_n532), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n527), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n501), .B1(new_n526), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n512), .B1(new_n522), .B2(new_n524), .ZN(new_n538));
  INV_X1    g352(.A(new_n501), .ZN(new_n539));
  NOR4_X1   g353(.A1(new_n538), .A2(new_n515), .A3(new_n539), .A4(new_n535), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n533), .A2(new_n534), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n392), .A2(new_n393), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n345), .B2(new_n346), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n346), .B1(new_n518), .B2(new_n519), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT66), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n404), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n545), .B1(new_n548), .B2(new_n520), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT73), .B1(new_n549), .B2(new_n512), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n513), .B1(new_n517), .B2(new_n521), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT73), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n427), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n553), .A3(new_n514), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n514), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n543), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n498), .B1(new_n541), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n523), .A2(new_n427), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n558), .B1(new_n562), .B2(new_n514), .ZN(new_n563));
  INV_X1    g377(.A(new_n559), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT29), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n542), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(G902), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n526), .B2(new_n543), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n543), .A2(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n554), .B2(new_n556), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n568), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n561), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n564), .B1(new_n554), .B2(new_n556), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n540), .A2(new_n537), .B1(new_n575), .B2(new_n543), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT32), .B1(new_n576), .B2(new_n495), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT74), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n576), .A2(new_n498), .B1(new_n572), .B2(G472), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n557), .A2(new_n559), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n516), .B1(new_n511), .B2(new_n513), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n549), .B2(new_n516), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n536), .B(new_n514), .C1(new_n582), .C2(new_n512), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n539), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n526), .A2(new_n501), .A3(new_n536), .ZN(new_n585));
  AOI22_X1  g399(.A1(new_n580), .A2(new_n542), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n497), .B1(new_n586), .B2(new_n496), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n579), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n209), .A2(G221), .A3(G234), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT79), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT22), .B(G137), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT76), .ZN(new_n594));
  INV_X1    g408(.A(G110), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(KEYINPUT24), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT24), .B(G110), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT76), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n263), .A2(G119), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n420), .A2(G128), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT75), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n598), .A2(new_n600), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT23), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT23), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT77), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n601), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n611), .A2(new_n614), .A3(G110), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n197), .B(new_n227), .C1(new_n607), .C2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n605), .A2(new_n598), .A3(new_n600), .A4(new_n606), .ZN(new_n617));
  OAI21_X1  g431(.A(G110), .B1(new_n611), .B2(new_n614), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n228), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n616), .A2(new_n619), .A3(KEYINPUT80), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT80), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n593), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n592), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n591), .B(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT80), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n616), .A2(new_n619), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n622), .A2(new_n248), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT25), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT25), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n622), .A2(new_n630), .A3(new_n248), .A4(new_n627), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n285), .B1(G234), .B2(new_n248), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT81), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n622), .A2(new_n627), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n632), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n622), .A2(KEYINPUT81), .A3(new_n627), .A4(new_n636), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n633), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n578), .A2(new_n589), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n642), .A2(KEYINPUT82), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(KEYINPUT82), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n494), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT94), .B(G101), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G3));
  AND2_X1   g461(.A1(new_n388), .A2(new_n389), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n548), .A2(new_n520), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n512), .B1(new_n649), .B2(new_n513), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n515), .B1(new_n650), .B2(new_n552), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n555), .B1(new_n651), .B2(new_n550), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n542), .B1(new_n652), .B2(new_n564), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n584), .A2(new_n585), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n496), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n586), .B2(G902), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n648), .A2(new_n656), .A3(new_n641), .A4(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n296), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n294), .A2(new_n659), .A3(new_n660), .A4(new_n295), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n260), .A2(G902), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n665), .A2(new_n666), .B1(new_n260), .B2(new_n289), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n667), .B1(new_n252), .B2(new_n259), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n391), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n467), .B2(KEYINPUT95), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT95), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n488), .A2(new_n489), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n658), .A2(new_n310), .A3(new_n669), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n221), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  OR2_X1    g492(.A1(new_n298), .A2(new_n301), .ZN(new_n679));
  INV_X1    g493(.A(new_n310), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n252), .A2(new_n259), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n391), .B1(new_n489), .B2(new_n672), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n467), .A2(new_n485), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(new_n672), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n658), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT35), .B(G107), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  OAI21_X1  g504(.A(KEYINPUT99), .B1(new_n624), .B2(KEYINPUT36), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT36), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n593), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n619), .A2(new_n691), .A3(new_n616), .A4(new_n694), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n691), .A2(new_n694), .B1(new_n619), .B2(new_n616), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n636), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n633), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n576), .A2(new_n248), .ZN(new_n700));
  AOI211_X1 g514(.A(new_n655), .B(new_n699), .C1(G472), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n493), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT37), .B(G110), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G12));
  NAND3_X1  g518(.A1(new_n388), .A2(new_n698), .A3(new_n389), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n674), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n252), .A2(new_n259), .A3(new_n679), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n306), .B1(new_n308), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AND4_X1   g524(.A1(new_n578), .A2(new_n706), .A3(new_n589), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n263), .ZN(G30));
  XOR2_X1   g526(.A(new_n709), .B(KEYINPUT39), .Z(new_n713));
  NAND2_X1  g527(.A1(new_n648), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT101), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT40), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n543), .B1(new_n538), .B2(new_n515), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n542), .A2(new_n514), .A3(new_n562), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n248), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G472), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n587), .A2(new_n561), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n490), .B(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n252), .A2(new_n259), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n679), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n699), .A2(new_n391), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n717), .A2(new_n718), .A3(new_n723), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  AOI211_X1 g546(.A(new_n667), .B(new_n709), .C1(new_n252), .C2(new_n259), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n578), .A2(new_n706), .A3(new_n589), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NOR3_X1   g549(.A1(new_n574), .A2(new_n577), .A3(KEYINPUT74), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n588), .B1(new_n579), .B2(new_n587), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n669), .A2(new_n674), .A3(new_n310), .ZN(new_n739));
  INV_X1    g553(.A(new_n389), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n248), .B1(new_n375), .B2(new_n381), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(KEYINPUT102), .A3(new_n382), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n744), .A3(G469), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n740), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n738), .A2(new_n641), .A3(new_n739), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NOR2_X1   g563(.A1(new_n686), .A2(new_n687), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n738), .A2(new_n750), .A3(new_n641), .A4(new_n746), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  NOR2_X1   g566(.A1(new_n312), .A2(new_n699), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n746), .A2(new_n685), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n738), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n382), .A2(KEYINPUT102), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n365), .A2(new_n369), .A3(new_n374), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n348), .B1(new_n376), .B2(KEYINPUT84), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n379), .A2(new_n759), .B1(new_n362), .B2(new_n364), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n758), .B1(new_n760), .B2(new_n369), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n313), .B1(new_n761), .B2(new_n248), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n745), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n680), .B(new_n389), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n671), .A2(new_n727), .A3(new_n679), .A4(new_n673), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n565), .A2(new_n543), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n496), .B1(new_n654), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n700), .B2(G472), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n641), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n733), .A3(new_n698), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n746), .A2(new_n685), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n495), .B1(new_n541), .B2(new_n768), .ZN(new_n779));
  AOI21_X1  g593(.A(G902), .B1(new_n653), .B2(new_n654), .ZN(new_n780));
  INV_X1    g594(.A(G472), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n698), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n709), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n668), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT103), .A3(new_n685), .A4(new_n746), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n778), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G125), .ZN(G27));
  NOR2_X1   g602(.A1(new_n740), .A2(new_n670), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n684), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT106), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n386), .A2(KEYINPUT104), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT104), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n365), .A2(new_n380), .A3(new_n793), .A4(new_n369), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n792), .A2(G469), .A3(new_n385), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT105), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n382), .B(new_n383), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n791), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n382), .A2(new_n383), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n795), .A2(new_n796), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT106), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n790), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n642), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n784), .A2(KEYINPUT42), .ZN(new_n807));
  AOI211_X1 g621(.A(KEYINPUT107), .B(new_n640), .C1(new_n579), .C2(new_n587), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT107), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n561), .B(new_n573), .C1(new_n655), .C2(KEYINPUT32), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n641), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n804), .B(new_n733), .C1(new_n808), .C2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n806), .A2(new_n807), .B1(new_n812), .B2(KEYINPUT42), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G131), .ZN(G33));
  NAND4_X1  g628(.A1(new_n738), .A2(new_n641), .A3(new_n710), .A4(new_n804), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G134), .ZN(G36));
  NAND2_X1  g630(.A1(new_n385), .A2(new_n386), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT45), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n313), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n792), .A2(KEYINPUT45), .A3(new_n385), .A4(new_n794), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n383), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT46), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(KEYINPUT46), .A3(new_n383), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n382), .A3(new_n827), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n389), .A3(new_n713), .ZN(new_n829));
  INV_X1    g643(.A(new_n727), .ZN(new_n830));
  INV_X1    g644(.A(new_n667), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT43), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(KEYINPUT109), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g648(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n835));
  NAND3_X1  g649(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n699), .B1(new_n657), .B2(new_n656), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(KEYINPUT44), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT44), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n490), .A2(new_n670), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT110), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n829), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(G137), .ZN(G39));
  NAND2_X1  g659(.A1(new_n578), .A2(new_n589), .ZN(new_n846));
  INV_X1    g660(.A(new_n841), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n784), .A2(new_n847), .A3(new_n641), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n828), .A2(KEYINPUT47), .A3(new_n389), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT47), .B1(new_n828), .B2(new_n389), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G140), .ZN(G42));
  NOR4_X1   g669(.A1(new_n725), .A2(new_n832), .A3(new_n670), .A4(new_n740), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n723), .A2(new_n640), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n743), .A2(new_n745), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT49), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n491), .B1(new_n490), .B2(new_n391), .ZN(new_n862));
  AOI211_X1 g676(.A(KEYINPUT89), .B(new_n670), .C1(new_n488), .C2(new_n489), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n680), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n658), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n707), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n707), .A2(new_n866), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n668), .A2(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(KEYINPUT112), .B(new_n667), .C1(new_n252), .C2(new_n259), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n867), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n865), .A2(new_n872), .B1(new_n767), .B2(new_n772), .ZN(new_n873));
  AOI22_X1  g687(.A1(new_n738), .A2(new_n754), .B1(new_n493), .B2(new_n701), .ZN(new_n874));
  AND4_X1   g688(.A1(new_n747), .A2(new_n873), .A3(new_n874), .A4(new_n751), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n643), .A2(new_n644), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n493), .ZN(new_n877));
  INV_X1    g691(.A(new_n705), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n578), .A2(new_n589), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n679), .A2(new_n709), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n830), .A2(new_n841), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT114), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n830), .A2(new_n841), .A3(new_n883), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n879), .A2(new_n885), .B1(new_n785), .B2(new_n804), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n886), .A2(new_n815), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n875), .A2(new_n877), .A3(new_n887), .A4(new_n813), .ZN(new_n888));
  INV_X1    g702(.A(new_n711), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n787), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n799), .A2(new_n803), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n698), .B2(new_n709), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n633), .A2(new_n697), .A3(KEYINPUT115), .A4(new_n783), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n740), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n766), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n891), .A2(new_n723), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n734), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT52), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n711), .B1(new_n778), .B2(new_n786), .ZN(new_n900));
  INV_X1    g714(.A(new_n898), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n861), .B1(new_n888), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n900), .B2(new_n901), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n812), .A2(KEYINPUT42), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n738), .A2(new_n641), .A3(new_n804), .A4(new_n807), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n886), .A3(new_n910), .A4(new_n815), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n874), .A2(new_n873), .A3(new_n751), .A4(new_n747), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n645), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n908), .A2(new_n913), .A3(KEYINPUT53), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n905), .A2(new_n914), .A3(KEYINPUT117), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n916), .B(new_n861), .C1(new_n888), .C2(new_n904), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OR4_X1    g735(.A1(KEYINPUT116), .A2(new_n888), .A3(new_n904), .A4(new_n861), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n905), .A2(new_n914), .A3(KEYINPUT116), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(KEYINPUT54), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT54), .B1(new_n915), .B2(new_n917), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n926), .A2(new_n919), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n305), .B1(new_n834), .B2(new_n836), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n772), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n852), .A2(new_n853), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n858), .A2(new_n740), .ZN(new_n931));
  AOI211_X1 g745(.A(new_n842), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n746), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n847), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n698), .B(new_n771), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n933), .A2(new_n725), .A3(new_n391), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT50), .B1(new_n929), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n306), .A3(new_n857), .ZN(new_n942));
  OR3_X1    g756(.A1(new_n942), .A2(new_n727), .A3(new_n831), .ZN(new_n943));
  OR3_X1    g757(.A1(new_n929), .A2(new_n940), .A3(KEYINPUT50), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n938), .A2(new_n941), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT119), .B1(new_n932), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT51), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT51), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT119), .B(new_n948), .C1(new_n932), .C2(new_n945), .ZN(new_n949));
  OAI221_X1 g763(.A(new_n303), .B1(new_n942), .B2(new_n669), .C1(new_n929), .C2(new_n777), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n808), .A2(new_n811), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n936), .B2(new_n937), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n952), .A2(KEYINPUT48), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(KEYINPUT48), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n947), .A2(new_n949), .A3(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n925), .A2(new_n927), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(G952), .A2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n860), .B1(new_n957), .B2(new_n959), .ZN(G75));
  NOR2_X1   g774(.A1(new_n469), .A2(new_n482), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n468), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT55), .Z(new_n963));
  NOR2_X1   g777(.A1(new_n918), .A2(new_n248), .ZN(new_n964));
  AOI211_X1 g778(.A(KEYINPUT56), .B(new_n963), .C1(new_n964), .C2(G210), .ZN(new_n965));
  INV_X1    g779(.A(new_n963), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n915), .A2(new_n917), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(G210), .A3(G902), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT56), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n209), .A2(G952), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n965), .A2(new_n970), .A3(new_n971), .ZN(G51));
  XOR2_X1   g786(.A(new_n383), .B(KEYINPUT57), .Z(new_n973));
  AND3_X1   g787(.A1(new_n915), .A2(KEYINPUT54), .A3(new_n917), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n926), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n761), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n823), .B(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n964), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n976), .B2(new_n978), .ZN(G54));
  NAND4_X1  g793(.A1(new_n967), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n980));
  INV_X1    g794(.A(new_n244), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n982), .A2(new_n983), .A3(new_n971), .ZN(G60));
  NAND2_X1  g798(.A1(G478), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT59), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n665), .B(new_n987), .C1(new_n974), .C2(new_n926), .ZN(new_n988));
  INV_X1    g802(.A(new_n971), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n925), .B2(new_n927), .ZN(new_n991));
  INV_X1    g805(.A(new_n665), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G63));
  OR2_X1    g807(.A1(new_n695), .A2(new_n696), .ZN(new_n994));
  NAND2_X1  g808(.A1(G217), .A2(G902), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT60), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n967), .A2(new_n994), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n635), .B1(new_n918), .B2(new_n996), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n998), .A2(new_n989), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n999), .A4(new_n989), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(G66));
  INV_X1    g818(.A(G224), .ZN(new_n1005));
  OAI21_X1  g819(.A(G953), .B1(new_n309), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n912), .A2(new_n645), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(new_n307), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT123), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n961), .B1(G898), .B2(new_n209), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NAND3_X1  g825(.A1(new_n829), .A2(new_n896), .A3(new_n951), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n900), .A2(new_n734), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(new_n813), .A3(new_n815), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n854), .A2(new_n844), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n209), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n708), .B2(new_n209), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n239), .A2(new_n240), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT124), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n525), .B(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT125), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT62), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n731), .A2(new_n1013), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n872), .ZN(new_n1026));
  NOR3_X1   g840(.A1(new_n1026), .A2(new_n714), .A3(new_n847), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n876), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g842(.A1(new_n1025), .A2(new_n844), .A3(new_n854), .A4(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n731), .A2(new_n1013), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1023), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  AND3_X1   g847(.A1(new_n854), .A2(new_n844), .A3(new_n1028), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1034), .A2(KEYINPUT125), .A3(new_n1031), .A4(new_n1025), .ZN(new_n1035));
  AOI211_X1 g849(.A(new_n307), .B(new_n1021), .C1(new_n1033), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n209), .B1(G227), .B2(G900), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n1022), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G227), .A2(G900), .ZN(new_n1039));
  AND4_X1   g853(.A1(new_n307), .A2(new_n1018), .A3(new_n1039), .A4(new_n1021), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n1038), .A2(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT126), .Z(new_n1044));
  AOI21_X1  g858(.A(new_n1044), .B1(new_n1016), .B2(new_n1007), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n526), .A2(new_n542), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n989), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1033), .A2(new_n1007), .A3(new_n1035), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1044), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n719), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1046), .A2(new_n719), .A3(new_n1043), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n922), .A2(new_n923), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g866(.A(KEYINPUT127), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OR2_X1    g868(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  AOI211_X1 g869(.A(new_n1047), .B(new_n1050), .C1(new_n1054), .C2(new_n1055), .ZN(G57));
endmodule


