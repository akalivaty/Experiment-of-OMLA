//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1209, new_n1210, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266, new_n1267;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n223), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT64), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT21), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n247), .A2(new_n212), .B1(G20), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G283), .ZN(new_n250));
  INV_X1    g0050(.A(G97), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n250), .B(new_n206), .C1(G33), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n249), .A2(KEYINPUT20), .A3(new_n252), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n248), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n247), .A2(new_n212), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n258), .C1(G1), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(new_n248), .ZN(new_n265));
  OAI21_X1  g0065(.A(G169), .B1(new_n257), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  INV_X1    g0068(.A(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT5), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT5), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT67), .B1(new_n274), .B2(new_n212), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G1), .A4(G13), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n273), .A2(new_n275), .A3(G270), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n275), .A2(G274), .A3(new_n278), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G257), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G264), .A2(G1698), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OR2_X1    g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(G303), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n274), .A2(new_n212), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT82), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT82), .A4(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n281), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n246), .B1(new_n266), .B2(new_n297), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n299), .A2(G274), .A3(new_n275), .A4(new_n278), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n300), .A2(new_n279), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n296), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n255), .A2(new_n256), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n304), .B(new_n260), .C1(new_n248), .C2(new_n264), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT21), .A4(G169), .ZN(new_n306));
  INV_X1    g0106(.A(new_n305), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n302), .A3(G179), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n298), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G200), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n307), .B1(new_n297), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G190), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n206), .A2(new_n263), .A3(KEYINPUT69), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT69), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(G20), .B2(G33), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G150), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT8), .B(G58), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n206), .A2(G33), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n206), .B2(new_n201), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n261), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n258), .A2(G50), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n261), .B1(new_n205), .B2(G20), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G50), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n213), .A2(new_n276), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n288), .A2(new_n290), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G223), .A2(G1698), .ZN(new_n332));
  INV_X1    g0132(.A(G222), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n202), .B2(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT68), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n337), .B2(new_n336), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g0140(.A1(KEYINPUT65), .A2(G45), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT65), .A2(G45), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n342), .A2(new_n343), .A3(G41), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n340), .B1(new_n344), .B2(G1), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n275), .A2(G274), .A3(new_n278), .ZN(new_n346));
  OR2_X1    g0146(.A1(KEYINPUT65), .A2(G45), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(new_n269), .A3(new_n341), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT66), .A3(new_n205), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n275), .A2(new_n278), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(G226), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n339), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n329), .B1(new_n354), .B2(G179), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n354), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n354), .A2(G200), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT72), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n325), .A2(KEYINPUT9), .A3(new_n328), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n362), .B1(new_n329), .B2(new_n363), .ZN(new_n364));
  AOI211_X1 g0164(.A(KEYINPUT71), .B(KEYINPUT9), .C1(new_n325), .C2(new_n328), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n361), .B1(new_n364), .B2(new_n365), .C1(new_n354), .C2(new_n312), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT10), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT10), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n360), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n357), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  MUX2_X1   g0172(.A(new_n223), .B(new_n225), .S(G1698), .Z(new_n373));
  AOI21_X1  g0173(.A(new_n330), .B1(new_n373), .B2(new_n331), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n285), .A2(new_n286), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(G244), .A2(new_n352), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n350), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n356), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n327), .A2(G77), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT15), .B(G87), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n385), .A2(new_n323), .B1(new_n206), .B2(new_n202), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n316), .A2(new_n318), .ZN(new_n387));
  INV_X1    g0187(.A(new_n322), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI221_X1 g0189(.A(new_n384), .B1(G77), .B2(new_n258), .C1(new_n389), .C2(new_n262), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n382), .A2(new_n383), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n379), .B2(G200), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(KEYINPUT70), .B1(G190), .B2(new_n380), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n393), .B1(KEYINPUT70), .B2(new_n392), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n372), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n259), .A2(new_n224), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT12), .ZN(new_n397));
  INV_X1    g0197(.A(new_n327), .ZN(new_n398));
  INV_X1    g0198(.A(G50), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n319), .A2(new_n399), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n323), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n261), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT11), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n397), .B1(new_n224), .B2(new_n398), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n403), .B2(new_n402), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n348), .A2(KEYINPUT66), .A3(new_n205), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT66), .B1(new_n348), .B2(new_n205), .ZN(new_n407));
  NOR3_X1   g0207(.A1(new_n406), .A2(new_n407), .A3(new_n280), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n275), .A2(G238), .A3(new_n278), .A4(new_n351), .ZN(new_n409));
  NOR2_X1   g0209(.A1(G226), .A2(G1698), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n223), .B2(G1698), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n331), .B1(G33), .B2(G97), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n409), .B1(new_n412), .B2(new_n330), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT13), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n223), .A2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G226), .B2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n417), .B2(new_n375), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n352), .A2(G238), .B1(new_n418), .B2(new_n292), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n350), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n414), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n405), .B(new_n423), .C1(new_n312), .C2(new_n422), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT73), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n405), .B(KEYINPUT76), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT14), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n408), .A2(new_n413), .A3(KEYINPUT13), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n420), .B1(new_n419), .B2(new_n350), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT74), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT74), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n422), .A2(new_n432), .A3(new_n427), .A4(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n427), .B1(new_n422), .B2(G169), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n422), .A2(new_n381), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n434), .A2(KEYINPUT75), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT75), .B1(new_n434), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n426), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n352), .A2(G232), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n350), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT77), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n350), .A2(new_n445), .A3(new_n442), .ZN(new_n446));
  OR2_X1    g0246(.A1(G223), .A2(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n331), .B(new_n447), .C1(G226), .C2(new_n282), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G87), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n330), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n444), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n356), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT16), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT7), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n331), .B2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n375), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n224), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n387), .A2(G159), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n222), .A2(new_n224), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G58), .A2(G68), .ZN(new_n461));
  OAI21_X1  g0261(.A(G20), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n454), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n331), .A2(new_n455), .A3(G20), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT7), .B1(new_n375), .B2(new_n206), .ZN(new_n466));
  OAI21_X1  g0266(.A(G68), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n463), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT16), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n464), .A2(new_n469), .A3(new_n261), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n322), .A2(new_n259), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n398), .B2(new_n322), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n450), .B1(new_n443), .B2(KEYINPUT77), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n381), .A3(new_n446), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n453), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT18), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT18), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n453), .A2(new_n479), .A3(new_n474), .A4(new_n476), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n452), .A2(new_n310), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n475), .A2(new_n312), .A3(new_n446), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n467), .A2(new_n468), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n262), .B1(new_n485), .B2(new_n454), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n472), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n481), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AOI211_X1 g0288(.A(KEYINPUT17), .B(new_n474), .C1(new_n482), .C2(new_n483), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n478), .B(new_n480), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NOR4_X1   g0290(.A1(new_n395), .A2(new_n425), .A3(new_n441), .A4(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n219), .B1(new_n288), .B2(new_n290), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT79), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g0294(.A(G1698), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G244), .B1(new_n285), .B2(new_n286), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n496), .A2(new_n494), .B1(G33), .B2(G283), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT4), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n331), .A2(G244), .A3(new_n282), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(KEYINPUT79), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n292), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(new_n278), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n300), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT80), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n217), .B1(new_n288), .B2(new_n290), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n493), .B1(new_n508), .B2(new_n282), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n495), .B(new_n497), .C1(new_n509), .C2(new_n499), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n504), .B1(new_n510), .B2(new_n292), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT80), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n507), .A2(G200), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n515), .A2(new_n251), .A3(G107), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n518), .A2(new_n206), .B1(new_n202), .B2(new_n319), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n376), .B1(new_n456), .B2(new_n457), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n261), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n258), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT78), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n522), .B(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n264), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(G97), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(G190), .B2(new_n511), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n511), .A2(new_n381), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n506), .A2(new_n356), .B1(new_n521), .B2(new_n526), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n514), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n273), .A2(new_n275), .A3(new_n278), .ZN(new_n532));
  OAI211_X1 g0332(.A(G250), .B(new_n282), .C1(new_n285), .C2(new_n286), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G294), .ZN(new_n534));
  AND2_X1   g0334(.A1(G257), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n285), .B2(new_n286), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n532), .A2(G264), .B1(new_n537), .B2(new_n292), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n381), .A3(new_n300), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n292), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n273), .A2(new_n275), .A3(G264), .A4(new_n278), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n300), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n356), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n206), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  AOI21_X1  g0350(.A(G20), .B1(new_n288), .B2(new_n290), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G87), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n206), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n549), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT24), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n331), .A2(new_n550), .A3(new_n206), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n559), .A2(new_n560), .A3(new_n549), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n262), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n258), .A2(new_n563), .A3(G107), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n563), .B1(new_n258), .B2(G107), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n525), .A2(G107), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n539), .B(new_n543), .C1(new_n562), .C2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n267), .A2(G1), .A3(G274), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n219), .B1(new_n267), .B2(G1), .ZN(new_n572));
  AND4_X1   g0372(.A1(new_n275), .A2(new_n571), .A3(new_n278), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n225), .A2(new_n282), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n217), .A2(G1698), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n285), .C2(new_n286), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n330), .B1(new_n576), .B2(new_n544), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n570), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n275), .A2(new_n571), .A3(new_n278), .A4(new_n572), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G238), .A2(G1698), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n217), .B2(G1698), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n581), .A2(new_n331), .B1(G33), .B2(G116), .ZN(new_n582));
  OAI211_X1 g0382(.A(KEYINPUT81), .B(new_n579), .C1(new_n582), .C2(new_n330), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n356), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n551), .A2(G68), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n218), .A2(new_n251), .A3(new_n376), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n415), .A2(new_n206), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT19), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n323), .B2(new_n251), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n261), .B1(new_n259), .B2(new_n385), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n264), .B2(new_n385), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n585), .B(new_n594), .C1(G179), .C2(new_n584), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n538), .A2(new_n312), .A3(new_n300), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n542), .A2(new_n310), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n559), .A2(new_n560), .A3(new_n549), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n560), .B1(new_n559), .B2(new_n549), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n261), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n598), .A2(new_n601), .A3(new_n567), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n584), .A2(G200), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n578), .A2(new_n583), .A3(G190), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n525), .A2(G87), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n603), .A2(new_n593), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  AND4_X1   g0406(.A1(new_n569), .A2(new_n595), .A3(new_n602), .A4(new_n606), .ZN(new_n607));
  AND4_X1   g0407(.A1(new_n315), .A2(new_n491), .A3(new_n531), .A4(new_n607), .ZN(G372));
  OAI21_X1  g0408(.A(new_n579), .B1(new_n582), .B2(new_n330), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n356), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n594), .B(new_n610), .C1(G179), .C2(new_n584), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(G200), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n604), .A2(new_n593), .A3(new_n605), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n530), .A2(new_n529), .ZN(new_n615));
  OR3_X1    g0415(.A1(new_n614), .A2(new_n615), .A3(KEYINPUT26), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n595), .A2(new_n606), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT26), .B1(new_n617), .B2(new_n615), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n616), .A2(KEYINPUT83), .A3(new_n611), .A4(new_n618), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n531), .A2(new_n602), .A3(new_n611), .A4(new_n613), .ZN(new_n623));
  INV_X1    g0423(.A(new_n309), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n569), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n491), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n478), .A2(new_n480), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT73), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n424), .B(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n391), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n441), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n488), .A2(new_n489), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n369), .A2(new_n371), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n357), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n629), .A2(new_n639), .ZN(G369));
  INV_X1    g0440(.A(new_n569), .ZN(new_n641));
  INV_X1    g0441(.A(new_n602), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n601), .A2(new_n567), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(G213), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n649), .B(KEYINPUT85), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G343), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n643), .B1(new_n645), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n651), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n641), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n305), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n315), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n624), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g0458(.A(KEYINPUT86), .B(G330), .Z(new_n659));
  AND3_X1   g0459(.A1(new_n658), .A2(KEYINPUT87), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(KEYINPUT87), .B1(new_n658), .B2(new_n659), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n641), .A2(new_n651), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n624), .A2(new_n653), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n643), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(G399));
  INV_X1    g0466(.A(new_n209), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G41), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n215), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n587), .A2(G116), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n668), .A2(new_n672), .A3(new_n205), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n670), .B1(new_n674), .B2(KEYINPUT88), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(KEYINPUT88), .B2(new_n674), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n619), .A2(new_n620), .B1(new_n623), .B2(new_n625), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n653), .B1(new_n678), .B2(new_n622), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT29), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR3_X1    g0481(.A1(new_n617), .A2(new_n615), .A3(KEYINPUT26), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT26), .B1(new_n614), .B2(new_n615), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n626), .A2(new_n611), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n651), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n511), .A2(new_n538), .A3(new_n578), .A4(new_n583), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT89), .B1(new_n297), .B2(G179), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT90), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT89), .A4(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT30), .A4(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n308), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n578), .A2(new_n538), .A3(new_n583), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n511), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT90), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n542), .A2(new_n381), .A3(new_n609), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n701), .A2(new_n511), .A3(new_n297), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n698), .B2(new_n699), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n694), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n653), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n607), .A2(new_n315), .A3(new_n531), .A4(new_n651), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n705), .A2(KEYINPUT31), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n704), .A2(new_n653), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT31), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n707), .A2(new_n706), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n659), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n688), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n677), .B1(new_n716), .B2(G1), .ZN(G364));
  AOI21_X1  g0517(.A(new_n212), .B1(G20), .B2(new_n356), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n310), .A2(G179), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n206), .A2(G190), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(G283), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n206), .A2(new_n312), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n381), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G322), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n721), .A2(new_n726), .ZN(new_n729));
  INV_X1    g0529(.A(G311), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n727), .A2(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G179), .A2(G200), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI211_X1 g0534(.A(new_n724), .B(new_n731), .C1(G329), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n206), .B1(new_n732), .B2(G190), .ZN(new_n736));
  INV_X1    g0536(.A(G294), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n725), .A2(new_n720), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n375), .B1(new_n739), .B2(new_n289), .ZN(new_n740));
  NAND3_X1  g0540(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n312), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n738), .B(new_n740), .C1(G326), .C2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n741), .A2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT96), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT33), .B(G317), .Z(new_n750));
  OAI211_X1 g0550(.A(new_n735), .B(new_n743), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n202), .A2(new_n729), .B1(new_n722), .B2(new_n376), .ZN(new_n752));
  INV_X1    g0552(.A(new_n742), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n753), .A2(new_n399), .B1(new_n736), .B2(new_n251), .ZN(new_n754));
  INV_X1    g0554(.A(new_n727), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n752), .B(new_n754), .C1(G58), .C2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n331), .B1(new_n739), .B2(new_n218), .ZN(new_n757));
  XOR2_X1   g0557(.A(new_n757), .B(KEYINPUT95), .Z(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n733), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  OAI21_X1  g0561(.A(G68), .B1(new_n747), .B2(new_n748), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n756), .A2(new_n758), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n719), .B1(new_n751), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G13), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n205), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n668), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT92), .Z(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT94), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n718), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n244), .A2(new_n267), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n667), .A2(new_n331), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n347), .A2(new_n341), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n215), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n776), .B1(new_n779), .B2(KEYINPUT93), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(KEYINPUT93), .B2(new_n779), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n667), .A2(new_n375), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G355), .B1(new_n248), .B2(new_n667), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n764), .B(new_n771), .C1(new_n775), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT97), .Z(new_n786));
  INV_X1    g0586(.A(new_n774), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n658), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT98), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n660), .A2(new_n661), .ZN(new_n790));
  INV_X1    g0590(.A(new_n769), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(new_n659), .C2(new_n658), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n718), .A2(new_n772), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n771), .B1(new_n202), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n749), .A2(KEYINPUT100), .ZN(new_n799));
  OAI21_X1  g0599(.A(G283), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n375), .B1(new_n736), .B2(new_n251), .C1(new_n218), .C2(new_n722), .ZN(new_n801));
  INV_X1    g0601(.A(new_n729), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G116), .A2(new_n802), .B1(new_n734), .B2(G311), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n803), .B1(new_n376), .B2(new_n739), .C1(new_n737), .C2(new_n727), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n801), .B(new_n804), .C1(G303), .C2(new_n742), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G143), .A2(new_n755), .B1(new_n802), .B2(G159), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n807), .B2(new_n753), .C1(new_n749), .C2(new_n320), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n720), .A2(new_n721), .A3(G68), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n331), .ZN(new_n811));
  INV_X1    g0611(.A(G132), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n739), .A2(new_n399), .B1(new_n733), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n736), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n813), .C1(G58), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n800), .A2(new_n805), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n653), .A2(new_n390), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n394), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n391), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n634), .A2(new_n651), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n797), .B1(new_n719), .B2(new_n816), .C1(new_n822), .C2(new_n773), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n627), .A2(new_n822), .A3(new_n651), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n821), .B(KEYINPUT101), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n679), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n769), .B1(new_n827), .B2(new_n714), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n827), .A2(new_n714), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n823), .B1(new_n829), .B2(new_n830), .ZN(G384));
  OAI21_X1  g0631(.A(G77), .B1(new_n222), .B2(new_n224), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n832), .A2(new_n215), .B1(G50), .B2(new_n224), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(G1), .A3(new_n765), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT102), .ZN(new_n835));
  INV_X1    g0635(.A(new_n518), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n248), .B(new_n214), .C1(new_n836), .C2(KEYINPUT35), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT35), .B2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT36), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n434), .A2(new_n437), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT75), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n434), .A2(KEYINPUT75), .A3(new_n437), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n426), .B(new_n653), .C1(new_n846), .C2(new_n425), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n426), .A2(new_n653), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n440), .A2(new_n633), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n820), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n824), .B2(new_n851), .ZN(new_n852));
  AND4_X1   g0652(.A1(new_n312), .A2(new_n444), .A3(new_n446), .A4(new_n451), .ZN(new_n853));
  AOI21_X1  g0653(.A(G200), .B1(new_n475), .B2(new_n446), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n487), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n474), .A2(new_n650), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n477), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT37), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n855), .A2(new_n477), .A3(new_n859), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT103), .ZN(new_n862));
  INV_X1    g0662(.A(new_n650), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n487), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n861), .A2(new_n862), .B1(new_n490), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n860), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n484), .B2(new_n487), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n859), .B1(new_n868), .B2(new_n477), .ZN(new_n869));
  INV_X1    g0669(.A(new_n860), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n862), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n864), .B1(new_n636), .B2(new_n630), .ZN(new_n872));
  AND4_X1   g0672(.A1(KEYINPUT38), .A2(new_n871), .A3(new_n866), .A4(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n852), .A2(new_n874), .B1(new_n631), .B2(new_n650), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n872), .A3(new_n866), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n865), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n858), .A2(KEYINPUT104), .A3(new_n860), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n857), .A2(new_n884), .A3(KEYINPUT37), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(KEYINPUT105), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n872), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT105), .B1(new_n883), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n880), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n882), .B1(new_n890), .B2(KEYINPUT39), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n440), .A2(new_n653), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n875), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n687), .A2(new_n491), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n639), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n821), .B1(new_n847), .B2(new_n849), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n711), .A2(KEYINPUT106), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT106), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n709), .A2(new_n899), .A3(new_n710), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n708), .A2(new_n898), .A3(new_n712), .A4(new_n900), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n897), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT40), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n901), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n904), .B1(new_n874), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n491), .A2(new_n901), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n659), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n896), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n205), .B2(new_n766), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n896), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n841), .B1(new_n913), .B2(new_n914), .ZN(G367));
  NAND2_X1  g0715(.A1(new_n653), .A2(new_n527), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n531), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n641), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n653), .B1(new_n918), .B2(new_n615), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n615), .A2(new_n651), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(new_n665), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n922), .B2(KEYINPUT42), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(KEYINPUT42), .B2(new_n922), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n651), .B1(new_n593), .B2(new_n605), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n614), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n611), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n925), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n931), .B(new_n932), .Z(new_n933));
  INV_X1    g0733(.A(new_n662), .ZN(new_n934));
  INV_X1    g0734(.A(new_n921), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n933), .B(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n668), .B(KEYINPUT41), .Z(new_n938));
  OAI21_X1  g0738(.A(new_n665), .B1(new_n655), .B2(new_n664), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n790), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n790), .A2(new_n939), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n688), .A2(new_n714), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n665), .A2(new_n663), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n921), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT44), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n921), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT45), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n946), .A2(new_n662), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n948), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n934), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n943), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n938), .B1(new_n955), .B2(new_n716), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n937), .B1(new_n956), .B2(new_n768), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n929), .A2(new_n787), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n777), .A2(new_n236), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(new_n775), .C1(new_n209), .C2(new_n385), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n727), .A2(new_n320), .B1(new_n729), .B2(new_n399), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n739), .A2(new_n222), .B1(new_n733), .B2(new_n807), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n736), .A2(new_n224), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n331), .B1(new_n722), .B2(new_n202), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G143), .C2(new_n742), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n798), .A2(new_n799), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n963), .B(new_n966), .C1(new_n967), .C2(new_n759), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n727), .A2(new_n289), .B1(new_n729), .B2(new_n723), .ZN(new_n969));
  INV_X1    g0769(.A(new_n739), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(G116), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT46), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n375), .B1(new_n722), .B2(new_n251), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n969), .B(new_n973), .C1(G317), .C2(new_n734), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n971), .A2(new_n972), .B1(new_n742), .B2(G311), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n376), .C2(new_n736), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n967), .A2(new_n737), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI211_X1 g0779(.A(new_n770), .B(new_n960), .C1(new_n979), .C2(new_n719), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT108), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n958), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n957), .A2(new_n983), .ZN(G387));
  AOI21_X1  g0784(.A(new_n331), .B1(new_n734), .B2(G326), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n739), .A2(new_n737), .B1(new_n736), .B2(new_n723), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G317), .A2(new_n755), .B1(new_n802), .B2(G303), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n728), .B2(new_n753), .C1(new_n967), .C2(new_n730), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT48), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n989), .B2(new_n988), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT49), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n985), .B1(new_n248), .B2(new_n722), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n749), .A2(new_n322), .B1(new_n224), .B2(new_n729), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT109), .Z(new_n996));
  NAND2_X1  g0796(.A1(new_n970), .A2(G77), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n733), .B2(new_n320), .C1(new_n399), .C2(new_n727), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n736), .A2(new_n385), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n331), .B1(new_n722), .B2(new_n251), .C1(new_n753), .C2(new_n759), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n996), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n718), .B1(new_n994), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n233), .A2(new_n778), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1003), .A2(new_n777), .B1(new_n672), .B2(new_n782), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n388), .A2(new_n399), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT50), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n267), .B1(new_n224), .B2(new_n202), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1006), .A2(new_n672), .A3(new_n1007), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1004), .A2(new_n1008), .B1(G107), .B2(new_n209), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n771), .B1(new_n1009), .B2(new_n775), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1002), .B(new_n1010), .C1(new_n655), .C2(new_n787), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n940), .A2(new_n768), .A3(new_n941), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n716), .B1(new_n940), .B2(new_n941), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n942), .A2(new_n668), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(G393));
  NAND3_X1  g0815(.A1(new_n952), .A2(new_n768), .A3(new_n949), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n775), .B1(new_n251), .B2(new_n209), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n240), .B2(new_n777), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n331), .B1(new_n736), .B2(new_n202), .C1(new_n218), .C2(new_n722), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n734), .A2(G143), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n224), .B2(new_n739), .C1(new_n322), .C2(new_n729), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n755), .A2(G159), .B1(G150), .B2(new_n742), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1019), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n1022), .B2(new_n1023), .C1(new_n967), .C2(new_n399), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n742), .A2(G317), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n730), .B2(new_n727), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n739), .A2(new_n723), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n729), .A2(new_n737), .B1(new_n733), .B2(new_n728), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n375), .B1(new_n736), .B2(new_n248), .C1(new_n376), .C2(new_n722), .ZN(new_n1034));
  NOR4_X1   g0834(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n1028), .B2(new_n1030), .C1(new_n967), .C2(new_n289), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1025), .A2(KEYINPUT111), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1026), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n771), .B(new_n1018), .C1(new_n1038), .C2(new_n718), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n935), .B2(new_n787), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1016), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n952), .A2(new_n949), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n942), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1043), .B(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n955), .A2(new_n668), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1041), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G390));
  AOI21_X1  g0848(.A(new_n851), .B1(new_n679), .B2(new_n822), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n850), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(KEYINPUT114), .B1(new_n1051), .B2(new_n892), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n888), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n872), .A3(new_n886), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n873), .B1(new_n1054), .B2(new_n878), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n881), .B1(new_n1055), .B2(new_n876), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT114), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n892), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n852), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1052), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n685), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n851), .B1(new_n1061), .B2(new_n819), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n890), .B(new_n1058), .C1(new_n1062), .C2(new_n1050), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n713), .A2(new_n850), .A3(new_n659), .A4(new_n822), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n901), .A2(G330), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n897), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1065), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n491), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n895), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1050), .B1(new_n714), .B2(new_n821), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n851), .B2(new_n824), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1067), .A2(new_n826), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1062), .B(new_n1064), .C1(new_n1076), .C2(new_n850), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1069), .A2(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1068), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1079), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1080), .A2(new_n1085), .A3(new_n668), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n768), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n770), .B1(new_n388), .B2(new_n795), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n375), .B1(new_n739), .B2(new_n218), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n810), .B1(new_n733), .B2(new_n737), .C1(new_n251), .C2(new_n729), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G283), .C2(new_n742), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n727), .A2(new_n248), .B1(new_n736), .B2(new_n202), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT116), .Z(new_n1093));
  OAI211_X1 g0893(.A(new_n1091), .B(new_n1093), .C1(new_n967), .C2(new_n376), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n967), .A2(new_n807), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n729), .A2(new_n1096), .B1(new_n733), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n753), .A2(new_n1099), .B1(new_n736), .B2(new_n759), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(G132), .C2(new_n755), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n970), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT53), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n739), .B2(new_n320), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n331), .B1(new_n722), .B2(new_n399), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1102), .A2(new_n1104), .B1(KEYINPUT115), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1101), .B(new_n1106), .C1(KEYINPUT115), .C2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1094), .B1(new_n1095), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1088), .B1(new_n1108), .B2(new_n718), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n891), .B2(new_n773), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1086), .A2(new_n1087), .A3(new_n1110), .ZN(G378));
  NAND2_X1  g0911(.A1(new_n1085), .A2(new_n1072), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n372), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n372), .A2(new_n1114), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n650), .A2(new_n329), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1115), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AND4_X1   g0921(.A1(G330), .A2(new_n903), .A3(new_n906), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(G330), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n897), .B(new_n901), .C1(new_n867), .C2(new_n873), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n904), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1121), .B1(new_n1125), .B2(new_n903), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n893), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n903), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1121), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n879), .A2(new_n880), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1051), .A2(new_n1131), .B1(new_n630), .B2(new_n863), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1125), .A2(new_n903), .A3(new_n1121), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1127), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(KEYINPUT57), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n669), .B1(new_n1112), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1071), .B1(new_n1083), .B2(new_n1078), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(KEYINPUT120), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1130), .A2(new_n1133), .A3(new_n1142), .A4(new_n1134), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(KEYINPUT119), .A3(new_n1127), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1127), .A2(KEYINPUT119), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n1146), .B2(new_n1133), .ZN(new_n1147));
  AND4_X1   g0947(.A1(new_n1142), .A2(new_n1130), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1140), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1139), .B1(new_n1150), .B2(KEYINPUT57), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n791), .B1(new_n399), .B2(new_n794), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT118), .Z(new_n1153));
  NOR2_X1   g0953(.A1(new_n749), .A2(new_n251), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n742), .A2(G116), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n964), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n331), .A2(G41), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n997), .A4(new_n1157), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n722), .A2(new_n222), .B1(new_n733), .B2(new_n723), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n727), .A2(new_n376), .B1(new_n729), .B2(new_n385), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1154), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1161), .A2(KEYINPUT58), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(G33), .A2(G41), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1157), .A2(G50), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT117), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n1099), .A2(new_n727), .B1(new_n739), .B2(new_n1096), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G137), .B2(new_n802), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n814), .A2(G150), .B1(G125), .B2(new_n742), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n749), .C2(new_n812), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  INV_X1    g0971(.A(G124), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1163), .B1(new_n733), .B2(new_n1172), .C1(new_n759), .C2(new_n722), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1170), .B2(KEYINPUT59), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1171), .A2(new_n1174), .B1(new_n1161), .B2(KEYINPUT58), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1166), .A2(new_n1175), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1153), .B1(new_n719), .B2(new_n1176), .C1(new_n1129), .C2(new_n773), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1149), .A2(new_n1144), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n768), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1151), .A2(new_n1180), .ZN(G375));
  NAND2_X1  g0981(.A1(new_n1050), .A2(new_n772), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n331), .B1(new_n736), .B2(new_n399), .C1(new_n222), .C2(new_n722), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G137), .A2(new_n755), .B1(new_n734), .B2(G128), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n320), .B2(new_n729), .C1(new_n759), .C2(new_n739), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n1183), .B(new_n1185), .C1(G132), .C2(new_n742), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n967), .B2(new_n1096), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n999), .B1(G283), .B2(new_n755), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT121), .Z(new_n1189));
  OAI22_X1  g0989(.A1(new_n729), .A2(new_n376), .B1(new_n733), .B2(new_n289), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n375), .B1(new_n722), .B2(new_n202), .C1(new_n753), .C2(new_n737), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(G97), .C2(new_n970), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1189), .B(new_n1192), .C1(new_n248), .C2(new_n967), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n719), .B1(new_n1187), .B2(new_n1193), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n771), .B(new_n1194), .C1(new_n224), .C2(new_n796), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT122), .Z(new_n1196));
  AOI22_X1  g0996(.A1(new_n1078), .A2(new_n768), .B1(new_n1182), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n938), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1079), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1072), .A2(new_n1078), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(G381));
  XNOR2_X1  g1001(.A(G375), .B(KEYINPUT123), .ZN(new_n1202));
  INV_X1    g1002(.A(G378), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n957), .A2(new_n1047), .A3(new_n983), .ZN(new_n1204));
  OR2_X1    g1004(.A1(G393), .A2(G396), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1204), .A2(G381), .A3(G384), .A4(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1202), .A2(new_n1203), .A3(new_n1206), .ZN(G407));
  INV_X1    g1007(.A(G213), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(G343), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1202), .A2(new_n1203), .A3(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(G407), .A2(new_n1210), .A3(G213), .ZN(G409));
  AOI21_X1  g1011(.A(new_n1047), .B1(new_n957), .B2(new_n983), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  XOR2_X1   g1013(.A(G393), .B(G396), .Z(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1213), .A2(new_n1215), .A3(KEYINPUT126), .A4(new_n1204), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1204), .A2(KEYINPUT126), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1214), .B1(new_n1217), .B2(new_n1212), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT61), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1200), .A2(KEYINPUT60), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1200), .A2(KEYINPUT60), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n668), .A3(new_n1079), .A4(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1197), .ZN(new_n1224));
  INV_X1    g1024(.A(G384), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(G384), .A3(new_n1197), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1209), .A2(G2897), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1228), .B(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1150), .A2(new_n1198), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1178), .B1(new_n1136), .B2(new_n768), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G378), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT57), .B1(new_n1179), .B2(new_n1112), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n668), .B1(new_n1140), .B2(new_n1137), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G378), .B(new_n1180), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT124), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1151), .A2(new_n1238), .A3(G378), .A4(new_n1180), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1233), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1230), .B1(new_n1240), .B2(new_n1209), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1240), .A2(new_n1209), .A3(new_n1228), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1220), .B(new_n1241), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1233), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1209), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1228), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1219), .B1(new_n1244), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT125), .B1(new_n1242), .B2(KEYINPUT63), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1250), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1216), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1258), .B1(new_n1259), .B2(new_n1230), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1242), .A2(KEYINPUT63), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1253), .A2(new_n1256), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1252), .A2(new_n1262), .ZN(G405));
  AOI21_X1  g1063(.A(G378), .B1(new_n1151), .B2(new_n1180), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1245), .A2(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(new_n1219), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1267), .B(new_n1249), .ZN(G402));
endmodule


