//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039, new_n1040;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(G43gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(G43gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT89), .ZN(new_n218));
  NAND2_X1  g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(KEYINPUT89), .B1(new_n215), .B2(new_n217), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n212), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n223), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n215), .A2(new_n217), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n209), .B2(new_n210), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT90), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n215), .A2(new_n217), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n230), .A3(KEYINPUT17), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT91), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n222), .A2(new_n230), .A3(KEYINPUT91), .A4(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G15gat), .B(G22gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT16), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(G1gat), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G1gat), .B2(new_n236), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G8gat), .ZN(new_n240));
  INV_X1    g039(.A(G8gat), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n238), .B(new_n241), .C1(G1gat), .C2(new_n236), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n222), .A2(new_n230), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n235), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT92), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n235), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n243), .A2(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(G229gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT18), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NOR3_X1   g056(.A1(new_n252), .A2(new_n257), .A3(new_n254), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n235), .A2(new_n246), .A3(new_n249), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n249), .B1(new_n235), .B2(new_n246), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n243), .B(new_n244), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n263), .B(new_n253), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n207), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n257), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n269), .A2(new_n261), .A3(new_n265), .A4(new_n206), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n267), .A2(new_n270), .A3(KEYINPUT94), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT94), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n207), .C1(new_n256), .C2(new_n266), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G225gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT76), .B(G162gat), .ZN(new_n277));
  INV_X1    g076(.A(G155gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT2), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G141gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .A4(G148gat), .ZN(new_n289));
  OR2_X1    g088(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(G141gat), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT73), .B(G141gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n288), .B1(new_n294), .B2(G148gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n279), .B(new_n283), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n284), .A2(G148gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(KEYINPUT2), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n282), .A2(KEYINPUT72), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(G155gat), .A3(G162gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n281), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(G134gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G127gat), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n307), .A2(KEYINPUT1), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G113gat), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n296), .A2(new_n306), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n285), .A2(new_n287), .A3(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n292), .A3(new_n289), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n281), .A2(new_n282), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT76), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G162gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n280), .A2(KEYINPUT76), .ZN(new_n330));
  OAI21_X1  g129(.A(G155gat), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n331), .B2(KEYINPUT2), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n305), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n276), .B1(new_n323), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n335), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n321), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n280), .A2(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n328), .A2(G162gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n278), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT2), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n283), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n289), .A2(new_n292), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n325), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n347), .B2(new_n305), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n275), .B1(new_n348), .B2(new_n322), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT81), .B1(new_n349), .B2(new_n337), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n293), .A2(new_n295), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n351), .B(new_n306), .C1(new_n352), .C2(new_n345), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n296), .A2(new_n306), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n321), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n276), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n322), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n361), .B1(new_n333), .B2(new_n321), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT79), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n333), .A2(new_n368), .A3(new_n321), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n364), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n339), .A2(new_n350), .B1(new_n360), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT82), .B(KEYINPUT0), .Z(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT83), .ZN(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G57gat), .B(G85gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AND4_X1   g177(.A1(new_n355), .A2(new_n296), .A3(new_n351), .A4(new_n306), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n355), .B1(new_n333), .B2(new_n351), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n359), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n322), .A2(new_n368), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n333), .A2(new_n321), .A3(new_n362), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n338), .A2(new_n276), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT84), .B1(new_n371), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n369), .B1(new_n365), .B2(new_n366), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n363), .A2(KEYINPUT79), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n381), .B(new_n275), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n336), .B1(new_n335), .B2(new_n338), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n349), .A2(KEYINPUT81), .A3(new_n337), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n382), .A2(new_n383), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n357), .B2(new_n359), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n377), .B1(new_n397), .B2(new_n385), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n388), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n386), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n377), .B1(new_n371), .B2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n388), .A2(new_n399), .A3(KEYINPUT85), .A4(new_n400), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT86), .B1(new_n405), .B2(new_n400), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n378), .B1(new_n394), .B2(new_n386), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT86), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT6), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  INV_X1    g214(.A(G190gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(G183gat), .ZN(new_n417));
  INV_X1    g216(.A(G183gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(G190gat), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT24), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G169gat), .ZN(new_n421));
  INV_X1    g220(.A(G176gat), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT64), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT64), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(G169gat), .A3(G176gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT23), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(new_n421), .A3(new_n422), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(G183gat), .A2(G190gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(KEYINPUT24), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n415), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(G183gat), .B(G190gat), .Z(new_n436));
  AOI22_X1  g235(.A1(new_n436), .A2(KEYINPUT24), .B1(new_n423), .B2(new_n425), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT24), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n429), .A2(new_n430), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(KEYINPUT25), .A3(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT27), .B(G183gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n416), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n418), .A2(KEYINPUT27), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G183gat), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n446), .A3(new_n416), .ZN(new_n447));
  XNOR2_X1  g246(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(G169gat), .A2(G176gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT26), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n432), .B1(new_n452), .B2(new_n426), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n435), .A2(new_n440), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT69), .B(KEYINPUT29), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n414), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n426), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n458), .A2(new_n449), .A3(new_n433), .A4(new_n443), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT25), .B1(new_n437), .B2(new_n439), .ZN(new_n460));
  AND4_X1   g259(.A1(KEYINPUT25), .A2(new_n439), .A3(new_n420), .A4(new_n426), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n414), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G211gat), .B(G218gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n467));
  XNOR2_X1  g266(.A(G197gat), .B(G204gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(G211gat), .A2(G218gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT22), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT68), .B(new_n466), .C1(new_n473), .C2(new_n474), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n465), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G8gat), .B(G36gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(G64gat), .B(G92gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n481), .B(new_n482), .Z(new_n483));
  NOR3_X1   g282(.A1(new_n454), .A2(KEYINPUT70), .A3(new_n414), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT29), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n463), .B1(new_n462), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n462), .B2(new_n463), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n480), .B(new_n483), .C1(new_n490), .C2(new_n479), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT30), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(KEYINPUT71), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n479), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n457), .B2(new_n464), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n462), .A2(new_n488), .A3(new_n463), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n464), .A2(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n486), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n500), .B2(new_n496), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n501), .A2(new_n483), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n493), .A2(new_n495), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n496), .B1(new_n357), .B2(new_n455), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n477), .A2(new_n485), .A3(new_n478), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n333), .B1(new_n507), .B2(new_n351), .ZN(new_n508));
  OAI211_X1 g307(.A(G228gat), .B(G233gat), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n351), .B1(new_n479), .B2(new_n456), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n358), .ZN(new_n511));
  NAND2_X1  g310(.A1(G228gat), .A2(G233gat), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n456), .B1(new_n354), .B2(new_n356), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n511), .B(new_n512), .C1(new_n496), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G78gat), .B(G106gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n516), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n357), .A2(new_n455), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n508), .B1(new_n521), .B2(new_n479), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n514), .B(new_n520), .C1(new_n522), .C2(new_n512), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n519), .ZN(new_n525));
  INV_X1    g324(.A(new_n523), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n520), .B1(new_n509), .B2(new_n514), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT34), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(G15gat), .B(G43gat), .Z(new_n533));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(G227gat), .ZN(new_n536));
  INV_X1    g335(.A(G233gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n462), .A2(new_n340), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n459), .B(new_n321), .C1(new_n460), .C2(new_n461), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n535), .B1(new_n542), .B2(KEYINPUT33), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  AOI221_X4 g346(.A(new_n544), .B1(KEYINPUT33), .B2(new_n535), .C1(new_n547), .C2(new_n538), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n532), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI22_X1  g348(.A1(new_n547), .A2(new_n538), .B1(KEYINPUT66), .B2(KEYINPUT34), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n541), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n435), .A2(new_n440), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n321), .B1(new_n553), .B2(new_n459), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n538), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT32), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n558), .A3(new_n535), .ZN(new_n559));
  INV_X1    g358(.A(new_n532), .ZN(new_n560));
  INV_X1    g359(.A(new_n535), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n555), .B(KEYINPUT32), .C1(new_n557), .C2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n549), .A2(new_n551), .A3(new_n563), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n546), .A2(new_n532), .A3(new_n548), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n560), .B1(new_n559), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n550), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n529), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n413), .A2(new_n505), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n504), .B1(new_n564), .B2(new_n567), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n529), .A2(KEYINPUT35), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n388), .A2(new_n405), .A3(new_n399), .A4(new_n400), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n408), .A3(new_n411), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n348), .A2(new_n322), .A3(new_n275), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT39), .B(new_n577), .C1(new_n397), .C2(new_n275), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n381), .A2(new_n384), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n276), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n378), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n578), .A2(KEYINPUT40), .A3(new_n581), .A4(new_n378), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n587), .A2(new_n405), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n583), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n504), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n529), .ZN(new_n591));
  INV_X1    g390(.A(new_n483), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n480), .B1(new_n490), .B2(new_n479), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(KEYINPUT37), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n501), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT38), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n483), .B1(new_n501), .B2(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n500), .A2(new_n479), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n595), .B1(new_n465), .B2(new_n496), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT38), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT88), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT88), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n491), .B(new_n597), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n590), .B(new_n591), .C1(new_n604), .C2(new_n574), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT36), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n565), .A2(new_n566), .A3(new_n550), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n551), .B1(new_n549), .B2(new_n563), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n567), .A2(KEYINPUT36), .A3(new_n564), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n504), .B1(new_n407), .B2(new_n412), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n605), .B(new_n612), .C1(new_n613), .C2(new_n591), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n274), .B1(new_n576), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n244), .A2(new_n245), .ZN(new_n619));
  XOR2_X1   g418(.A(G99gat), .B(G106gat), .Z(new_n620));
  NAND2_X1  g419(.A1(G85gat), .A2(G92gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT98), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .A4(KEYINPUT7), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT8), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT100), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G85gat), .ZN(new_n632));
  INV_X1    g431(.A(G92gat), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n626), .A2(new_n628), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT99), .B1(new_n621), .B2(KEYINPUT7), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT7), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n637), .B1(new_n621), .B2(KEYINPUT98), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n624), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n620), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n624), .ZN(new_n641));
  INV_X1    g440(.A(new_n636), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT100), .B(G85gat), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n644), .A2(new_n633), .B1(KEYINPUT8), .B2(new_n627), .ZN(new_n645));
  INV_X1    g444(.A(new_n620), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n646), .A4(new_n626), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n235), .A2(new_n619), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n648), .ZN(new_n650));
  AND2_X1   g449(.A1(G232gat), .A2(G233gat), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n650), .A2(new_n244), .B1(KEYINPUT41), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n618), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n649), .A2(new_n618), .A3(new_n652), .ZN(new_n655));
  XOR2_X1   g454(.A(G134gat), .B(G162gat), .Z(new_n656));
  NOR2_X1   g455(.A1(new_n651), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(KEYINPUT102), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n655), .B2(new_n653), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(KEYINPUT101), .B(new_n658), .C1(new_n655), .C2(new_n653), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(G57gat), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT95), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT95), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G57gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n671), .A3(G64gat), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n668), .B2(G64gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(G71gat), .A2(G78gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT9), .ZN(new_n675));
  INV_X1    g474(.A(G71gat), .ZN(new_n676));
  INV_X1    g475(.A(G78gat), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n668), .A2(G64gat), .ZN(new_n679));
  INV_X1    g478(.A(G64gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(G57gat), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT9), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(G71gat), .B(G78gat), .Z(new_n683));
  AOI22_X1  g482(.A1(new_n673), .A2(new_n678), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(KEYINPUT21), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n243), .B1(KEYINPUT21), .B2(new_n684), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  XNOR2_X1  g488(.A(G127gat), .B(G155gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g490(.A1(G231gat), .A2(G233gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT96), .Z(new_n693));
  XNOR2_X1  g492(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(G183gat), .B(G211gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n689), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n667), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(G230gat), .A2(G233gat), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n640), .A2(new_n684), .A3(new_n647), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n684), .B1(new_n640), .B2(new_n647), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT10), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n640), .A2(new_n684), .A3(new_n647), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT10), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n699), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n699), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n700), .B2(new_n701), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g508(.A(G120gat), .B(G148gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT103), .ZN(new_n711));
  XOR2_X1   g510(.A(G176gat), .B(G204gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n713), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n616), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n408), .A2(new_n411), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n409), .B1(new_n401), .B2(new_n402), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(new_n406), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g524(.A(KEYINPUT16), .B(G8gat), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n615), .A2(new_n504), .A3(new_n718), .A4(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n728), .A2(KEYINPUT105), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT105), .B1(new_n728), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT35), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n613), .B2(new_n568), .ZN(new_n734));
  INV_X1    g533(.A(new_n575), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n614), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n274), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n736), .A2(new_n504), .A3(new_n737), .A4(new_n718), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n729), .B1(new_n738), .B2(new_n726), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT104), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(G8gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n732), .A2(new_n740), .A3(new_n741), .ZN(G1325gat));
  INV_X1    g541(.A(G15gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n567), .A2(new_n564), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n720), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n616), .A2(new_n612), .A3(new_n719), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n743), .B2(new_n746), .ZN(G1326gat));
  NAND2_X1  g546(.A1(new_n720), .A2(new_n529), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT43), .B(G22gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1327gat));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n529), .B1(new_n723), .B2(new_n504), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n598), .A2(new_n601), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT88), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT88), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n598), .B1(new_n595), .B2(new_n501), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n758), .A2(KEYINPUT38), .B1(new_n501), .B2(new_n483), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n412), .A2(new_n757), .A3(new_n759), .A4(new_n573), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n587), .A2(new_n405), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n502), .B1(new_n492), .B2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n495), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n582), .A2(KEYINPUT87), .A3(new_n583), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT87), .B1(new_n582), .B2(new_n583), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n529), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n611), .B1(new_n760), .B2(new_n767), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n570), .A2(new_n575), .B1(new_n752), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n751), .B1(new_n769), .B2(new_n667), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n666), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n717), .B(KEYINPUT107), .Z(new_n773));
  INV_X1    g572(.A(new_n697), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n737), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT108), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(G29gat), .B1(new_n777), .B2(new_n413), .ZN(new_n778));
  INV_X1    g577(.A(new_n717), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n666), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT106), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n736), .A2(new_n737), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n213), .A3(new_n723), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n778), .A2(new_n784), .ZN(G1328gat));
  OAI21_X1  g584(.A(G36gat), .B1(new_n777), .B2(new_n505), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n214), .A3(new_n504), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(G1329gat));
  NAND4_X1  g589(.A1(new_n770), .A2(new_n611), .A3(new_n771), .A4(new_n776), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G43gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n744), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(G43gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n736), .A2(new_n737), .A3(new_n781), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(KEYINPUT47), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n615), .A2(KEYINPUT109), .A3(new_n781), .A4(new_n794), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(G43gat), .B2(new_n791), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n796), .B1(new_n801), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g601(.A1(new_n770), .A2(new_n529), .A3(new_n771), .A4(new_n776), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G50gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n591), .A2(G50gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n736), .A2(new_n737), .A3(new_n781), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n804), .A2(KEYINPUT48), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n615), .A2(new_n808), .A3(new_n781), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n806), .A2(KEYINPUT110), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(G50gat), .B2(new_n803), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n812), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g612(.A1(new_n773), .A2(new_n737), .A3(new_n698), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT111), .Z(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n769), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n723), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n669), .A2(new_n671), .ZN(new_n818));
  XOR2_X1   g617(.A(new_n817), .B(new_n818), .Z(G1332gat));
  AOI21_X1  g618(.A(new_n505), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n822), .A2(new_n826), .A3(new_n824), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1333gat));
  AOI21_X1  g629(.A(new_n676), .B1(new_n816), .B2(new_n611), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n815), .A2(new_n769), .A3(G71gat), .A4(new_n793), .ZN(new_n833));
  OR3_X1    g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n831), .B2(new_n833), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1334gat));
  NAND2_X1  g635(.A1(new_n816), .A2(new_n529), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g637(.A(new_n667), .B1(new_n576), .B2(new_n614), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n737), .A2(new_n697), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT51), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND4_X1   g640(.A1(KEYINPUT51), .A2(new_n736), .A3(new_n666), .A4(new_n840), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT113), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n736), .A2(new_n666), .ZN(new_n846));
  INV_X1    g645(.A(new_n840), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n839), .A2(KEYINPUT51), .A3(new_n840), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n723), .A2(new_n644), .A3(new_n717), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n847), .A2(new_n779), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n772), .A2(new_n723), .A3(new_n853), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n851), .A2(new_n852), .B1(new_n854), .B2(new_n644), .ZN(G1336gat));
  NAND4_X1  g654(.A1(new_n770), .A2(new_n504), .A3(new_n771), .A4(new_n853), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(G92gat), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n773), .A2(G92gat), .A3(new_n505), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n841), .B2(new_n842), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT52), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n857), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n861), .A2(new_n863), .ZN(G1337gat));
  NAND3_X1  g663(.A1(new_n772), .A2(new_n611), .A3(new_n853), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G99gat), .ZN(new_n866));
  OR3_X1    g665(.A1(new_n793), .A2(G99gat), .A3(new_n779), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n866), .B1(new_n851), .B2(new_n867), .ZN(G1338gat));
  NAND4_X1  g667(.A1(new_n770), .A2(new_n529), .A3(new_n771), .A4(new_n853), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G106gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n773), .A2(G106gat), .A3(new_n591), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n841), .B2(new_n842), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n848), .A2(new_n849), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n871), .B(KEYINPUT114), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n875), .A2(new_n876), .B1(new_n869), .B2(G106gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n877), .B2(new_n873), .ZN(G1339gat));
  INV_X1    g677(.A(new_n684), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n648), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n704), .A3(new_n703), .ZN(new_n881));
  INV_X1    g680(.A(new_n705), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n699), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n713), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n882), .A3(new_n707), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n706), .A2(KEYINPUT54), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n884), .B1(new_n883), .B2(new_n699), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n890), .A3(new_n887), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n885), .A2(KEYINPUT55), .A3(new_n713), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n714), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n271), .A2(new_n895), .A3(new_n273), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n252), .B1(new_n248), .B2(new_n250), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n253), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n259), .A2(new_n260), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT116), .B(new_n254), .C1(new_n905), .C2(new_n252), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n262), .A2(new_n264), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n205), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n270), .A3(new_n717), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n666), .B1(new_n901), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n666), .A3(new_n900), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n270), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n774), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n718), .A2(new_n274), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n723), .A2(new_n591), .A3(new_n571), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G113gat), .B1(new_n920), .B2(new_n274), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n917), .A2(new_n568), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n413), .A3(new_n504), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n737), .A2(new_n315), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT117), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n921), .A2(new_n926), .ZN(G1340gat));
  AOI21_X1  g726(.A(G120gat), .B1(new_n923), .B2(new_n717), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n920), .A2(new_n313), .A3(new_n773), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1341gat));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n308), .A3(new_n697), .ZN(new_n931));
  OAI21_X1  g730(.A(G127gat), .B1(new_n920), .B2(new_n774), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1342gat));
  AOI21_X1  g732(.A(new_n310), .B1(new_n919), .B2(new_n666), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT118), .Z(new_n935));
  NAND3_X1  g734(.A1(new_n505), .A2(new_n310), .A3(new_n666), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n922), .A2(new_n413), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1343gat));
  NAND2_X1  g738(.A1(new_n917), .A2(new_n529), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT57), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n591), .B1(new_n915), .B2(new_n916), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT57), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n413), .A2(new_n611), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n505), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n945), .A2(new_n948), .A3(new_n505), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n941), .A2(new_n737), .A3(new_n944), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT121), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n943), .B1(new_n917), .B2(new_n529), .ZN(new_n953));
  AOI211_X1 g752(.A(KEYINPUT57), .B(new_n591), .C1(new_n915), .C2(new_n916), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n737), .A4(new_n950), .ZN(new_n957));
  INV_X1    g756(.A(new_n294), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n945), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n274), .A2(G141gat), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT120), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n960), .A2(new_n504), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(KEYINPUT58), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n951), .A2(new_n958), .ZN(new_n966));
  OAI21_X1  g765(.A(KEYINPUT58), .B1(new_n966), .B2(new_n963), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1344gat));
  NOR2_X1   g767(.A1(new_n960), .A2(new_n504), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n969), .A2(new_n290), .A3(new_n291), .A4(new_n717), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n717), .A3(new_n950), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT59), .B1(new_n290), .B2(new_n291), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT59), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n971), .B2(G148gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n970), .B1(new_n973), .B2(new_n975), .ZN(G1345gat));
  NAND2_X1  g775(.A1(new_n955), .A2(new_n950), .ZN(new_n977));
  OAI21_X1  g776(.A(G155gat), .B1(new_n977), .B2(new_n774), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n278), .A3(new_n697), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1346gat));
  NOR2_X1   g779(.A1(new_n977), .A2(new_n667), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n505), .A2(new_n277), .A3(new_n666), .ZN(new_n982));
  OAI22_X1  g781(.A1(new_n981), .A2(new_n277), .B1(new_n960), .B2(new_n982), .ZN(G1347gat));
  NAND2_X1  g782(.A1(new_n413), .A2(new_n504), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n922), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT122), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n421), .A3(new_n737), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n737), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G169gat), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n989), .A2(KEYINPUT123), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n987), .B1(new_n990), .B2(new_n991), .ZN(G1348gat));
  NOR4_X1   g791(.A1(new_n922), .A2(new_n422), .A3(new_n773), .A4(new_n984), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT124), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n986), .A2(new_n717), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(new_n422), .ZN(G1349gat));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n997));
  AOI21_X1  g796(.A(G183gat), .B1(new_n985), .B2(new_n697), .ZN(new_n998));
  NOR4_X1   g797(.A1(new_n922), .A2(new_n442), .A3(new_n774), .A4(new_n984), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n998), .A2(new_n999), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  OAI211_X1 g803(.A(KEYINPUT126), .B(new_n997), .C1(new_n998), .C2(new_n999), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(G1350gat));
  NAND3_X1  g805(.A1(new_n986), .A2(new_n416), .A3(new_n666), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n985), .A2(new_n666), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1008), .A2(G190gat), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n1009), .A2(KEYINPUT61), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1009), .A2(KEYINPUT61), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(G1351gat));
  NOR2_X1   g811(.A1(new_n611), .A2(new_n505), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1014), .A2(new_n1015), .A3(new_n591), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT127), .B1(new_n1013), .B2(new_n529), .ZN(new_n1017));
  NOR3_X1   g816(.A1(new_n1016), .A2(new_n723), .A3(new_n1017), .ZN(new_n1018));
  AND2_X1   g817(.A1(new_n1018), .A2(new_n917), .ZN(new_n1019));
  AOI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n737), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1014), .A2(new_n723), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n955), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n737), .A2(G197gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(G1352gat));
  NOR2_X1   g824(.A1(new_n779), .A2(G204gat), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g826(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  OAI21_X1  g827(.A(G204gat), .B1(new_n1022), .B2(new_n773), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(G1353gat));
  INV_X1    g830(.A(G211gat), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1019), .A2(new_n1032), .A3(new_n697), .ZN(new_n1033));
  NAND3_X1  g832(.A1(new_n955), .A2(new_n697), .A3(new_n1021), .ZN(new_n1034));
  AND3_X1   g833(.A1(new_n1034), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1035));
  AOI21_X1  g834(.A(KEYINPUT63), .B1(new_n1034), .B2(G211gat), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(G1354gat));
  OAI21_X1  g836(.A(G218gat), .B1(new_n1022), .B2(new_n667), .ZN(new_n1038));
  INV_X1    g837(.A(G218gat), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n1019), .A2(new_n1039), .A3(new_n666), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1038), .A2(new_n1040), .ZN(G1355gat));
endmodule


