

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n753), .A2(n752), .ZN(n724) );
  INV_X1 U555 ( .A(n724), .ZN(n697) );
  XNOR2_X1 U556 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U557 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n686) );
  XNOR2_X1 U558 ( .A(n687), .B(n686), .ZN(n689) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n690) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n719) );
  XNOR2_X1 U561 ( .A(n719), .B(KEYINPUT94), .ZN(n720) );
  XNOR2_X1 U562 ( .A(n721), .B(n720), .ZN(n722) );
  OR2_X1 U563 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U564 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n523) );
  OR2_X1 U565 ( .A1(n804), .A2(n803), .ZN(n819) );
  AND2_X1 U566 ( .A1(n522), .A2(G2104), .ZN(n894) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n528), .Z(n895) );
  AND2_X1 U568 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U569 ( .A1(G651), .A2(n631), .ZN(n635) );
  NOR2_X1 U570 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U571 ( .A(G2105), .ZN(n522) );
  NAND2_X1 U572 ( .A1(G101), .A2(n894), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n522), .ZN(n890) );
  NAND2_X1 U574 ( .A1(n890), .A2(G125), .ZN(n525) );
  NAND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U576 ( .A(KEYINPUT66), .B(n527), .ZN(n532) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n895), .A2(G137), .ZN(n530) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U580 ( .A1(n891), .A2(G113), .ZN(n529) );
  NAND2_X1 U581 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U583 ( .A1(G85), .A2(n638), .ZN(n534) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  INV_X1 U585 ( .A(G651), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n631), .A2(n535), .ZN(n639) );
  NAND2_X1 U587 ( .A1(G72), .A2(n639), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n536), .Z(n634) );
  NAND2_X1 U591 ( .A1(G60), .A2(n634), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G47), .A2(n635), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  OR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G290) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U596 ( .A(G57), .ZN(G237) );
  NAND2_X1 U597 ( .A1(n638), .A2(G89), .ZN(n541) );
  XNOR2_X1 U598 ( .A(KEYINPUT4), .B(n541), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n639), .A2(G76), .ZN(n542) );
  XOR2_X1 U600 ( .A(KEYINPUT73), .B(n542), .Z(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U602 ( .A(n545), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n634), .A2(G63), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT74), .ZN(n548) );
  NAND2_X1 U605 ( .A1(G51), .A2(n635), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U611 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n554) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n554), .B(n553), .ZN(G223) );
  XOR2_X1 U614 ( .A(G223), .B(KEYINPUT70), .Z(n824) );
  NAND2_X1 U615 ( .A1(n824), .A2(G567), .ZN(n555) );
  XOR2_X1 U616 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  NAND2_X1 U617 ( .A1(n634), .A2(G56), .ZN(n556) );
  XNOR2_X1 U618 ( .A(n556), .B(KEYINPUT14), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G43), .A2(n635), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n638), .A2(G81), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT12), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G68), .A2(n639), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U625 ( .A(KEYINPUT13), .B(n562), .ZN(n563) );
  XNOR2_X1 U626 ( .A(KEYINPUT71), .B(n563), .ZN(n564) );
  NOR2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n1010) );
  NAND2_X1 U628 ( .A1(n1010), .A2(G860), .ZN(G153) );
  NAND2_X1 U629 ( .A1(G90), .A2(n638), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G77), .A2(n639), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n573) );
  NAND2_X1 U634 ( .A1(G64), .A2(n634), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G52), .A2(n635), .ZN(n570) );
  AND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G92), .A2(n638), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G79), .A2(n639), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G66), .A2(n634), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G54), .A2(n635), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n1004) );
  NOR2_X1 U647 ( .A1(n1004), .A2(G868), .ZN(n583) );
  INV_X1 U648 ( .A(G868), .ZN(n645) );
  NOR2_X1 U649 ( .A1(n645), .A2(G301), .ZN(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G91), .A2(n638), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G78), .A2(n639), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n634), .A2(G65), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT68), .B(n586), .Z(n587) );
  NOR2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n635), .A2(G53), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n645), .ZN(n592) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U662 ( .A(G860), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n593), .A2(G559), .ZN(n594) );
  INV_X1 U664 ( .A(n1004), .ZN(n610) );
  NAND2_X1 U665 ( .A1(n594), .A2(n610), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U667 ( .A1(n1010), .A2(n645), .ZN(n596) );
  XNOR2_X1 U668 ( .A(KEYINPUT75), .B(n596), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G868), .A2(n610), .ZN(n597) );
  NOR2_X1 U670 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G111), .A2(n891), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G135), .A2(n895), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U675 ( .A1(n890), .A2(G123), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n894), .A2(G99), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n974) );
  XOR2_X1 U680 ( .A(G2096), .B(KEYINPUT76), .Z(n607) );
  XNOR2_X1 U681 ( .A(n974), .B(n607), .ZN(n609) );
  INV_X1 U682 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U684 ( .A1(n610), .A2(G559), .ZN(n611) );
  XOR2_X1 U685 ( .A(n1010), .B(n611), .Z(n653) );
  NOR2_X1 U686 ( .A1(n653), .A2(G860), .ZN(n618) );
  NAND2_X1 U687 ( .A1(G67), .A2(n634), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G55), .A2(n635), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U690 ( .A1(G93), .A2(n638), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G80), .A2(n639), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n649) );
  XNOR2_X1 U694 ( .A(n618), .B(n649), .ZN(G145) );
  NAND2_X1 U695 ( .A1(G86), .A2(n638), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G61), .A2(n634), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U698 ( .A(KEYINPUT78), .B(n621), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n639), .A2(G73), .ZN(n622) );
  XOR2_X1 U700 ( .A(KEYINPUT2), .B(n622), .Z(n623) );
  NOR2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n635), .A2(G48), .ZN(n625) );
  NAND2_X1 U703 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U704 ( .A1(G49), .A2(n635), .ZN(n628) );
  NAND2_X1 U705 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U707 ( .A1(n634), .A2(n629), .ZN(n630) );
  XOR2_X1 U708 ( .A(KEYINPUT77), .B(n630), .Z(n633) );
  NAND2_X1 U709 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G62), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G50), .A2(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G88), .A2(n638), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G75), .A2(n639), .ZN(n640) );
  NAND2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(KEYINPUT79), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(n645), .A2(n649), .ZN(n656) );
  XNOR2_X1 U721 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n647) );
  XNOR2_X1 U722 ( .A(G290), .B(G166), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(G299), .ZN(n651) );
  XNOR2_X1 U726 ( .A(G288), .B(n651), .ZN(n652) );
  XNOR2_X1 U727 ( .A(G305), .B(n652), .ZN(n846) );
  XNOR2_X1 U728 ( .A(n846), .B(n653), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n654), .A2(G868), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n657), .B(KEYINPUT81), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n661), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U738 ( .A1(G69), .A2(G120), .ZN(n662) );
  NOR2_X1 U739 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G108), .A2(n663), .ZN(n830) );
  NAND2_X1 U741 ( .A1(G567), .A2(n830), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT83), .B(n664), .Z(n670) );
  NAND2_X1 U743 ( .A1(G132), .A2(G82), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n665), .B(KEYINPUT22), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT82), .ZN(n667) );
  NOR2_X1 U746 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G96), .A2(n668), .ZN(n831) );
  NAND2_X1 U748 ( .A1(G2106), .A2(n831), .ZN(n669) );
  NAND2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U750 ( .A(KEYINPUT84), .B(n671), .Z(G319) );
  INV_X1 U751 ( .A(G319), .ZN(n913) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n672) );
  NOR2_X1 U753 ( .A1(n913), .A2(n672), .ZN(n829) );
  NAND2_X1 U754 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(n895), .A2(G138), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G102), .A2(n894), .ZN(n673) );
  XOR2_X1 U757 ( .A(KEYINPUT85), .B(n673), .Z(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n679) );
  NAND2_X1 U759 ( .A1(G126), .A2(n890), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G114), .A2(n891), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U762 ( .A1(n679), .A2(n678), .ZN(G164) );
  INV_X1 U763 ( .A(G301), .ZN(G171) );
  NOR2_X1 U764 ( .A1(G1976), .A2(G288), .ZN(n742) );
  INV_X1 U765 ( .A(n742), .ZN(n1016) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n753) );
  NAND2_X1 U767 ( .A1(G40), .A2(G160), .ZN(n681) );
  INV_X1 U768 ( .A(KEYINPUT86), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n681), .B(n680), .ZN(n752) );
  NAND2_X1 U770 ( .A1(G8), .A2(n724), .ZN(n797) );
  OR2_X1 U771 ( .A1(n1016), .A2(n797), .ZN(n682) );
  AND2_X1 U772 ( .A1(n682), .A2(KEYINPUT33), .ZN(n750) );
  XOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .Z(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT91), .B(n683), .ZN(n955) );
  NOR2_X1 U775 ( .A1(n724), .A2(n955), .ZN(n685) );
  INV_X1 U776 ( .A(G1961), .ZN(n940) );
  NOR2_X1 U777 ( .A1(n697), .A2(n940), .ZN(n684) );
  NOR2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n713), .A2(G171), .ZN(n712) );
  NAND2_X1 U780 ( .A1(G2072), .A2(n697), .ZN(n687) );
  AND2_X1 U781 ( .A1(G1956), .A2(n724), .ZN(n688) );
  NOR2_X1 U782 ( .A1(n689), .A2(n688), .ZN(n692) );
  INV_X1 U783 ( .A(G299), .ZN(n1005) );
  NOR2_X1 U784 ( .A1(n692), .A2(n1005), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n691), .B(n690), .ZN(n708) );
  NAND2_X1 U786 ( .A1(n692), .A2(n1005), .ZN(n706) );
  NAND2_X1 U787 ( .A1(G1348), .A2(n724), .ZN(n694) );
  NAND2_X1 U788 ( .A1(G2067), .A2(n697), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n1004), .A2(n702), .ZN(n696) );
  NAND2_X1 U791 ( .A1(G1341), .A2(n724), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n697), .A2(G1996), .ZN(n698) );
  XNOR2_X1 U794 ( .A(n698), .B(KEYINPUT26), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n699), .A2(n1010), .ZN(n700) );
  NOR2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n1004), .A2(n702), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n710) );
  XNOR2_X1 U801 ( .A(KEYINPUT93), .B(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U802 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n723) );
  NOR2_X1 U804 ( .A1(G171), .A2(n713), .ZN(n718) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n797), .ZN(n736) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n724), .ZN(n733) );
  NOR2_X1 U807 ( .A1(n736), .A2(n733), .ZN(n714) );
  NAND2_X1 U808 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U810 ( .A1(G168), .A2(n716), .ZN(n717) );
  NOR2_X1 U811 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n734) );
  NAND2_X1 U813 ( .A1(n734), .A2(G286), .ZN(n731) );
  INV_X1 U814 ( .A(G8), .ZN(n729) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n797), .ZN(n726) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n727), .A2(G303), .ZN(n728) );
  OR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT32), .ZN(n794) );
  NAND2_X1 U822 ( .A1(G8), .A2(n733), .ZN(n738) );
  INV_X1 U823 ( .A(n734), .ZN(n735) );
  NOR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n793) );
  NAND2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  INV_X1 U827 ( .A(n1015), .ZN(n739) );
  OR2_X1 U828 ( .A1(n739), .A2(n797), .ZN(n744) );
  INV_X1 U829 ( .A(n744), .ZN(n740) );
  AND2_X1 U830 ( .A1(n793), .A2(n740), .ZN(n741) );
  NAND2_X1 U831 ( .A1(n794), .A2(n741), .ZN(n746) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n1012) );
  NOR2_X1 U833 ( .A1(n742), .A2(n1012), .ZN(n743) );
  OR2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U836 ( .A(n747), .B(KEYINPUT64), .Z(n748) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n748), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U839 ( .A(KEYINPUT95), .B(n751), .ZN(n786) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n1024) );
  INV_X1 U841 ( .A(n752), .ZN(n754) );
  NOR2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n816) );
  NAND2_X1 U843 ( .A1(G104), .A2(n894), .ZN(n756) );
  NAND2_X1 U844 ( .A1(G140), .A2(n895), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U846 ( .A(KEYINPUT34), .B(n757), .ZN(n762) );
  NAND2_X1 U847 ( .A1(G128), .A2(n890), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G116), .A2(n891), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U850 ( .A(KEYINPUT35), .B(n760), .Z(n761) );
  NOR2_X1 U851 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U852 ( .A(KEYINPUT36), .B(n763), .ZN(n904) );
  XNOR2_X1 U853 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U854 ( .A1(n904), .A2(n805), .ZN(n978) );
  NAND2_X1 U855 ( .A1(n816), .A2(n978), .ZN(n813) );
  XNOR2_X1 U856 ( .A(n816), .B(KEYINPUT88), .ZN(n780) );
  NAND2_X1 U857 ( .A1(G107), .A2(n891), .ZN(n765) );
  NAND2_X1 U858 ( .A1(G131), .A2(n895), .ZN(n764) );
  NAND2_X1 U859 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G119), .A2(n890), .ZN(n767) );
  NAND2_X1 U861 ( .A1(G95), .A2(n894), .ZN(n766) );
  NAND2_X1 U862 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n887) );
  NAND2_X1 U864 ( .A1(G1991), .A2(n887), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G117), .A2(n891), .ZN(n771) );
  NAND2_X1 U866 ( .A1(G141), .A2(n895), .ZN(n770) );
  NAND2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U868 ( .A1(G105), .A2(n894), .ZN(n772) );
  XNOR2_X1 U869 ( .A(n772), .B(KEYINPUT38), .ZN(n773) );
  XNOR2_X1 U870 ( .A(n773), .B(KEYINPUT87), .ZN(n774) );
  NOR2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n890), .A2(G129), .ZN(n776) );
  NAND2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n907) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n907), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n970) );
  NAND2_X1 U876 ( .A1(n780), .A2(n970), .ZN(n781) );
  XNOR2_X1 U877 ( .A(KEYINPUT89), .B(n781), .ZN(n809) );
  INV_X1 U878 ( .A(n809), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n813), .A2(n782), .ZN(n783) );
  XOR2_X1 U880 ( .A(n783), .B(KEYINPUT90), .Z(n788) );
  AND2_X1 U881 ( .A1(n1024), .A2(n788), .ZN(n784) );
  XNOR2_X1 U882 ( .A(G1986), .B(G290), .ZN(n1011) );
  NAND2_X1 U883 ( .A1(n1011), .A2(n816), .ZN(n787) );
  AND2_X1 U884 ( .A1(n784), .A2(n787), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n821) );
  INV_X1 U886 ( .A(n787), .ZN(n804) );
  INV_X1 U887 ( .A(n788), .ZN(n802) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U889 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  OR2_X1 U890 ( .A1(n797), .A2(n790), .ZN(n800) );
  NOR2_X1 U891 ( .A1(G2090), .A2(G303), .ZN(n791) );
  XNOR2_X1 U892 ( .A(KEYINPUT96), .B(n791), .ZN(n792) );
  NAND2_X1 U893 ( .A1(n792), .A2(G8), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n904), .A2(n805), .ZN(n969) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n907), .ZN(n981) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n887), .ZN(n806) );
  XOR2_X1 U902 ( .A(KEYINPUT97), .B(n806), .Z(n973) );
  NOR2_X1 U903 ( .A1(n807), .A2(n973), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n981), .A2(n810), .ZN(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT98), .B(n811), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n969), .A2(n815), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n823) );
  XOR2_X1 U912 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n822) );
  XNOR2_X1 U913 ( .A(n823), .B(n822), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n824), .ZN(G217) );
  INV_X1 U915 ( .A(G661), .ZN(n826) );
  NAND2_X1 U916 ( .A1(G2), .A2(G15), .ZN(n825) );
  NOR2_X1 U917 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U918 ( .A(KEYINPUT102), .B(n827), .Z(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G82), .ZN(G220) );
  INV_X1 U925 ( .A(G69), .ZN(G235) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U927 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U928 ( .A(KEYINPUT100), .B(G2454), .ZN(n840) );
  XNOR2_X1 U929 ( .A(G2430), .B(G2435), .ZN(n838) );
  XOR2_X1 U930 ( .A(G2451), .B(G2427), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2438), .B(G2446), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n834), .B(G2443), .Z(n836) );
  XNOR2_X1 U934 ( .A(G1348), .B(G1341), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n841), .A2(G14), .ZN(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT101), .B(n842), .ZN(G401) );
  XOR2_X1 U940 ( .A(G286), .B(n1004), .Z(n844) );
  XNOR2_X1 U941 ( .A(G171), .B(n1010), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(n846), .B(n845), .Z(n847) );
  NOR2_X1 U944 ( .A1(G37), .A2(n847), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT111), .B(n848), .Z(G397) );
  XOR2_X1 U946 ( .A(G2100), .B(KEYINPUT103), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT104), .B(KEYINPUT43), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(KEYINPUT42), .B(G2090), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2678), .B(G2096), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U955 ( .A(G2084), .B(G2078), .Z(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1971), .B(G1956), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1991), .B(G1961), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U960 ( .A(G1976), .B(G1981), .Z(n862) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1966), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U963 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U964 ( .A(KEYINPUT105), .B(G2474), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n868) );
  XOR2_X1 U966 ( .A(G1996), .B(KEYINPUT41), .Z(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U968 ( .A1(G112), .A2(n891), .ZN(n869) );
  XNOR2_X1 U969 ( .A(n869), .B(KEYINPUT106), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G124), .A2(n890), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n870), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G100), .A2(n894), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G136), .A2(n895), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(G162) );
  XOR2_X1 U977 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  XNOR2_X1 U978 ( .A(KEYINPUT110), .B(KEYINPUT109), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n889) );
  NAND2_X1 U980 ( .A1(G103), .A2(n894), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G139), .A2(n895), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G127), .A2(n890), .ZN(n882) );
  NAND2_X1 U984 ( .A1(G115), .A2(n891), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n987) );
  XOR2_X1 U988 ( .A(G160), .B(n987), .Z(n886) );
  XNOR2_X1 U989 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U990 ( .A(n889), .B(n888), .ZN(n906) );
  NAND2_X1 U991 ( .A1(G130), .A2(n890), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G118), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n902) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n900) );
  NAND2_X1 U995 ( .A1(n894), .A2(G106), .ZN(n898) );
  NAND2_X1 U996 ( .A1(n895), .A2(G142), .ZN(n896) );
  XOR2_X1 U997 ( .A(KEYINPUT107), .B(n896), .Z(n897) );
  NAND2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U999 ( .A(n900), .B(n899), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(G162), .B(n907), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n908), .B(n974), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(G164), .B(n909), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n912), .ZN(G395) );
  NOR2_X1 U1008 ( .A1(n913), .A2(G401), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G397), .A2(n915), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n918), .A2(G395), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1015 ( .A(G308), .ZN(G225) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1018 ( .A(G1986), .B(G24), .Z(n923) );
  XNOR2_X1 U1019 ( .A(G1971), .B(G22), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G23), .B(G1976), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n925), .B(n924), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(G1348), .B(KEYINPUT59), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(G4), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G20), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(G19), .B(G1341), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1031 ( .A(KEYINPUT125), .B(G1981), .Z(n931) );
  XNOR2_X1 U1032 ( .A(G6), .B(n931), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1034 ( .A(n934), .B(KEYINPUT60), .Z(n935) );
  XNOR2_X1 U1035 ( .A(KEYINPUT126), .B(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G21), .B(G1966), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1039 ( .A(G5), .B(n940), .Z(n941) );
  XNOR2_X1 U1040 ( .A(KEYINPUT124), .B(n941), .ZN(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT61), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G16), .B(KEYINPUT123), .ZN(n945) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(G11), .A2(n947), .ZN(n1001) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1048 ( .A1(n949), .A2(n948), .ZN(n954) );
  XOR2_X1 U1049 ( .A(G1991), .B(G25), .Z(n950) );
  NAND2_X1 U1050 ( .A1(n950), .A2(G28), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1054 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n958), .B(KEYINPUT117), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(KEYINPUT53), .ZN(n962) );
  XOR2_X1 U1058 ( .A(G2084), .B(G34), .Z(n960) );
  XNOR2_X1 U1059 ( .A(KEYINPUT54), .B(n960), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(n965), .B(KEYINPUT118), .ZN(n966) );
  XOR2_X1 U1064 ( .A(KEYINPUT55), .B(KEYINPUT116), .Z(n995) );
  XNOR2_X1 U1065 ( .A(n966), .B(n995), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(G29), .A2(n967), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(n968), .B(KEYINPUT119), .ZN(n999) );
  INV_X1 U1068 ( .A(n969), .ZN(n971) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n986) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1073 ( .A(KEYINPUT113), .B(n976), .Z(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1075 ( .A(KEYINPUT114), .B(n979), .Z(n984) );
  XOR2_X1 U1076 ( .A(G2090), .B(G162), .Z(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT51), .B(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G2072), .B(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(G164), .B(G2078), .ZN(n988) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1084 ( .A(KEYINPUT115), .B(n990), .Z(n991) );
  XNOR2_X1 U1085 ( .A(KEYINPUT50), .B(n991), .ZN(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(G29), .A2(n997), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1032) );
  XNOR2_X1 U1092 ( .A(G171), .B(G1961), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(G1971), .A2(G303), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(n1004), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1096 ( .A(n1005), .B(G1956), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1021) );
  XNOR2_X1 U1099 ( .A(n1010), .B(G1341), .ZN(n1014) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1019) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT121), .B(n1017), .Z(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1027) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G168), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT120), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1025), .Z(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT122), .B(n1028), .Z(n1030) );
  XNOR2_X1 U1112 ( .A(G16), .B(KEYINPUT56), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

