

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U554 ( .A(KEYINPUT32), .B(n739), .ZN(n816) );
  XNOR2_X1 U555 ( .A(n710), .B(n709), .ZN(n716) );
  NAND2_X1 U556 ( .A1(n561), .A2(n521), .ZN(n562) );
  AND2_X1 U557 ( .A1(n560), .A2(n559), .ZN(n521) );
  NOR2_X1 U558 ( .A1(n826), .A2(n806), .ZN(n522) );
  AND2_X1 U559 ( .A1(G137), .A2(n882), .ZN(n523) );
  NOR2_X1 U560 ( .A1(n812), .A2(n752), .ZN(n524) );
  AND2_X1 U561 ( .A1(n754), .A2(n753), .ZN(n525) );
  XOR2_X1 U562 ( .A(KEYINPUT95), .B(n721), .Z(n526) );
  NOR2_X1 U563 ( .A1(n993), .A2(n694), .ZN(n697) );
  INV_X1 U564 ( .A(KEYINPUT94), .ZN(n695) );
  XNOR2_X1 U565 ( .A(n696), .B(n695), .ZN(n703) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n709) );
  XNOR2_X1 U567 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U568 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U569 ( .A1(G1966), .A2(n812), .ZN(n743) );
  NAND2_X1 U570 ( .A1(n777), .A2(n778), .ZN(n729) );
  NOR2_X1 U571 ( .A1(n524), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  NOR2_X2 U573 ( .A1(G2105), .A2(n530), .ZN(n880) );
  NOR2_X1 U574 ( .A1(G651), .A2(n640), .ZN(n645) );
  NOR2_X1 U575 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U576 ( .A1(G102), .A2(n880), .ZN(n529) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n527), .Z(n882) );
  NAND2_X1 U578 ( .A1(G138), .A2(n882), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n538) );
  INV_X1 U580 ( .A(KEYINPUT83), .ZN(n536) );
  INV_X1 U581 ( .A(G2104), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n530), .A2(G2105), .ZN(n531) );
  XNOR2_X2 U583 ( .A(n531), .B(KEYINPUT65), .ZN(n889) );
  NAND2_X1 U584 ( .A1(n889), .A2(G126), .ZN(n532) );
  XNOR2_X1 U585 ( .A(n532), .B(KEYINPUT82), .ZN(n534) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U587 ( .A1(G114), .A2(n886), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U589 ( .A(n536), .B(n535), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U591 ( .A1(n647), .A2(G89), .ZN(n539) );
  XNOR2_X1 U592 ( .A(n539), .B(KEYINPUT4), .ZN(n541) );
  XOR2_X1 U593 ( .A(G543), .B(KEYINPUT0), .Z(n640) );
  INV_X1 U594 ( .A(G651), .ZN(n543) );
  NOR2_X1 U595 ( .A1(n640), .A2(n543), .ZN(n648) );
  NAND2_X1 U596 ( .A1(G76), .A2(n648), .ZN(n540) );
  NAND2_X1 U597 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U598 ( .A(n542), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G51), .A2(n645), .ZN(n546) );
  NOR2_X1 U600 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n544), .Z(n651) );
  NAND2_X1 U602 ( .A1(G63), .A2(n651), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G85), .A2(n647), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G60), .A2(n651), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G72), .A2(n648), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G47), .A2(n645), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G290) );
  NAND2_X1 U615 ( .A1(G101), .A2(n880), .ZN(n557) );
  XOR2_X1 U616 ( .A(KEYINPUT23), .B(n557), .Z(n558) );
  XNOR2_X1 U617 ( .A(n558), .B(KEYINPUT66), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G113), .A2(n886), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G125), .A2(n889), .ZN(n559) );
  NOR2_X1 U620 ( .A1(n562), .A2(n523), .ZN(n563) );
  XNOR2_X1 U621 ( .A(KEYINPUT64), .B(n563), .ZN(G160) );
  INV_X1 U622 ( .A(G57), .ZN(G237) );
  NAND2_X1 U623 ( .A1(G94), .A2(G452), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(n564), .Z(G173) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U627 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n567) );
  INV_X1 U628 ( .A(G223), .ZN(n833) );
  NAND2_X1 U629 ( .A1(G567), .A2(n833), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n567), .B(n566), .ZN(G234) );
  NAND2_X1 U631 ( .A1(n651), .A2(G56), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n568), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n647), .A2(G81), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G68), .A2(n648), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(n572), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(n575), .B(KEYINPUT71), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n645), .A2(G43), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n993) );
  INV_X1 U642 ( .A(G860), .ZN(n605) );
  OR2_X1 U643 ( .A1(n993), .A2(n605), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G52), .A2(n645), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT67), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G90), .A2(n647), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G77), .A2(n648), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U649 ( .A(KEYINPUT9), .B(n581), .Z(n582) );
  NOR2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n651), .A2(G64), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G92), .A2(n647), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G66), .A2(n651), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G79), .A2(n648), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G54), .A2(n645), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n592), .Z(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT72), .B(n593), .ZN(n980) );
  INV_X1 U662 ( .A(G868), .ZN(n665) );
  AND2_X1 U663 ( .A1(n980), .A2(n665), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n665), .A2(G301), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G91), .A2(n647), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G65), .A2(n651), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G78), .A2(n648), .ZN(n598) );
  XNOR2_X1 U670 ( .A(KEYINPUT69), .B(n598), .ZN(n599) );
  NOR2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n645), .A2(G53), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G299) );
  NOR2_X1 U674 ( .A1(G286), .A2(n665), .ZN(n604) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n606), .A2(n980), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n993), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT73), .B(n608), .Z(n611) );
  NAND2_X1 U682 ( .A1(G868), .A2(n980), .ZN(n609) );
  NOR2_X1 U683 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G99), .A2(n880), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G111), .A2(n886), .ZN(n612) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n889), .A2(G123), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT18), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G135), .A2(n882), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n926) );
  XNOR2_X1 U693 ( .A(n926), .B(G2096), .ZN(n620) );
  INV_X1 U694 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U695 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G559), .A2(n980), .ZN(n663) );
  XNOR2_X1 U697 ( .A(n993), .B(n663), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n621), .A2(G860), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G55), .A2(n645), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G67), .A2(n651), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G93), .A2(n647), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G80), .A2(n648), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n666) );
  XOR2_X1 U706 ( .A(n628), .B(n666), .Z(G145) );
  NAND2_X1 U707 ( .A1(G86), .A2(n647), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G61), .A2(n651), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n648), .A2(G73), .ZN(n631) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n631), .Z(n632) );
  NOR2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n645), .A2(G48), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(G305) );
  NAND2_X1 U715 ( .A1(G651), .A2(G74), .ZN(n636) );
  XNOR2_X1 U716 ( .A(n636), .B(KEYINPUT74), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G49), .A2(n645), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n639), .B(KEYINPUT75), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G87), .A2(n640), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U722 ( .A1(n651), .A2(n643), .ZN(n644) );
  XOR2_X1 U723 ( .A(KEYINPUT76), .B(n644), .Z(G288) );
  NAND2_X1 U724 ( .A1(G50), .A2(n645), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n646), .B(KEYINPUT78), .ZN(n656) );
  NAND2_X1 U726 ( .A1(G88), .A2(n647), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G75), .A2(n648), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U729 ( .A1(G62), .A2(n651), .ZN(n652) );
  XNOR2_X1 U730 ( .A(KEYINPUT77), .B(n652), .ZN(n653) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U732 ( .A1(n656), .A2(n655), .ZN(G303) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(n666), .ZN(n657) );
  XNOR2_X1 U734 ( .A(G290), .B(n657), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n658), .B(G305), .ZN(n661) );
  INV_X1 U736 ( .A(G299), .ZN(n979) );
  XNOR2_X1 U737 ( .A(n979), .B(G288), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n659), .B(G303), .ZN(n660) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(n993), .ZN(n901) );
  XNOR2_X1 U741 ( .A(n901), .B(n663), .ZN(n664) );
  NOR2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U743 ( .A1(G868), .A2(n666), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U749 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XOR2_X1 U750 ( .A(KEYINPUT79), .B(G44), .Z(n673) );
  XNOR2_X1 U751 ( .A(KEYINPUT3), .B(n673), .ZN(G218) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G108), .A2(n675), .ZN(n921) );
  NAND2_X1 U755 ( .A1(G567), .A2(n921), .ZN(n682) );
  NAND2_X1 U756 ( .A1(G132), .A2(G82), .ZN(n676) );
  XNOR2_X1 U757 ( .A(n676), .B(KEYINPUT80), .ZN(n677) );
  XNOR2_X1 U758 ( .A(n677), .B(KEYINPUT22), .ZN(n678) );
  NOR2_X1 U759 ( .A1(G218), .A2(n678), .ZN(n679) );
  XOR2_X1 U760 ( .A(KEYINPUT81), .B(n679), .Z(n680) );
  NAND2_X1 U761 ( .A1(G96), .A2(n680), .ZN(n920) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n920), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n682), .A2(n681), .ZN(n838) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U765 ( .A1(n838), .A2(n683), .ZN(n836) );
  NAND2_X1 U766 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U767 ( .A(G303), .ZN(G166) );
  INV_X1 U768 ( .A(G301), .ZN(G171) );
  AND2_X1 U769 ( .A1(G40), .A2(G160), .ZN(n777) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n778) );
  INV_X2 U771 ( .A(n729), .ZN(n712) );
  NAND2_X1 U772 ( .A1(n712), .A2(G2072), .ZN(n685) );
  XNOR2_X1 U773 ( .A(n685), .B(KEYINPUT27), .ZN(n687) );
  AND2_X1 U774 ( .A1(G1956), .A2(n729), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n704) );
  NOR2_X1 U776 ( .A1(n704), .A2(n979), .ZN(n689) );
  XOR2_X1 U777 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n688) );
  XNOR2_X1 U778 ( .A(n689), .B(n688), .ZN(n708) );
  AND2_X1 U779 ( .A1(n712), .A2(G1996), .ZN(n691) );
  XNOR2_X1 U780 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n729), .A2(G1341), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n697), .A2(n980), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n980), .ZN(n701) );
  NOR2_X1 U786 ( .A1(G2067), .A2(n729), .ZN(n699) );
  NOR2_X1 U787 ( .A1(n712), .A2(G1348), .ZN(n698) );
  NOR2_X1 U788 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U790 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n704), .A2(n979), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U794 ( .A1(n712), .A2(G1961), .ZN(n711) );
  XNOR2_X1 U795 ( .A(n711), .B(KEYINPUT91), .ZN(n714) );
  XNOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U797 ( .A1(n712), .A2(n955), .ZN(n713) );
  NAND2_X1 U798 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U799 ( .A1(n717), .A2(G171), .ZN(n715) );
  NAND2_X1 U800 ( .A1(n716), .A2(n715), .ZN(n728) );
  NOR2_X1 U801 ( .A1(G171), .A2(n717), .ZN(n722) );
  NAND2_X1 U802 ( .A1(G8), .A2(n729), .ZN(n812) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n729), .ZN(n740) );
  NOR2_X1 U804 ( .A1(n743), .A2(n740), .ZN(n718) );
  NAND2_X1 U805 ( .A1(G8), .A2(n718), .ZN(n719) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n719), .ZN(n720) );
  NOR2_X1 U807 ( .A1(G168), .A2(n720), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n526), .ZN(n726) );
  XOR2_X1 U809 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n724) );
  INV_X1 U810 ( .A(KEYINPUT31), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n728), .A2(n727), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n741), .A2(G286), .ZN(n735) );
  NOR2_X1 U813 ( .A1(G2090), .A2(n729), .ZN(n730) );
  XNOR2_X1 U814 ( .A(n730), .B(KEYINPUT98), .ZN(n732) );
  NOR2_X1 U815 ( .A1(n812), .A2(G1971), .ZN(n731) );
  NOR2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U817 ( .A1(n733), .A2(G303), .ZN(n734) );
  NAND2_X1 U818 ( .A1(n735), .A2(n734), .ZN(n737) );
  INV_X1 U819 ( .A(KEYINPUT99), .ZN(n736) );
  XNOR2_X1 U820 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n738), .A2(G8), .ZN(n739) );
  NAND2_X1 U822 ( .A1(G8), .A2(n740), .ZN(n745) );
  INV_X1 U823 ( .A(n741), .ZN(n742) );
  NOR2_X1 U824 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U825 ( .A1(n745), .A2(n744), .ZN(n814) );
  NAND2_X1 U826 ( .A1(G288), .A2(G1976), .ZN(n973) );
  AND2_X1 U827 ( .A1(n814), .A2(n973), .ZN(n746) );
  NAND2_X1 U828 ( .A1(n816), .A2(n746), .ZN(n754) );
  INV_X1 U829 ( .A(n973), .ZN(n751) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n747) );
  XNOR2_X1 U831 ( .A(KEYINPUT101), .B(n747), .ZN(n749) );
  NOR2_X1 U832 ( .A1(G288), .A2(G1976), .ZN(n748) );
  XOR2_X1 U833 ( .A(KEYINPUT100), .B(n748), .Z(n972) );
  AND2_X1 U834 ( .A1(n749), .A2(n972), .ZN(n750) );
  OR2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n752) );
  INV_X1 U836 ( .A(KEYINPUT102), .ZN(n755) );
  XNOR2_X1 U837 ( .A(n525), .B(n755), .ZN(n809) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n976) );
  NOR2_X1 U839 ( .A1(n812), .A2(n972), .ZN(n756) );
  NAND2_X1 U840 ( .A1(KEYINPUT33), .A2(n756), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n976), .A2(n757), .ZN(n807) );
  NAND2_X1 U842 ( .A1(G117), .A2(n886), .ZN(n759) );
  NAND2_X1 U843 ( .A1(G129), .A2(n889), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U845 ( .A1(G105), .A2(n880), .ZN(n760) );
  XNOR2_X1 U846 ( .A(n760), .B(KEYINPUT38), .ZN(n761) );
  XNOR2_X1 U847 ( .A(n761), .B(KEYINPUT89), .ZN(n762) );
  NOR2_X1 U848 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n882), .A2(G141), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(n875) );
  NOR2_X1 U851 ( .A1(G1996), .A2(n875), .ZN(n924) );
  NAND2_X1 U852 ( .A1(n880), .A2(G95), .ZN(n766) );
  XOR2_X1 U853 ( .A(KEYINPUT87), .B(n766), .Z(n768) );
  NAND2_X1 U854 ( .A1(n882), .A2(G131), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U856 ( .A(KEYINPUT88), .B(n769), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n886), .A2(G107), .ZN(n770) );
  XOR2_X1 U858 ( .A(KEYINPUT86), .B(n770), .Z(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n889), .A2(G119), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n872) );
  AND2_X1 U862 ( .A1(n872), .A2(G1991), .ZN(n776) );
  AND2_X1 U863 ( .A1(n875), .A2(G1996), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n934) );
  INV_X1 U865 ( .A(n777), .ZN(n779) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U867 ( .A(n780), .B(KEYINPUT84), .ZN(n803) );
  XOR2_X1 U868 ( .A(KEYINPUT90), .B(n803), .Z(n781) );
  NOR2_X1 U869 ( .A1(n934), .A2(n781), .ZN(n800) );
  NOR2_X1 U870 ( .A1(G1986), .A2(G290), .ZN(n782) );
  NOR2_X1 U871 ( .A1(G1991), .A2(n872), .ZN(n927) );
  NOR2_X1 U872 ( .A1(n782), .A2(n927), .ZN(n783) );
  NOR2_X1 U873 ( .A1(n800), .A2(n783), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n924), .A2(n784), .ZN(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT39), .B(n785), .ZN(n796) );
  NAND2_X1 U876 ( .A1(G104), .A2(n880), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G140), .A2(n882), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(KEYINPUT34), .B(n788), .ZN(n794) );
  NAND2_X1 U880 ( .A1(n889), .A2(G128), .ZN(n789) );
  XOR2_X1 U881 ( .A(KEYINPUT85), .B(n789), .Z(n791) );
  NAND2_X1 U882 ( .A1(n886), .A2(G116), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U884 ( .A(KEYINPUT35), .B(n792), .Z(n793) );
  NOR2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n795), .ZN(n897) );
  XNOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .ZN(n797) );
  NOR2_X1 U888 ( .A1(n897), .A2(n797), .ZN(n944) );
  NAND2_X1 U889 ( .A1(n944), .A2(n803), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n796), .A2(n801), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n897), .A2(n797), .ZN(n941) );
  NAND2_X1 U892 ( .A1(n798), .A2(n941), .ZN(n799) );
  AND2_X1 U893 ( .A1(n799), .A2(n803), .ZN(n826) );
  INV_X1 U894 ( .A(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n805) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n990) );
  AND2_X1 U897 ( .A1(n990), .A2(n803), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U899 ( .A1(n807), .A2(n522), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n830) );
  NOR2_X1 U901 ( .A1(G1981), .A2(G305), .ZN(n810) );
  XOR2_X1 U902 ( .A(n810), .B(KEYINPUT24), .Z(n811) );
  OR2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n820) );
  INV_X1 U904 ( .A(n820), .ZN(n813) );
  OR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n817) );
  AND2_X1 U906 ( .A1(n814), .A2(n817), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n825) );
  INV_X1 U908 ( .A(n817), .ZN(n823) );
  NAND2_X1 U909 ( .A1(G8), .A2(G166), .ZN(n818) );
  NOR2_X1 U910 ( .A1(G2090), .A2(n818), .ZN(n819) );
  XNOR2_X1 U911 ( .A(n819), .B(KEYINPUT103), .ZN(n821) );
  AND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  OR2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n825), .A2(n824), .ZN(n827) );
  NOR2_X1 U915 ( .A1(n827), .A2(n826), .ZN(n828) );
  OR2_X1 U916 ( .A1(n828), .A2(n522), .ZN(n829) );
  NAND2_X1 U917 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U918 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n831) );
  XNOR2_X1 U919 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U922 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n835) );
  XNOR2_X1 U924 ( .A(KEYINPUT106), .B(n835), .ZN(n837) );
  NAND2_X1 U925 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U926 ( .A(n838), .ZN(G319) );
  XOR2_X1 U927 ( .A(KEYINPUT107), .B(G2090), .Z(n840) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2084), .ZN(n839) );
  XNOR2_X1 U929 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U930 ( .A(n841), .B(G2100), .Z(n843) );
  XNOR2_X1 U931 ( .A(G2072), .B(G2067), .ZN(n842) );
  XNOR2_X1 U932 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT43), .Z(n845) );
  XNOR2_X1 U934 ( .A(G2678), .B(KEYINPUT42), .ZN(n844) );
  XNOR2_X1 U935 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U936 ( .A(n847), .B(n846), .Z(G227) );
  XOR2_X1 U937 ( .A(G1976), .B(G1981), .Z(n849) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1971), .ZN(n848) );
  XNOR2_X1 U939 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U940 ( .A(n850), .B(G2474), .Z(n852) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U942 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1986), .Z(n854) );
  XNOR2_X1 U944 ( .A(G1961), .B(G1956), .ZN(n853) );
  XNOR2_X1 U945 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U946 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U947 ( .A1(G100), .A2(n880), .ZN(n858) );
  NAND2_X1 U948 ( .A1(G112), .A2(n886), .ZN(n857) );
  NAND2_X1 U949 ( .A1(n858), .A2(n857), .ZN(n863) );
  NAND2_X1 U950 ( .A1(n889), .A2(G124), .ZN(n859) );
  XNOR2_X1 U951 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U952 ( .A1(G136), .A2(n882), .ZN(n860) );
  NAND2_X1 U953 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U954 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U955 ( .A1(G115), .A2(n886), .ZN(n865) );
  NAND2_X1 U956 ( .A1(G127), .A2(n889), .ZN(n864) );
  NAND2_X1 U957 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U958 ( .A(n866), .B(KEYINPUT47), .ZN(n868) );
  NAND2_X1 U959 ( .A1(G139), .A2(n882), .ZN(n867) );
  NAND2_X1 U960 ( .A1(n868), .A2(n867), .ZN(n871) );
  NAND2_X1 U961 ( .A1(n880), .A2(G103), .ZN(n869) );
  XOR2_X1 U962 ( .A(KEYINPUT110), .B(n869), .Z(n870) );
  NOR2_X1 U963 ( .A1(n871), .A2(n870), .ZN(n935) );
  XOR2_X1 U964 ( .A(n872), .B(n935), .Z(n879) );
  XNOR2_X1 U965 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U966 ( .A(n873), .B(KEYINPUT48), .ZN(n874) );
  XOR2_X1 U967 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U968 ( .A(G160), .B(G164), .ZN(n876) );
  XNOR2_X1 U969 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U970 ( .A(n879), .B(n878), .ZN(n894) );
  NAND2_X1 U971 ( .A1(n880), .A2(G106), .ZN(n881) );
  XOR2_X1 U972 ( .A(KEYINPUT109), .B(n881), .Z(n884) );
  NAND2_X1 U973 ( .A1(n882), .A2(G142), .ZN(n883) );
  NAND2_X1 U974 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U975 ( .A(n885), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U976 ( .A1(G118), .A2(n886), .ZN(n887) );
  NAND2_X1 U977 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U978 ( .A1(n889), .A2(G130), .ZN(n890) );
  XOR2_X1 U979 ( .A(KEYINPUT108), .B(n890), .Z(n891) );
  NOR2_X1 U980 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U981 ( .A(n894), .B(n893), .Z(n896) );
  XNOR2_X1 U982 ( .A(G162), .B(n926), .ZN(n895) );
  XNOR2_X1 U983 ( .A(n896), .B(n895), .ZN(n898) );
  XNOR2_X1 U984 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U985 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U986 ( .A(G286), .B(KEYINPUT112), .Z(n900) );
  XNOR2_X1 U987 ( .A(n980), .B(n900), .ZN(n903) );
  XOR2_X1 U988 ( .A(G301), .B(n901), .Z(n902) );
  XNOR2_X1 U989 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U990 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U991 ( .A(G2430), .B(G2451), .Z(n906) );
  XNOR2_X1 U992 ( .A(G2446), .B(G2427), .ZN(n905) );
  XNOR2_X1 U993 ( .A(n906), .B(n905), .ZN(n913) );
  XOR2_X1 U994 ( .A(G2438), .B(KEYINPUT105), .Z(n908) );
  XNOR2_X1 U995 ( .A(G2443), .B(G2454), .ZN(n907) );
  XNOR2_X1 U996 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U997 ( .A(n909), .B(G2435), .Z(n911) );
  XNOR2_X1 U998 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U999 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1000 ( .A(n913), .B(n912), .ZN(n914) );
  NAND2_X1 U1001 ( .A1(n914), .A2(G14), .ZN(n922) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n922), .ZN(n917) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1005 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1007 ( .A1(n919), .A2(n918), .ZN(G225) );
  XNOR2_X1 U1008 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(G132), .ZN(G219) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  INV_X1 U1012 ( .A(G96), .ZN(G221) );
  INV_X1 U1013 ( .A(G82), .ZN(G220) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  INV_X1 U1017 ( .A(G108), .ZN(G238) );
  INV_X1 U1018 ( .A(n922), .ZN(G401) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n925), .Z(n929) );
  NOR2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n930) );
  XNOR2_X1 U1025 ( .A(KEYINPUT114), .B(n930), .ZN(n931) );
  NOR2_X1 U1026 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1028 ( .A(G2072), .B(n935), .Z(n937) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n936) );
  NOR2_X1 U1030 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n938), .Z(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1035 ( .A(KEYINPUT52), .B(n945), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(KEYINPUT55), .B(KEYINPUT115), .ZN(n968) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n968), .ZN(n947) );
  NAND2_X1 U1038 ( .A1(n947), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G35), .ZN(n963) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(G2067), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(n948), .B(G26), .ZN(n954) );
  XOR2_X1 U1042 ( .A(G2072), .B(G33), .Z(n949) );
  NAND2_X1 U1043 ( .A1(G28), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G25), .B(G1991), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT116), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n960) );
  XOR2_X1 U1048 ( .A(n955), .B(G27), .Z(n957) );
  XNOR2_X1 U1049 ( .A(G32), .B(G1996), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT118), .B(n958), .Z(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n961), .ZN(n962) );
  NOR2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1055 ( .A(G2084), .B(KEYINPUT54), .Z(n964) );
  XNOR2_X1 U1056 ( .A(G34), .B(n964), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n970) );
  INV_X1 U1059 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n971), .ZN(n1030) );
  XNOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  NAND2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(n974), .B(KEYINPUT121), .ZN(n997) );
  XOR2_X1 U1065 ( .A(G1966), .B(G168), .Z(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT119), .B(n975), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n978), .B(KEYINPUT57), .ZN(n992) );
  XNOR2_X1 U1069 ( .A(n979), .B(G1956), .ZN(n988) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(G1348), .B(n980), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT120), .ZN(n986) );
  XOR2_X1 U1074 ( .A(G1971), .B(G166), .Z(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT122), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G1341), .B(n993), .ZN(n994) );
  NOR2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1028) );
  INV_X1 U1084 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1085 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1024) );
  XNOR2_X1 U1086 ( .A(G1986), .B(G24), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n1000), .B(KEYINPUT124), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT125), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT126), .ZN(n1022) );
  XOR2_X1 U1095 ( .A(G1961), .B(G5), .Z(n1018) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(n1008), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1956), .B(G20), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1981), .B(G6), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT123), .B(G1341), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G19), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(KEYINPUT60), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G21), .B(G1966), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1114 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

