

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U323 ( .A(KEYINPUT48), .B(n514), .Z(n542) );
  NOR2_X1 U324 ( .A1(n513), .A2(n512), .ZN(n514) );
  AND2_X1 U325 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U326 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n431) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n543) );
  XNOR2_X1 U328 ( .A(n432), .B(n431), .ZN(n436) );
  XNOR2_X1 U329 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U330 ( .A(n441), .B(n291), .ZN(n442) );
  XNOR2_X1 U331 ( .A(n443), .B(n442), .ZN(n537) );
  XNOR2_X1 U332 ( .A(KEYINPUT94), .B(n406), .ZN(n546) );
  XNOR2_X1 U333 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n448) );
  XOR2_X1 U334 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n293) );
  XNOR2_X1 U335 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n294), .B(G155GAT), .Z(n296) );
  XNOR2_X1 U338 ( .A(G141GAT), .B(G148GAT), .ZN(n295) );
  XNOR2_X1 U339 ( .A(n296), .B(n295), .ZN(n363) );
  XOR2_X1 U340 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n298) );
  XNOR2_X1 U341 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n297) );
  XNOR2_X1 U342 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U343 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n300) );
  XNOR2_X1 U344 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U346 ( .A(n302), .B(n301), .Z(n312) );
  XNOR2_X1 U347 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n303), .B(KEYINPUT77), .ZN(n304) );
  XOR2_X1 U349 ( .A(n304), .B(KEYINPUT0), .Z(n306) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(G127GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n379) );
  XOR2_X1 U352 ( .A(G120GAT), .B(G57GAT), .Z(n338) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n307), .B(G85GAT), .ZN(n438) );
  XOR2_X1 U355 ( .A(n338), .B(n438), .Z(n309) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n379), .B(n310), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n363), .B(n313), .ZN(n406) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G141GAT), .Z(n315) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(G197GAT), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n332) );
  XOR2_X1 U364 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n317) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U366 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U367 ( .A(n318), .B(KEYINPUT30), .Z(n327) );
  INV_X1 U368 ( .A(KEYINPUT7), .ZN(n319) );
  NAND2_X1 U369 ( .A1(n319), .A2(G43GAT), .ZN(n322) );
  INV_X1 U370 ( .A(G43GAT), .ZN(n320) );
  NAND2_X1 U371 ( .A1(n320), .A2(KEYINPUT7), .ZN(n321) );
  NAND2_X1 U372 ( .A1(n322), .A2(n321), .ZN(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n432) );
  XNOR2_X1 U375 ( .A(G22GAT), .B(G15GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n325), .B(G1GAT), .ZN(n418) );
  XNOR2_X1 U377 ( .A(n432), .B(n418), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U379 ( .A(G169GAT), .B(G8GAT), .Z(n398) );
  XOR2_X1 U380 ( .A(n328), .B(n398), .Z(n330) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(G36GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U383 ( .A(n332), .B(n331), .Z(n475) );
  INV_X1 U384 ( .A(n475), .ZN(n570) );
  XOR2_X1 U385 ( .A(G99GAT), .B(G106GAT), .Z(n441) );
  XOR2_X1 U386 ( .A(KEYINPUT32), .B(G92GAT), .Z(n334) );
  XNOR2_X1 U387 ( .A(G148GAT), .B(G85GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U389 ( .A(n441), .B(n335), .Z(n340) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G204GAT), .Z(n337) );
  XNOR2_X1 U391 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n353) );
  XNOR2_X1 U393 ( .A(n353), .B(n338), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n347) );
  XOR2_X1 U395 ( .A(KEYINPUT69), .B(KEYINPUT31), .Z(n342) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U398 ( .A(n343), .B(KEYINPUT33), .Z(n345) );
  XOR2_X1 U399 ( .A(G176GAT), .B(G64GAT), .Z(n395) );
  XOR2_X1 U400 ( .A(G71GAT), .B(KEYINPUT13), .Z(n414) );
  XNOR2_X1 U401 ( .A(n395), .B(n414), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n575) );
  NAND2_X1 U404 ( .A1(n570), .A2(n575), .ZN(n462) );
  XOR2_X1 U405 ( .A(G211GAT), .B(KEYINPUT21), .Z(n349) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n392) );
  XOR2_X1 U408 ( .A(G50GAT), .B(G162GAT), .Z(n433) );
  XOR2_X1 U409 ( .A(n392), .B(n433), .Z(n351) );
  NAND2_X1 U410 ( .A1(G228GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U412 ( .A(n352), .B(KEYINPUT23), .Z(n355) );
  XNOR2_X1 U413 ( .A(n353), .B(KEYINPUT22), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U415 ( .A(KEYINPUT91), .B(KEYINPUT85), .Z(n357) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(G106GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U418 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U419 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n361) );
  XNOR2_X1 U420 ( .A(G22GAT), .B(KEYINPUT87), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n547) );
  XOR2_X1 U424 ( .A(G71GAT), .B(G190GAT), .Z(n367) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G134GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U427 ( .A(G43GAT), .B(G99GAT), .Z(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n383) );
  XOR2_X1 U429 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n371) );
  XNOR2_X1 U430 ( .A(G15GAT), .B(G176GAT), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U432 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n373) );
  XNOR2_X1 U433 ( .A(G120GAT), .B(KEYINPUT80), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U435 ( .A(n375), .B(n374), .Z(n381) );
  XOR2_X1 U436 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n377) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U439 ( .A(KEYINPUT19), .B(n378), .Z(n397) );
  XNOR2_X1 U440 ( .A(n397), .B(n379), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n385) );
  NAND2_X1 U443 ( .A1(G227GAT), .A2(G233GAT), .ZN(n384) );
  XOR2_X2 U444 ( .A(n385), .B(n384), .Z(n551) );
  NOR2_X1 U445 ( .A1(n547), .A2(n551), .ZN(n386) );
  XOR2_X1 U446 ( .A(KEYINPUT26), .B(n386), .Z(n567) );
  XOR2_X1 U447 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n388) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n388), .B(n387), .ZN(n391) );
  XOR2_X1 U450 ( .A(G92GAT), .B(G218GAT), .Z(n390) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G190GAT), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n390), .B(n389), .ZN(n437) );
  XOR2_X1 U453 ( .A(n391), .B(n437), .Z(n394) );
  XNOR2_X1 U454 ( .A(G204GAT), .B(n392), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U456 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n541) );
  XOR2_X1 U459 ( .A(n541), .B(KEYINPUT27), .Z(n407) );
  NOR2_X1 U460 ( .A1(n567), .A2(n407), .ZN(n527) );
  NAND2_X1 U461 ( .A1(n541), .A2(n551), .ZN(n401) );
  NAND2_X1 U462 ( .A1(n547), .A2(n401), .ZN(n402) );
  XNOR2_X1 U463 ( .A(KEYINPUT25), .B(n402), .ZN(n403) );
  NOR2_X1 U464 ( .A1(n527), .A2(n403), .ZN(n404) );
  XOR2_X1 U465 ( .A(KEYINPUT97), .B(n404), .Z(n405) );
  NOR2_X1 U466 ( .A1(n406), .A2(n405), .ZN(n410) );
  XOR2_X1 U467 ( .A(n547), .B(KEYINPUT28), .Z(n496) );
  NOR2_X1 U468 ( .A1(n407), .A2(n496), .ZN(n408) );
  NAND2_X1 U469 ( .A1(n546), .A2(n408), .ZN(n516) );
  NOR2_X1 U470 ( .A1(n551), .A2(n516), .ZN(n409) );
  NOR2_X1 U471 ( .A1(n410), .A2(n409), .ZN(n411) );
  XOR2_X1 U472 ( .A(KEYINPUT98), .B(n411), .Z(n459) );
  XOR2_X1 U473 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n445) );
  XOR2_X1 U474 ( .A(G57GAT), .B(G211GAT), .Z(n413) );
  XNOR2_X1 U475 ( .A(G127GAT), .B(G78GAT), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U477 ( .A(n415), .B(n414), .Z(n417) );
  XNOR2_X1 U478 ( .A(G183GAT), .B(G155GAT), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U480 ( .A(n418), .B(KEYINPUT12), .Z(n420) );
  NAND2_X1 U481 ( .A1(G231GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U483 ( .A(n422), .B(n421), .Z(n430) );
  XOR2_X1 U484 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n424) );
  XNOR2_X1 U485 ( .A(G8GAT), .B(G64GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n426) );
  XNOR2_X1 U488 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n578) );
  XNOR2_X1 U492 ( .A(n433), .B(KEYINPUT9), .ZN(n434) );
  XOR2_X1 U493 ( .A(n434), .B(KEYINPUT70), .Z(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n443) );
  XNOR2_X1 U497 ( .A(KEYINPUT71), .B(n537), .ZN(n561) );
  NAND2_X1 U498 ( .A1(n578), .A2(n561), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n459), .A2(n446), .ZN(n476) );
  NOR2_X1 U501 ( .A1(n462), .A2(n476), .ZN(n454) );
  NAND2_X1 U502 ( .A1(n546), .A2(n454), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(G1324GAT) );
  XOR2_X1 U504 ( .A(G8GAT), .B(KEYINPUT99), .Z(n450) );
  NAND2_X1 U505 ( .A1(n454), .A2(n541), .ZN(n449) );
  XNOR2_X1 U506 ( .A(n450), .B(n449), .ZN(G1325GAT) );
  XOR2_X1 U507 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n452) );
  NAND2_X1 U508 ( .A1(n454), .A2(n551), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U510 ( .A(G15GAT), .B(n453), .ZN(G1326GAT) );
  XOR2_X1 U511 ( .A(G22GAT), .B(KEYINPUT101), .Z(n456) );
  NAND2_X1 U512 ( .A1(n454), .A2(n496), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(G1327GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT102), .B(KEYINPUT39), .Z(n465) );
  XNOR2_X1 U515 ( .A(KEYINPUT37), .B(KEYINPUT103), .ZN(n457) );
  XNOR2_X1 U516 ( .A(n457), .B(KEYINPUT104), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT36), .B(n561), .ZN(n502) );
  NOR2_X1 U518 ( .A1(n502), .A2(n578), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n461), .B(n460), .ZN(n489) );
  NOR2_X1 U521 ( .A1(n462), .A2(n489), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT38), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n546), .A2(n470), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U525 ( .A(G29GAT), .B(n466), .ZN(G1328GAT) );
  NAND2_X1 U526 ( .A1(n470), .A2(n541), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U528 ( .A1(n470), .A2(n551), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT40), .ZN(n469) );
  XNOR2_X1 U530 ( .A(G43GAT), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U531 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n472) );
  NAND2_X1 U532 ( .A1(n496), .A2(n470), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U534 ( .A(G50GAT), .B(n473), .ZN(G1331GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n479) );
  XNOR2_X1 U536 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n474) );
  XNOR2_X1 U537 ( .A(n575), .B(n474), .ZN(n554) );
  NAND2_X1 U538 ( .A1(n475), .A2(n554), .ZN(n488) );
  NOR2_X1 U539 ( .A1(n488), .A2(n476), .ZN(n477) );
  XOR2_X1 U540 ( .A(KEYINPUT107), .B(n477), .Z(n485) );
  NAND2_X1 U541 ( .A1(n485), .A2(n546), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U543 ( .A(G57GAT), .B(n480), .Z(G1332GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n482) );
  NAND2_X1 U545 ( .A1(n485), .A2(n541), .ZN(n481) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U547 ( .A(G64GAT), .B(n483), .ZN(G1333GAT) );
  NAND2_X1 U548 ( .A1(n551), .A2(n485), .ZN(n484) );
  XNOR2_X1 U549 ( .A(n484), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U550 ( .A(G78GAT), .B(KEYINPUT43), .Z(n487) );
  NAND2_X1 U551 ( .A1(n485), .A2(n496), .ZN(n486) );
  XNOR2_X1 U552 ( .A(n487), .B(n486), .ZN(G1335GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n491) );
  NOR2_X1 U554 ( .A1(n489), .A2(n488), .ZN(n497) );
  NAND2_X1 U555 ( .A1(n497), .A2(n546), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U557 ( .A(G85GAT), .B(n492), .ZN(G1336GAT) );
  NAND2_X1 U558 ( .A1(n497), .A2(n541), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n493), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U560 ( .A(G99GAT), .B(KEYINPUT113), .Z(n495) );
  NAND2_X1 U561 ( .A1(n497), .A2(n551), .ZN(n494) );
  XNOR2_X1 U562 ( .A(n495), .B(n494), .ZN(G1338GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n499) );
  NAND2_X1 U564 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U566 ( .A(G106GAT), .B(n500), .Z(G1339GAT) );
  INV_X1 U567 ( .A(n578), .ZN(n501) );
  NOR2_X1 U568 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(KEYINPUT45), .ZN(n506) );
  INV_X1 U570 ( .A(n575), .ZN(n504) );
  NOR2_X1 U571 ( .A1(n570), .A2(n504), .ZN(n505) );
  AND2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n513) );
  NOR2_X1 U573 ( .A1(n537), .A2(n578), .ZN(n510) );
  XOR2_X1 U574 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n508) );
  AND2_X1 U575 ( .A1(n570), .A2(n554), .ZN(n507) );
  XOR2_X1 U576 ( .A(n508), .B(n507), .Z(n509) );
  NAND2_X1 U577 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(KEYINPUT47), .ZN(n512) );
  NAND2_X1 U579 ( .A1(n542), .A2(n551), .ZN(n515) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n570), .A2(n524), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(G120GAT), .B(KEYINPUT49), .Z(n519) );
  NAND2_X1 U584 ( .A1(n524), .A2(n554), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1341GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n521) );
  NAND2_X1 U587 ( .A1(n524), .A2(n578), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U589 ( .A(G127GAT), .B(n522), .Z(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n526) );
  INV_X1 U591 ( .A(n561), .ZN(n523) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  INV_X1 U594 ( .A(n546), .ZN(n529) );
  NAND2_X1 U595 ( .A1(n542), .A2(n527), .ZN(n528) );
  NOR2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n538), .A2(n570), .ZN(n530) );
  XNOR2_X1 U598 ( .A(G141GAT), .B(n530), .ZN(G1344GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n532) );
  NAND2_X1 U600 ( .A1(n538), .A2(n554), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n534) );
  XOR2_X1 U602 ( .A(G148GAT), .B(KEYINPUT117), .Z(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n578), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n535), .B(KEYINPUT118), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G155GAT), .B(n536), .ZN(G1346GAT) );
  XOR2_X1 U607 ( .A(G162GAT), .B(KEYINPUT119), .Z(n540) );
  NAND2_X1 U608 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n540), .B(n539), .ZN(G1347GAT) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n568) );
  NAND2_X1 U612 ( .A1(n568), .A2(n547), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT121), .ZN(n549) );
  XOR2_X1 U614 ( .A(n549), .B(KEYINPUT55), .Z(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n562) );
  INV_X1 U616 ( .A(n562), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n559), .A2(n570), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n552), .B(KEYINPUT122), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U620 ( .A1(n559), .A2(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .Z(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n559), .A2(n578), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n566) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(KEYINPUT124), .ZN(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT125), .B(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1351GAT) );
  INV_X1 U632 ( .A(n567), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n581) );
  INV_X1 U634 ( .A(n581), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n570), .A2(n579), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  OR2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n502), .A2(n581), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

