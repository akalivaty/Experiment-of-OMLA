//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n637, new_n638, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G57), .Z(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  OR2_X1    g039(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n472), .A3(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT72), .B1(new_n477), .B2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n482));
  OAI21_X1  g057(.A(G137), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n474), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(KEYINPUT73), .B(new_n474), .C1(new_n480), .C2(new_n483), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n471), .B1(new_n486), .B2(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n467), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n480), .A2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G124), .ZN(new_n493));
  XOR2_X1   g068(.A(new_n493), .B(KEYINPUT74), .Z(new_n494));
  INV_X1    g069(.A(new_n480), .ZN(new_n495));
  INV_X1    g070(.A(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n491), .B(new_n494), .C1(G136), .C2(new_n498), .ZN(G162));
  OAI211_X1 g074(.A(G126), .B(new_n476), .C1(new_n478), .C2(new_n479), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n467), .A2(new_n468), .A3(G138), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n504), .A2(new_n505), .B1(G102), .B2(new_n473), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n507), .B1(new_n465), .B2(new_n466), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n475), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n508), .A2(new_n511), .A3(KEYINPUT4), .A4(new_n476), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n503), .A2(new_n506), .A3(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(G164));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(new_n517), .B2(G651), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n519), .A2(KEYINPUT75), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT6), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT75), .B1(new_n519), .B2(KEYINPUT76), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n521), .A2(G543), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n521), .A2(new_n526), .A3(new_n524), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n515), .A2(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(G62), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(new_n531), .B1(G75), .B2(G543), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(KEYINPUT77), .A3(G62), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n529), .A2(new_n534), .ZN(G166));
  NAND3_X1  g110(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT78), .Z(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT7), .Z(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G651), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n523), .B1(new_n522), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT5), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT5), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n517), .A2(G651), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT6), .B1(new_n548), .B2(KEYINPUT75), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n542), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G89), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G51), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n540), .A2(new_n551), .A3(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  NAND2_X1  g130(.A1(new_n550), .A2(G90), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(G52), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n519), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G56), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n547), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n552), .A2(G43), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n550), .A2(G81), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  NAND4_X1  g149(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n524), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n521), .A2(G91), .A3(new_n526), .A4(new_n524), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n547), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n577), .A2(KEYINPUT79), .B1(G651), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n576), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT80), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n578), .A2(new_n582), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n585), .A2(new_n586), .A3(new_n576), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G166), .ZN(G303));
  INV_X1    g164(.A(G74), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n519), .B1(new_n547), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n552), .B2(G49), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT81), .ZN(new_n593));
  INV_X1    g168(.A(G87), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n527), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n550), .A2(KEYINPUT81), .A3(G87), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(KEYINPUT82), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G288));
  NAND4_X1  g176(.A1(new_n521), .A2(G86), .A3(new_n526), .A4(new_n524), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n521), .A2(G48), .A3(G543), .A4(new_n524), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n526), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n519), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n544), .A2(new_n546), .A3(G61), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n610), .A2(KEYINPUT83), .A3(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n604), .B1(new_n612), .B2(KEYINPUT84), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(G305));
  NAND2_X1  g191(.A1(new_n550), .A2(G85), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n552), .A2(G47), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n617), .B(new_n618), .C1(new_n519), .C2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(new_n550), .A2(G92), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n547), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n552), .A2(G54), .B1(G651), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(G301), .A2(G868), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n628), .A2(new_n629), .B1(KEYINPUT85), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(KEYINPUT85), .B2(new_n630), .ZN(G284));
  OAI21_X1  g207(.A(new_n631), .B1(KEYINPUT85), .B2(new_n630), .ZN(G321));
  NAND2_X1  g208(.A1(G299), .A2(new_n629), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(G168), .ZN(G280));
  XNOR2_X1  g210(.A(G280), .B(KEYINPUT86), .ZN(G297));
  AND2_X1   g211(.A1(new_n623), .A2(new_n627), .ZN(new_n637));
  INV_X1    g212(.A(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G860), .ZN(G148));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n492), .A2(G123), .ZN(new_n644));
  OAI221_X1 g219(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n467), .C2(G111), .ZN(new_n645));
  INV_X1    g220(.A(G135), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n644), .B(new_n645), .C1(new_n497), .C2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2096), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n468), .A2(new_n473), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2430), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2435), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(KEYINPUT14), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2451), .B(G2454), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  XOR2_X1   g242(.A(G1341), .B(G1348), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n669), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(KEYINPUT92), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n673), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n675), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n673), .B(KEYINPUT17), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n682), .B(new_n683), .C1(new_n681), .C2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G2096), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G227));
  XNOR2_X1  g263(.A(G1971), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT19), .ZN(new_n690));
  XOR2_X1   g265(.A(G1956), .B(G2474), .Z(new_n691));
  XOR2_X1   g266(.A(G1961), .B(G1966), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT20), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n691), .B2(new_n692), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n690), .A2(KEYINPUT93), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT94), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT95), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(G229));
  MUX2_X1   g284(.A(G6), .B(G305), .S(G16), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G23), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n710), .A2(new_n711), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1971), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n715), .A2(new_n716), .ZN(new_n723));
  NOR4_X1   g298(.A1(new_n717), .A2(new_n718), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT34), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n719), .A2(G24), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G290), .B2(G16), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1986), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n492), .A2(G119), .ZN(new_n730));
  OAI221_X1 g305(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n467), .C2(G107), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n497), .C2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G25), .B(new_n733), .S(G29), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT35), .B(G1991), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n728), .A2(G1986), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n725), .A2(new_n729), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT36), .ZN(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n741), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(G2090), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(G2090), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n719), .A2(G4), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n637), .B2(new_n719), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1348), .ZN(new_n749));
  NOR3_X1   g324(.A1(new_n745), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n719), .A2(G20), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n751), .B(new_n752), .C1(G299), .C2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  INV_X1    g329(.A(G1956), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n568), .A2(new_n719), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n719), .B2(G19), .ZN(new_n758));
  INV_X1    g333(.A(G1341), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  NAND2_X1  g335(.A1(G171), .A2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G5), .B2(G16), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n759), .B2(new_n758), .ZN(new_n764));
  NOR2_X1   g339(.A1(G168), .A2(new_n719), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n719), .B2(G21), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(G34), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G160), .B2(new_n741), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n762), .A2(new_n760), .B1(G2084), .B2(new_n774), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n764), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n741), .A2(G33), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n467), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT25), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n781), .B(new_n783), .C1(G139), .C2(new_n498), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n779), .B1(new_n784), .B2(new_n741), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G2072), .Z(new_n786));
  INV_X1    g361(.A(G28), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT30), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(KEYINPUT30), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n647), .B2(new_n741), .ZN(new_n793));
  NOR2_X1   g368(.A1(G29), .A2(G32), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n498), .A2(G141), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n492), .A2(G129), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n473), .A2(G105), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n798));
  NAND3_X1  g373(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n795), .A2(new_n796), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n794), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT27), .B(G1996), .Z(new_n805));
  AOI21_X1  g380(.A(new_n793), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n786), .B(new_n806), .C1(new_n804), .C2(new_n805), .ZN(new_n807));
  NOR2_X1   g382(.A1(G27), .A2(G29), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G164), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2078), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n766), .B2(new_n767), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n741), .A2(G26), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n492), .A2(G128), .ZN(new_n814));
  OAI221_X1 g389(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n467), .C2(G116), .ZN(new_n815));
  INV_X1    g390(.A(G140), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n814), .B(new_n815), .C1(new_n497), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n813), .B1(new_n817), .B2(G29), .ZN(new_n818));
  MUX2_X1   g393(.A(new_n813), .B(new_n818), .S(KEYINPUT28), .Z(new_n819));
  INV_X1    g394(.A(G2067), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n778), .A2(new_n807), .A3(new_n812), .A4(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n750), .A2(new_n756), .A3(new_n822), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n740), .A2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n740), .A2(new_n823), .ZN(G150));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  INV_X1    g401(.A(G80), .ZN(new_n827));
  OAI22_X1  g402(.A1(new_n547), .A2(new_n826), .B1(new_n827), .B2(new_n543), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI221_X1 g405(.A(KEYINPUT98), .B1(new_n827), .B2(new_n543), .C1(new_n547), .C2(new_n826), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(G651), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT99), .ZN(new_n834));
  AOI22_X1  g409(.A1(G55), .A2(new_n552), .B1(new_n550), .B2(G93), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n637), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n836), .A2(new_n568), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n833), .A2(new_n567), .A3(new_n834), .A4(new_n835), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n840), .B(new_n843), .Z(new_n844));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n845));
  AOI21_X1  g420(.A(G860), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(KEYINPUT100), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n847), .A2(KEYINPUT100), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n838), .B1(new_n848), .B2(new_n849), .ZN(G145));
  NAND2_X1  g425(.A1(new_n492), .A2(G130), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n467), .C2(G118), .ZN(new_n852));
  INV_X1    g427(.A(G142), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n851), .B(new_n852), .C1(new_n497), .C2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(new_n651), .Z(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n817), .B(new_n733), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n802), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n857), .A2(new_n802), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n817), .B(new_n733), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n803), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(new_n855), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(G138), .B1(new_n481), .B2(new_n482), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n477), .A2(G2104), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n510), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n505), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n473), .A2(G102), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n512), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT101), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n503), .A2(new_n506), .A3(new_n874), .A4(new_n512), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n865), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n861), .A2(new_n877), .A3(new_n864), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n784), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n784), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G160), .B(new_n647), .ZN(new_n884));
  XNOR2_X1  g459(.A(G162), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n881), .A2(new_n888), .A3(new_n885), .A4(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  XOR2_X1   g469(.A(G305), .B(G290), .Z(new_n895));
  XNOR2_X1  g470(.A(G166), .B(new_n597), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(KEYINPUT103), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n843), .B(new_n640), .ZN(new_n907));
  NOR2_X1   g482(.A1(G299), .A2(new_n628), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n637), .B1(new_n584), .B2(new_n587), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n908), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n628), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n637), .A2(new_n584), .A3(new_n587), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(KEYINPUT41), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n907), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n906), .A2(new_n912), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(new_n904), .A3(new_n905), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(G868), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n836), .A2(new_n629), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n894), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n925), .ZN(new_n927));
  AOI211_X1 g502(.A(KEYINPUT104), .B(new_n927), .C1(new_n923), .C2(G868), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g506(.A1(G286), .A2(G171), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n540), .A2(new_n551), .A3(new_n553), .A4(G301), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n843), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n841), .A2(new_n932), .A3(new_n842), .A4(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n914), .A2(new_n917), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n914), .A2(new_n937), .A3(new_n940), .A4(new_n917), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n935), .A2(new_n915), .A3(new_n916), .A4(new_n936), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n899), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n938), .A2(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n947), .B2(new_n900), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(KEYINPUT107), .A3(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n931), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n946), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n942), .A2(new_n945), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n900), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT44), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n931), .B1(new_n955), .B2(new_n957), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(KEYINPUT127), .ZN(new_n965));
  INV_X1    g540(.A(G1996), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n803), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n817), .B(G2067), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n802), .A2(G1996), .ZN(new_n969));
  OR3_X1    g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(new_n877), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n971), .B1(new_n972), .B2(G1384), .ZN(new_n973));
  INV_X1    g548(.A(new_n471), .ZN(new_n974));
  INV_X1    g549(.A(new_n487), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n511), .A2(G137), .A3(new_n467), .A4(new_n476), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT73), .B1(new_n976), .B2(new_n474), .ZN(new_n977));
  OAI211_X1 g552(.A(G40), .B(new_n974), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n970), .A2(KEYINPUT108), .A3(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n733), .B(new_n736), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT109), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  AND2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n979), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n871), .B2(new_n872), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n978), .B1(new_n971), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n877), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT56), .B(G2072), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n992), .C1(new_n871), .C2(new_n872), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(G160), .A3(G40), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n513), .B2(new_n992), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT117), .B(new_n755), .C1(new_n1000), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n993), .A2(new_n1001), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n1007), .B(new_n471), .C1(new_n486), .C2(new_n487), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1008), .A3(new_n999), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT117), .B1(new_n1009), .B2(new_n755), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n997), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n755), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1004), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(KEYINPUT119), .A3(new_n997), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT57), .B1(new_n576), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n583), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n585), .B(new_n576), .C1(new_n1019), .C2(KEYINPUT57), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1013), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n997), .B(new_n1023), .C1(new_n1005), .C2(new_n1010), .ZN(new_n1026));
  INV_X1    g601(.A(G1348), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n992), .B(new_n1002), .C1(new_n871), .C2(new_n872), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(G160), .A3(G40), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n998), .B1(new_n513), .B2(new_n992), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n978), .A2(new_n993), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n820), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n628), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1025), .B1(new_n1026), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1035), .A2(KEYINPUT60), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1031), .A2(KEYINPUT60), .A3(new_n1033), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT122), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n637), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1031), .A2(new_n1033), .A3(KEYINPUT60), .A4(new_n628), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n1039), .B2(new_n637), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT123), .B(new_n1038), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1039), .A2(new_n637), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT122), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1048), .A2(new_n1042), .A3(new_n1041), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT123), .B1(new_n1049), .B2(new_n1038), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1011), .A2(new_n1024), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1026), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT61), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n994), .A2(new_n995), .A3(new_n966), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT58), .B(G1341), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1032), .B2(new_n1057), .ZN(new_n1058));
  AND4_X1   g633(.A1(KEYINPUT120), .A2(new_n1058), .A3(KEYINPUT59), .A4(new_n568), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1058), .A2(new_n568), .B1(KEYINPUT120), .B2(KEYINPUT59), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1026), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1017), .A2(KEYINPUT121), .A3(new_n997), .A4(new_n1023), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(KEYINPUT61), .A3(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1055), .B(new_n1061), .C1(new_n1025), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1037), .B1(new_n1051), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n994), .A2(new_n995), .A3(new_n810), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1030), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n1008), .A3(new_n1028), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1069), .A2(new_n1070), .B1(new_n760), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1070), .A2(G2078), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n973), .A2(new_n1008), .A3(new_n995), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1076), .B2(G171), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n513), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n994), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(new_n1078), .A3(G301), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1072), .A2(new_n760), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n1080), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT124), .B1(new_n1084), .B2(G171), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1077), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(G171), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1073), .A2(G301), .A3(new_n1075), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n993), .A2(new_n971), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(new_n1008), .A3(new_n1079), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n768), .B1(new_n1092), .B2(new_n767), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G286), .A2(G8), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G8), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1093), .B2(G168), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT51), .B(new_n1094), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1089), .A2(new_n1068), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(G1971), .B1(new_n994), .B2(new_n995), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1009), .A2(G2090), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT115), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1104), .A2(new_n1111), .A3(new_n1108), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n713), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n1114));
  INV_X1    g689(.A(G1976), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n597), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(G160), .A2(G40), .A3(new_n992), .A4(new_n513), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1113), .A2(G8), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT52), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(KEYINPUT112), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1032), .A2(new_n1096), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1123), .A2(new_n1113), .A3(new_n1120), .A4(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1119), .A2(new_n1115), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n599), .B2(new_n600), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1122), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT83), .B1(new_n610), .B2(G651), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n605), .B(new_n519), .C1(new_n608), .C2(new_n609), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT84), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n602), .A2(new_n603), .ZN(new_n1132));
  INV_X1    g707(.A(G1981), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n615), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT113), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT113), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n613), .A2(new_n1136), .A3(new_n1133), .A4(new_n615), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n612), .B1(KEYINPUT114), .B2(new_n604), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n604), .A2(KEYINPUT114), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G1981), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1123), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1135), .A2(new_n1137), .B1(new_n1141), .B2(G1981), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1146), .A2(KEYINPUT49), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1128), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT116), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1110), .A2(new_n1112), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(G1971), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n971), .B(G1384), .C1(new_n873), .C2(new_n875), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1091), .A2(new_n1008), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OR3_X1    g729(.A1(new_n1029), .A2(new_n1030), .A3(G2090), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1096), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1123), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1146), .B2(KEYINPUT49), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1126), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1160), .A2(new_n1161), .B1(new_n1162), .B2(new_n1124), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1158), .B1(new_n1163), .B2(KEYINPUT116), .ZN(new_n1164));
  AND4_X1   g739(.A1(new_n1086), .A2(new_n1101), .A3(new_n1150), .A4(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1067), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1092), .A2(new_n767), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1071), .A2(new_n1008), .A3(new_n768), .A4(new_n1028), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1171), .A2(G8), .A3(G168), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1172), .A2(KEYINPUT63), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1163), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT63), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G288), .A2(G1976), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1159), .B1(new_n1180), .B2(new_n1138), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1148), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1174), .A2(new_n1178), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1098), .B(G8), .C1(new_n1171), .C2(G286), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1171), .A2(G8), .A3(G286), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1187), .A2(new_n1100), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT62), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1087), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1187), .A2(new_n1100), .A3(new_n1192), .A4(new_n1188), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1185), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n991), .B1(new_n1166), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n979), .A2(new_n988), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT48), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n987), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n979), .B1(new_n802), .B2(new_n968), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT126), .Z(new_n1202));
  INV_X1    g777(.A(KEYINPUT47), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n979), .A2(new_n966), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT46), .ZN(new_n1205));
  AND3_X1   g780(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1203), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1200), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n1209));
  NOR2_X1   g784(.A1(new_n733), .A2(new_n735), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n982), .A2(new_n983), .A3(new_n1210), .ZN(new_n1211));
  OR2_X1    g786(.A1(new_n817), .A2(G2067), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1209), .B1(new_n1213), .B2(new_n979), .ZN(new_n1214));
  INV_X1    g789(.A(new_n979), .ZN(new_n1215));
  AOI211_X1 g790(.A(KEYINPUT125), .B(new_n1215), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  OR2_X1    g792(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n965), .B1(new_n1197), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n991), .ZN(new_n1220));
  NAND4_X1  g795(.A1(new_n1101), .A2(new_n1150), .A3(new_n1086), .A4(new_n1164), .ZN(new_n1221));
  AOI21_X1  g796(.A(KEYINPUT61), .B1(new_n1052), .B2(new_n1026), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1222), .A2(new_n1060), .A3(new_n1059), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1013), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1224), .A2(KEYINPUT61), .A3(new_n1064), .A4(new_n1063), .ZN(new_n1225));
  OAI211_X1 g800(.A(new_n1223), .B(new_n1225), .C1(new_n1050), .C2(new_n1046), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1221), .B1(new_n1226), .B2(new_n1037), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT63), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1228), .B1(new_n1176), .B2(new_n1163), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1229), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1230));
  OAI211_X1 g805(.A(new_n1230), .B(new_n1174), .C1(new_n1186), .C2(new_n1194), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1220), .B1(new_n1227), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g807(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1232), .A2(KEYINPUT127), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1219), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g810(.A1(new_n961), .A2(new_n962), .ZN(new_n1237));
  NOR4_X1   g811(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n892), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1237), .A2(new_n1239), .ZN(G308));
  OR2_X1    g814(.A1(new_n1237), .A2(new_n1239), .ZN(G225));
endmodule


