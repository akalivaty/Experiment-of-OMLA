//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT70), .ZN(new_n205));
  AND2_X1   g004(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g012(.A(G127gat), .B(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n211), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT69), .B(G113gat), .ZN(new_n216));
  OAI211_X1 g015(.A(KEYINPUT70), .B(new_n215), .C1(new_n216), .C2(new_n208), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G134gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G127gat), .ZN(new_n220));
  INV_X1    g019(.A(G127gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G134gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n208), .A2(G113gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n213), .B1(new_n211), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT68), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT67), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT67), .B1(new_n220), .B2(new_n222), .ZN(new_n232));
  OAI211_X1 g031(.A(KEYINPUT68), .B(new_n229), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n218), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n229), .B1(new_n231), .B2(new_n232), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT71), .A3(new_n218), .ZN(new_n242));
  NAND2_X1  g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT65), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT24), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  AND2_X1   g048(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G169gat), .ZN(new_n253));
  INV_X1    g052(.A(G176gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258));
  AND4_X1   g057(.A1(KEYINPUT25), .A2(new_n255), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n247), .ZN(new_n262));
  INV_X1    g061(.A(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n260), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT26), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n272), .B(new_n243), .C1(new_n274), .C2(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT27), .ZN(new_n277));
  AOI21_X1  g076(.A(G190gat), .B1(new_n277), .B2(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT27), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT66), .B(new_n264), .C1(new_n263), .C2(KEYINPUT27), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n280), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n281), .A2(new_n278), .A3(new_n284), .A4(new_n279), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n276), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n237), .A2(new_n242), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n237), .B2(new_n242), .ZN(new_n291));
  OAI211_X1 g090(.A(G227gat), .B(G233gat), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n204), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n291), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n297), .B2(new_n289), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n294), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n292), .B(KEYINPUT32), .C1(new_n293), .C2(new_n204), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n296), .A3(new_n289), .ZN(new_n305));
  XOR2_X1   g104(.A(new_n305), .B(KEYINPUT34), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n312), .B(new_n311), .C1(new_n309), .C2(KEYINPUT2), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G197gat), .B(G204gat), .Z(new_n318));
  AOI21_X1  g117(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321));
  OR3_X1    g120(.A1(new_n320), .A2(KEYINPUT73), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n321), .B1(new_n320), .B2(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n317), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G228gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n324), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n326), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n323), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(KEYINPUT81), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  INV_X1    g137(.A(new_n336), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n338), .B1(new_n339), .B2(new_n327), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G22gat), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n320), .A2(new_n321), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n323), .B1(new_n320), .B2(new_n321), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n326), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n315), .A2(new_n316), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n333), .A2(new_n335), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n332), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n342), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n350), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G22gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n341), .A2(new_n355), .A3(new_n342), .A4(new_n350), .ZN(new_n356));
  XNOR2_X1  g155(.A(G78gat), .B(G106gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT31), .B(G50gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n352), .A2(new_n354), .A3(new_n356), .A4(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n359), .B(KEYINPUT80), .Z(new_n362));
  INV_X1    g161(.A(new_n351), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n342), .B1(new_n341), .B2(new_n350), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(KEYINPUT29), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n270), .A2(new_n369), .A3(new_n286), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n270), .B2(new_n286), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n270), .A2(new_n367), .A3(new_n286), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n333), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(new_n255), .A3(new_n258), .A4(new_n257), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(new_n261), .B1(new_n252), .B2(new_n259), .ZN(new_n378));
  INV_X1    g177(.A(new_n285), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n281), .A2(new_n284), .B1(new_n278), .B2(new_n279), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(new_n275), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT74), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(new_n367), .A3(new_n370), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n287), .A2(new_n368), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n383), .A2(new_n333), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n375), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n389), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n375), .B2(new_n385), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n386), .A2(KEYINPUT30), .A3(new_n389), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n306), .A2(new_n302), .A3(new_n303), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n308), .A2(new_n366), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  XOR2_X1   g199(.A(G1gat), .B(G29gat), .Z(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G57gat), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n317), .A4(new_n242), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n346), .B(new_n326), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n235), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n317), .B(new_n218), .C1(new_n230), .C2(new_n234), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n407), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n235), .A2(new_n346), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n412), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(new_n409), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n406), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n237), .A2(new_n413), .A3(new_n317), .A4(new_n242), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT77), .B1(new_n412), .B2(KEYINPUT4), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n412), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n411), .A2(new_n416), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT78), .B1(new_n424), .B2(new_n425), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n420), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n415), .A2(new_n419), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n425), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n430), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n400), .B(new_n428), .C1(new_n435), .C2(new_n405), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n429), .B1(new_n426), .B2(new_n427), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n406), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT35), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n399), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n395), .A2(new_n394), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n394), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n392), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n429), .A2(new_n405), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n433), .B2(new_n434), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT79), .B1(new_n449), .B2(KEYINPUT6), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n437), .A2(new_n406), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n452), .A3(new_n400), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n447), .B1(new_n454), .B2(new_n438), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n361), .A2(new_n365), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n306), .A2(new_n302), .A3(new_n303), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n306), .B1(new_n302), .B2(new_n303), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n442), .B1(new_n460), .B2(KEYINPUT35), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n457), .B2(new_n458), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n308), .A2(new_n398), .A3(KEYINPUT36), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n393), .A2(KEYINPUT37), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n394), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n333), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n383), .A2(new_n468), .A3(new_n384), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n469), .A2(KEYINPUT37), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n373), .A2(new_n374), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n333), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT38), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n383), .A2(new_n333), .A3(new_n384), .ZN(new_n476));
  INV_X1    g275(.A(new_n374), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n382), .A2(new_n370), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n477), .B1(new_n478), .B2(new_n368), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(new_n333), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n393), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT37), .B(new_n469), .C1(new_n479), .C2(new_n468), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT38), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n475), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n474), .A2(new_n485), .A3(new_n390), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n436), .A3(new_n438), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT86), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n486), .A2(new_n436), .A3(new_n489), .A4(new_n438), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n467), .B1(new_n491), .B2(new_n386), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT38), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n492), .B2(KEYINPUT38), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n488), .A2(new_n490), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n410), .A2(new_n235), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n424), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n409), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n417), .A2(new_n412), .A3(new_n408), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT39), .B1(new_n501), .B2(KEYINPUT84), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(KEYINPUT84), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n409), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n405), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n451), .A2(new_n396), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n508), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n456), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n465), .B1(new_n497), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n451), .A2(new_n400), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n428), .A2(new_n400), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n516), .A2(KEYINPUT79), .B1(new_n437), .B2(new_n406), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n515), .B1(new_n517), .B2(new_n453), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n456), .B1(new_n518), .B2(new_n447), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n461), .B1(new_n514), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G29gat), .A2(G36gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(KEYINPUT15), .A3(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n521), .B(KEYINPUT90), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n524), .A2(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n524), .A2(KEYINPUT89), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n523), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n527), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT17), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(G1gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G1gat), .B2(new_n537), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(G8gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n535), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT91), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT18), .B1(new_n546), .B2(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT93), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT92), .B1(new_n541), .B2(new_n535), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n545), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n544), .B(KEYINPUT13), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n546), .ZN(new_n556));
  XOR2_X1   g355(.A(G113gat), .B(G141gat), .Z(new_n557));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT12), .Z(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT93), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n565), .A3(new_n548), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n549), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n563), .B1(new_n568), .B2(new_n556), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n520), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT7), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT7), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(G85gat), .A3(G92gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n573), .A2(KEYINPUT97), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G99gat), .ZN(new_n579));
  INV_X1    g378(.A(G106gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT8), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(KEYINPUT96), .B(G85gat), .Z(new_n582));
  OAI211_X1 g381(.A(new_n578), .B(new_n581), .C1(G92gat), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n573), .A2(KEYINPUT97), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n536), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n586), .ZN(new_n589));
  AND2_X1   g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n589), .A2(new_n535), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G134gat), .ZN(new_n599));
  INV_X1    g398(.A(G162gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n594), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n597), .A2(new_n601), .B1(new_n602), .B2(new_n595), .ZN(new_n603));
  AND4_X1   g402(.A1(KEYINPUT98), .A2(new_n595), .A3(new_n602), .A4(new_n601), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G57gat), .B(G64gat), .Z(new_n607));
  INV_X1    g406(.A(KEYINPUT9), .ZN(new_n608));
  INV_X1    g407(.A(G71gat), .ZN(new_n609));
  INV_X1    g408(.A(G78gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G71gat), .B(G78gat), .Z(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G127gat), .B(G155gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT94), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n620), .B(new_n622), .Z(new_n623));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n616), .B(KEYINPUT95), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n542), .B1(new_n626), .B2(new_n617), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n606), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G230gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(new_n330), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n589), .A2(new_n616), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n585), .A2(new_n586), .A3(new_n615), .A4(new_n614), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n587), .A2(new_n626), .A3(new_n641), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n637), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n637), .A3(new_n639), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n635), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT10), .B1(new_n638), .B2(new_n639), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n587), .A2(new_n626), .A3(new_n641), .ZN(new_n649));
  OAI22_X1  g448(.A1(new_n648), .A2(new_n649), .B1(new_n636), .B2(new_n330), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n650), .A2(new_n651), .A3(new_n634), .A4(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT100), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n631), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n572), .A2(new_n518), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g461(.A1(new_n572), .A2(new_n660), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n397), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n396), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n669));
  AND3_X1   g468(.A1(new_n668), .A2(KEYINPUT102), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT102), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  OAI221_X1 g470(.A(new_n665), .B1(new_n666), .B2(new_n668), .C1(new_n670), .C2(new_n671), .ZN(G1325gat));
  NOR2_X1   g471(.A1(new_n457), .A2(new_n458), .ZN(new_n673));
  AOI21_X1  g472(.A(G15gat), .B1(new_n663), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT103), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n663), .A2(G15gat), .A3(new_n465), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n456), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n630), .ZN(new_n681));
  INV_X1    g480(.A(new_n659), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n571), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n487), .A2(KEYINPUT86), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n490), .A2(new_n496), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n513), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n463), .A2(new_n464), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n455), .B2(new_n366), .ZN(new_n691));
  OAI211_X1 g490(.A(KEYINPUT104), .B(new_n456), .C1(new_n518), .C2(new_n447), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n460), .A2(KEYINPUT35), .ZN(new_n694));
  INV_X1    g493(.A(new_n442), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n693), .A2(KEYINPUT105), .A3(new_n696), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n606), .A2(KEYINPUT44), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT44), .B1(new_n520), .B2(new_n606), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n685), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n518), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n520), .A2(new_n606), .A3(new_n685), .ZN(new_n708));
  INV_X1    g507(.A(G29gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n518), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT45), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n713), .A3(new_n396), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT106), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n705), .B2(new_n397), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n716), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(G1329gat));
  XOR2_X1   g519(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n721));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n704), .B2(new_n465), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(KEYINPUT108), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n683), .A2(G43gat), .A3(new_n606), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n572), .A2(new_n673), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT109), .Z(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n721), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n724), .A2(KEYINPUT47), .A3(new_n727), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n705), .A2(new_n366), .ZN(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n708), .A2(new_n736), .A3(new_n456), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n738), .B1(new_n735), .B2(new_n736), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OAI221_X1 g540(.A(new_n738), .B1(new_n734), .B2(KEYINPUT48), .C1(new_n735), .C2(new_n736), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n699), .A2(new_n700), .ZN(new_n744));
  NOR4_X1   g543(.A1(new_n744), .A2(new_n570), .A3(new_n631), .A4(new_n682), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n518), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g546(.A(new_n397), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT111), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n753), .B(new_n754), .ZN(G1333gat));
  NAND2_X1  g554(.A1(new_n745), .A2(new_n465), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n457), .A2(new_n458), .A3(G71gat), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n756), .A2(G71gat), .B1(new_n745), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n456), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n630), .A2(new_n570), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n682), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n766));
  INV_X1    g565(.A(new_n703), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n582), .B1(new_n768), .B2(new_n706), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n606), .B1(new_n693), .B2(new_n696), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n764), .B1(new_n770), .B2(KEYINPUT113), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n691), .A2(new_n692), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n461), .B1(new_n773), .B2(new_n514), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n606), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT51), .B1(new_n771), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR3_X1    g577(.A1(new_n706), .A2(new_n682), .A3(new_n582), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n769), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  OAI211_X1 g579(.A(new_n396), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n682), .A2(G92gat), .A3(new_n397), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n697), .A2(KEYINPUT113), .A3(new_n605), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n763), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n770), .A2(KEYINPUT113), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n775), .A3(KEYINPUT51), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n784), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n782), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n783), .B1(new_n776), .B2(new_n777), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT114), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT52), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n781), .B2(G92gat), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT115), .B1(new_n797), .B2(new_n794), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n797), .A2(KEYINPUT115), .A3(new_n794), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n768), .B2(new_n689), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n673), .A2(new_n659), .A3(new_n579), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(new_n778), .B2(new_n802), .ZN(G1338gat));
  NOR3_X1   g602(.A1(new_n682), .A2(G106gat), .A3(new_n366), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n776), .B2(new_n777), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT117), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807));
  INV_X1    g606(.A(new_n765), .ZN(new_n808));
  AOI211_X1 g607(.A(new_n366), .B(new_n808), .C1(new_n702), .C2(new_n703), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n809), .B2(new_n580), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n811), .B(new_n804), .C1(new_n776), .C2(new_n777), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n456), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT116), .A3(G106gat), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n806), .A2(new_n810), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n816));
  XNOR2_X1  g615(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n805), .B(new_n817), .C1(new_n580), .C2(new_n809), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n634), .B1(new_n644), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n642), .A2(new_n643), .A3(new_n637), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n650), .A3(KEYINPUT54), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT55), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  INV_X1    g624(.A(new_n654), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n570), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n552), .A2(new_n553), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OR3_X1    g631(.A1(new_n552), .A2(new_n830), .A3(new_n553), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n561), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n659), .A2(new_n567), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n605), .B1(new_n828), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n836), .A2(new_n567), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n827), .A3(new_n605), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n681), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n660), .A2(new_n571), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n518), .A3(new_n397), .A4(new_n459), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n571), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n706), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  INV_X1    g646(.A(new_n399), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n571), .A2(new_n216), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(G1340gat));
  NOR3_X1   g650(.A1(new_n845), .A2(new_n208), .A3(new_n682), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n847), .A2(new_n848), .A3(new_n659), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n208), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n845), .B2(new_n681), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n630), .A2(new_n221), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n849), .B2(new_n856), .ZN(G1342gat));
  NOR3_X1   g656(.A1(new_n606), .A2(G134gat), .A3(new_n396), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n847), .A2(new_n459), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT120), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n863));
  OAI21_X1  g662(.A(G134gat), .B1(new_n845), .B2(new_n606), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(G1343gat));
  NOR3_X1   g664(.A1(new_n465), .A2(new_n706), .A3(new_n396), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n366), .B1(new_n842), .B2(new_n843), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(KEYINPUT57), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G141gat), .B1(new_n871), .B2(new_n571), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n571), .A2(G141gat), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n465), .A2(new_n366), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n847), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT121), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(KEYINPUT121), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n878), .A2(new_n397), .A3(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n872), .B(new_n873), .C1(new_n875), .C2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n847), .A2(new_n397), .A3(new_n876), .A4(new_n874), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n872), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n883), .B2(new_n873), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(G148gat), .C1(new_n871), .C2(new_n682), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n888), .B1(new_n838), .B2(new_n841), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n839), .A2(new_n659), .B1(new_n827), .B2(new_n570), .ZN(new_n890));
  OAI211_X1 g689(.A(KEYINPUT122), .B(new_n840), .C1(new_n890), .C2(new_n605), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n891), .A3(new_n681), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n366), .B1(new_n892), .B2(new_n843), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n868), .B1(new_n893), .B2(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n866), .A2(new_n659), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n887), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n885), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n898), .A2(KEYINPUT123), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n897), .A2(new_n900), .A3(new_n885), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n886), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n880), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n887), .A3(new_n659), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1345gat));
  OAI21_X1  g704(.A(G155gat), .B1(new_n871), .B2(new_n681), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n681), .A2(G155gat), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n880), .B2(new_n908), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT124), .ZN(G1346gat));
  NOR3_X1   g709(.A1(new_n871), .A2(new_n600), .A3(new_n606), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n903), .A2(new_n605), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n600), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n518), .A2(new_n397), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n844), .A2(new_n459), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n571), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(new_n253), .ZN(G1348gat));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n682), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(new_n254), .ZN(G1349gat));
  INV_X1    g718(.A(new_n915), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n277), .A2(G183gat), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n279), .A4(new_n630), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G183gat), .B1(new_n915), .B2(new_n681), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT60), .ZN(G1350gat));
  OAI22_X1  g727(.A1(new_n915), .A2(new_n606), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1351gat));
  AND2_X1   g730(.A1(new_n914), .A2(new_n689), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n867), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n570), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n894), .A2(new_n932), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n570), .A2(G197gat), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(G1352gat));
  INV_X1    g736(.A(G204gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n933), .A2(new_n938), .A3(new_n659), .ZN(new_n939));
  AND2_X1   g738(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n940));
  NOR2_X1   g739(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n935), .A2(new_n659), .ZN(new_n943));
  OAI221_X1 g742(.A(new_n942), .B1(new_n940), .B2(new_n939), .C1(new_n943), .C2(new_n938), .ZN(G1353gat));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n933), .A2(new_n945), .A3(new_n630), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n894), .A2(new_n630), .A3(new_n932), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n947), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT63), .B1(new_n947), .B2(G211gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n946), .B(KEYINPUT127), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n933), .A2(new_n955), .A3(new_n605), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n935), .A2(new_n605), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n955), .ZN(G1355gat));
endmodule


