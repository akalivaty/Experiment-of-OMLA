

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788;

  OR2_X1 U369 ( .A1(n707), .A2(n706), .ZN(n540) );
  XNOR2_X1 U370 ( .A(n777), .B(G146), .ZN(n446) );
  INV_X2 U371 ( .A(G953), .ZN(n780) );
  XNOR2_X1 U372 ( .A(n544), .B(KEYINPUT42), .ZN(n596) );
  XNOR2_X2 U373 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X2 U374 ( .A(G125), .B(G146), .ZN(n470) );
  XNOR2_X2 U375 ( .A(n586), .B(n538), .ZN(n707) );
  XNOR2_X2 U376 ( .A(G128), .B(KEYINPUT82), .ZN(n431) );
  NOR2_X1 U377 ( .A1(n617), .A2(n713), .ZN(n618) );
  NAND2_X1 U378 ( .A1(n570), .A2(n569), .ZN(n758) );
  XNOR2_X1 U379 ( .A(n558), .B(KEYINPUT1), .ZN(n617) );
  XNOR2_X1 U380 ( .A(n446), .B(n439), .ZN(n684) );
  OR2_X1 U381 ( .A1(n696), .A2(KEYINPUT44), .ZN(n625) );
  XNOR2_X1 U382 ( .A(n628), .B(n627), .ZN(n757) );
  AND2_X1 U383 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U384 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U385 ( .A(n618), .B(KEYINPUT75), .ZN(n626) );
  INV_X1 U386 ( .A(n555), .ZN(n716) );
  OR2_X1 U387 ( .A1(n684), .A2(n428), .ZN(n427) );
  NAND2_X1 U388 ( .A1(n684), .A2(n424), .ZN(n423) );
  XNOR2_X1 U389 ( .A(n382), .B(n381), .ZN(n772) );
  XNOR2_X1 U390 ( .A(n442), .B(G110), .ZN(n382) );
  XNOR2_X1 U391 ( .A(KEYINPUT80), .B(KEYINPUT17), .ZN(n474) );
  XNOR2_X1 U392 ( .A(KEYINPUT18), .B(KEYINPUT79), .ZN(n469) );
  XNOR2_X1 U393 ( .A(KEYINPUT76), .B(G101), .ZN(n381) );
  XNOR2_X1 U394 ( .A(G113), .B(KEYINPUT68), .ZN(n400) );
  XNOR2_X1 U395 ( .A(G107), .B(G104), .ZN(n442) );
  BUF_X1 U396 ( .A(n660), .Z(n347) );
  INV_X1 U397 ( .A(n651), .ZN(n348) );
  XNOR2_X1 U398 ( .A(n371), .B(KEYINPUT32), .ZN(n660) );
  XNOR2_X1 U399 ( .A(n375), .B(n365), .ZN(n642) );
  AND2_X2 U400 ( .A1(n653), .A2(n700), .ZN(n349) );
  AND2_X2 U401 ( .A1(n653), .A2(n700), .ZN(n689) );
  NAND2_X1 U402 ( .A1(n400), .A2(n399), .ZN(n352) );
  NAND2_X1 U403 ( .A1(n350), .A2(n351), .ZN(n353) );
  NAND2_X1 U404 ( .A1(n352), .A2(n353), .ZN(n433) );
  INV_X1 U405 ( .A(n400), .ZN(n350) );
  INV_X1 U406 ( .A(n399), .ZN(n351) );
  XNOR2_X2 U407 ( .A(n354), .B(n355), .ZN(n586) );
  NOR2_X1 U408 ( .A1(n675), .A2(n637), .ZN(n354) );
  XOR2_X1 U409 ( .A(n486), .B(n485), .Z(n355) );
  AND2_X1 U410 ( .A1(n567), .A2(n568), .ZN(n752) );
  XNOR2_X1 U411 ( .A(n527), .B(KEYINPUT22), .ZN(n554) );
  XNOR2_X2 U412 ( .A(n472), .B(G134), .ZN(n505) );
  XNOR2_X1 U413 ( .A(n475), .B(G137), .ZN(n429) );
  AND2_X1 U414 ( .A1(n420), .A2(n417), .ZN(n416) );
  NOR2_X1 U415 ( .A1(n419), .A2(n418), .ZN(n417) );
  NAND2_X1 U416 ( .A1(n412), .A2(n421), .ZN(n420) );
  NOR2_X1 U417 ( .A1(n582), .A2(KEYINPUT30), .ZN(n418) );
  NOR2_X1 U418 ( .A1(n415), .A2(KEYINPUT30), .ZN(n414) );
  INV_X1 U419 ( .A(n423), .ZN(n415) );
  INV_X1 U420 ( .A(KEYINPUT66), .ZN(n367) );
  NOR2_X1 U421 ( .A1(n533), .A2(n716), .ZN(n368) );
  NAND2_X1 U422 ( .A1(n717), .A2(n366), .ZN(n557) );
  AND2_X1 U423 ( .A1(n702), .A2(n532), .ZN(n366) );
  INV_X1 U424 ( .A(G143), .ZN(n430) );
  AND2_X2 U425 ( .A1(n427), .A2(n426), .ZN(n425) );
  NAND2_X1 U426 ( .A1(n441), .A2(G902), .ZN(n426) );
  XNOR2_X1 U427 ( .A(G119), .B(G116), .ZN(n432) );
  XNOR2_X1 U428 ( .A(G107), .B(G116), .ZN(n500) );
  AND2_X1 U429 ( .A1(n406), .A2(n357), .ZN(n405) );
  NAND2_X1 U430 ( .A1(n404), .A2(n361), .ZN(n407) );
  NOR2_X1 U431 ( .A1(n585), .A2(n584), .ZN(n603) );
  NOR2_X2 U432 ( .A1(n554), .A2(n716), .ZN(n372) );
  NAND2_X1 U433 ( .A1(n582), .A2(KEYINPUT30), .ZN(n422) );
  XNOR2_X1 U434 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n475) );
  INV_X1 U435 ( .A(n425), .ZN(n412) );
  INV_X1 U436 ( .A(n422), .ZN(n421) );
  NOR2_X1 U437 ( .A1(n423), .A2(n422), .ZN(n419) );
  NAND2_X1 U438 ( .A1(n401), .A2(n610), .ZN(n648) );
  INV_X1 U439 ( .A(KEYINPUT88), .ZN(n380) );
  XNOR2_X1 U440 ( .A(G128), .B(G119), .ZN(n449) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n498) );
  XNOR2_X1 U442 ( .A(G143), .B(G122), .ZN(n514) );
  XOR2_X1 U443 ( .A(G113), .B(G104), .Z(n515) );
  XNOR2_X1 U444 ( .A(n772), .B(KEYINPUT70), .ZN(n483) );
  INV_X1 U445 ( .A(KEYINPUT39), .ZN(n411) );
  XNOR2_X1 U446 ( .A(n525), .B(KEYINPUT21), .ZN(n717) );
  AND2_X1 U447 ( .A1(n524), .A2(G221), .ZN(n525) );
  NOR2_X1 U448 ( .A1(n697), .A2(n638), .ZN(n641) );
  NAND2_X1 U449 ( .A1(n707), .A2(n411), .ZN(n409) );
  AND2_X1 U450 ( .A1(n385), .A2(n391), .ZN(n384) );
  AND2_X1 U451 ( .A1(n389), .A2(n387), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n562), .B(KEYINPUT78), .ZN(n592) );
  AND2_X1 U453 ( .A1(n537), .A2(n547), .ZN(n568) );
  XNOR2_X1 U454 ( .A(n481), .B(n438), .ZN(n439) );
  XNOR2_X1 U455 ( .A(n437), .B(n358), .ZN(n438) );
  XNOR2_X1 U456 ( .A(KEYINPUT16), .B(G122), .ZN(n479) );
  XNOR2_X1 U457 ( .A(n507), .B(n506), .ZN(n690) );
  NAND2_X1 U458 ( .A1(n656), .A2(G953), .ZN(n692) );
  XNOR2_X1 U459 ( .A(n595), .B(n594), .ZN(n787) );
  NAND2_X1 U460 ( .A1(n405), .A2(n407), .ZN(n595) );
  AND2_X1 U461 ( .A1(n589), .A2(n612), .ZN(n761) );
  NAND2_X1 U462 ( .A1(n372), .A2(n356), .ZN(n371) );
  XNOR2_X1 U463 ( .A(n370), .B(n369), .ZN(n613) );
  INV_X1 U464 ( .A(KEYINPUT105), .ZN(n369) );
  NAND2_X1 U465 ( .A1(n372), .A2(n362), .ZN(n370) );
  AND2_X1 U466 ( .A1(n359), .A2(n612), .ZN(n356) );
  AND2_X1 U467 ( .A1(n410), .A2(n409), .ZN(n357) );
  XOR2_X1 U468 ( .A(n436), .B(n435), .Z(n358) );
  XOR2_X1 U469 ( .A(n619), .B(KEYINPUT81), .Z(n359) );
  AND2_X1 U470 ( .A1(n708), .A2(n717), .ZN(n360) );
  NOR2_X1 U471 ( .A1(n707), .A2(n411), .ZN(n361) );
  NOR2_X1 U472 ( .A1(n720), .A2(n612), .ZN(n362) );
  XOR2_X1 U473 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n363) );
  XOR2_X1 U474 ( .A(n496), .B(KEYINPUT0), .Z(n364) );
  INV_X1 U475 ( .A(G902), .ZN(n520) );
  XNOR2_X1 U476 ( .A(n636), .B(KEYINPUT45), .ZN(n365) );
  INV_X1 U477 ( .A(n755), .ZN(n410) );
  XNOR2_X1 U478 ( .A(G902), .B(KEYINPUT15), .ZN(n643) );
  NAND2_X1 U479 ( .A1(n376), .A2(n379), .ZN(n375) );
  NAND2_X1 U480 ( .A1(n616), .A2(n615), .ZN(n378) );
  NAND2_X1 U481 ( .A1(n378), .A2(n377), .ZN(n376) );
  INV_X1 U482 ( .A(n624), .ZN(n616) );
  NAND2_X2 U483 ( .A1(n425), .A2(n423), .ZN(n720) );
  XNOR2_X2 U484 ( .A(n614), .B(KEYINPUT89), .ZN(n624) );
  NAND2_X1 U485 ( .A1(n586), .A2(n582), .ZN(n374) );
  XNOR2_X1 U486 ( .A(n368), .B(n367), .ZN(n585) );
  XNOR2_X1 U487 ( .A(n402), .B(n600), .ZN(n401) );
  NAND2_X1 U488 ( .A1(n660), .A2(n613), .ZN(n614) );
  XNOR2_X2 U489 ( .A(n373), .B(n364), .ZN(n526) );
  NAND2_X2 U490 ( .A1(n567), .A2(n495), .ZN(n373) );
  XNOR2_X2 U491 ( .A(n374), .B(KEYINPUT19), .ZN(n567) );
  NAND2_X1 U492 ( .A1(n348), .A2(n644), .ZN(n645) );
  NAND2_X1 U493 ( .A1(n348), .A2(n780), .ZN(n770) );
  NAND2_X1 U494 ( .A1(n624), .A2(n625), .ZN(n377) );
  XNOR2_X1 U495 ( .A(n635), .B(n380), .ZN(n379) );
  NAND2_X1 U496 ( .A1(n626), .A2(n363), .ZN(n396) );
  NAND2_X1 U497 ( .A1(n394), .A2(n391), .ZN(n703) );
  NAND2_X1 U498 ( .A1(n386), .A2(n383), .ZN(n622) );
  NAND2_X1 U499 ( .A1(n384), .A2(n394), .ZN(n383) );
  NOR2_X1 U500 ( .A1(n545), .A2(n620), .ZN(n385) );
  NAND2_X1 U501 ( .A1(n388), .A2(n620), .ZN(n387) );
  NAND2_X1 U502 ( .A1(n526), .A2(n391), .ZN(n388) );
  NAND2_X1 U503 ( .A1(n390), .A2(n620), .ZN(n389) );
  INV_X1 U504 ( .A(n394), .ZN(n390) );
  NOR2_X1 U505 ( .A1(n619), .A2(n363), .ZN(n392) );
  INV_X1 U506 ( .A(n626), .ZN(n393) );
  NAND2_X1 U507 ( .A1(n619), .A2(n363), .ZN(n395) );
  XNOR2_X1 U508 ( .A(n398), .B(n397), .ZN(n675) );
  INV_X1 U509 ( .A(n483), .ZN(n397) );
  XNOR2_X1 U510 ( .A(n771), .B(n482), .ZN(n398) );
  INV_X1 U511 ( .A(n526), .ZN(n545) );
  XNOR2_X2 U512 ( .A(n481), .B(n480), .ZN(n771) );
  NAND2_X1 U513 ( .A1(n403), .A2(n599), .ZN(n402) );
  XNOR2_X1 U514 ( .A(n598), .B(n597), .ZN(n403) );
  NAND2_X1 U515 ( .A1(n592), .A2(n411), .ZN(n406) );
  AND2_X1 U516 ( .A1(n406), .A2(n409), .ZN(n408) );
  INV_X1 U517 ( .A(n592), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n408), .A2(n407), .ZN(n602) );
  NAND2_X1 U519 ( .A1(n416), .A2(n413), .ZN(n560) );
  NAND2_X1 U520 ( .A1(n425), .A2(n414), .ZN(n413) );
  NOR2_X1 U521 ( .A1(n441), .A2(G902), .ZN(n424) );
  INV_X1 U522 ( .A(n441), .ZN(n428) );
  XNOR2_X2 U523 ( .A(n505), .B(n429), .ZN(n777) );
  XNOR2_X2 U524 ( .A(n431), .B(n430), .ZN(n472) );
  AND2_X1 U525 ( .A1(n779), .A2(n637), .ZN(n644) );
  XNOR2_X1 U526 ( .A(n446), .B(n445), .ZN(n669) );
  INV_X1 U527 ( .A(KEYINPUT46), .ZN(n597) );
  INV_X1 U528 ( .A(KEYINPUT23), .ZN(n451) );
  XNOR2_X1 U529 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U530 ( .A(n483), .B(n444), .ZN(n445) );
  XNOR2_X1 U531 ( .A(n454), .B(n453), .ZN(n455) );
  BUF_X1 U532 ( .A(n613), .Z(n556) );
  XNOR2_X2 U533 ( .A(n433), .B(n432), .ZN(n481) );
  NOR2_X1 U534 ( .A1(G953), .A2(G237), .ZN(n434) );
  XOR2_X1 U535 ( .A(KEYINPUT77), .B(n434), .Z(n509) );
  NAND2_X1 U536 ( .A1(n509), .A2(G210), .ZN(n437) );
  XOR2_X1 U537 ( .A(KEYINPUT99), .B(KEYINPUT5), .Z(n436) );
  XNOR2_X1 U538 ( .A(G101), .B(G131), .ZN(n435) );
  INV_X1 U539 ( .A(KEYINPUT71), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n440), .B(G472), .ZN(n441) );
  XNOR2_X1 U541 ( .A(n720), .B(KEYINPUT6), .ZN(n619) );
  XOR2_X1 U542 ( .A(G140), .B(G131), .Z(n512) );
  NAND2_X1 U543 ( .A1(G227), .A2(n780), .ZN(n443) );
  XNOR2_X1 U544 ( .A(n512), .B(n443), .ZN(n444) );
  NAND2_X1 U545 ( .A1(n669), .A2(n520), .ZN(n448) );
  INV_X1 U546 ( .A(G469), .ZN(n447) );
  XNOR2_X2 U547 ( .A(n448), .B(n447), .ZN(n558) );
  INV_X1 U548 ( .A(n617), .ZN(n612) );
  INV_X1 U549 ( .A(n612), .ZN(n714) );
  XOR2_X1 U550 ( .A(KEYINPUT84), .B(G137), .Z(n450) );
  XNOR2_X1 U551 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U552 ( .A(G110), .B(G140), .ZN(n452) );
  XNOR2_X1 U553 ( .A(n470), .B(KEYINPUT10), .ZN(n510) );
  XNOR2_X1 U554 ( .A(n455), .B(n510), .ZN(n460) );
  NAND2_X1 U555 ( .A1(G234), .A2(n780), .ZN(n456) );
  XOR2_X1 U556 ( .A(KEYINPUT8), .B(n456), .Z(n502) );
  NAND2_X1 U557 ( .A1(n502), .A2(G221), .ZN(n458) );
  XNOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT24), .ZN(n457) );
  XNOR2_X1 U559 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U560 ( .A(n460), .B(n459), .ZN(n655) );
  NAND2_X1 U561 ( .A1(n655), .A2(n520), .ZN(n467) );
  XOR2_X1 U562 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n462) );
  NAND2_X1 U563 ( .A1(G234), .A2(n643), .ZN(n461) );
  XNOR2_X1 U564 ( .A(n461), .B(n462), .ZN(n463) );
  XNOR2_X1 U565 ( .A(KEYINPUT96), .B(n463), .ZN(n524) );
  NAND2_X1 U566 ( .A1(G217), .A2(n524), .ZN(n464) );
  XNOR2_X1 U567 ( .A(KEYINPUT98), .B(n464), .ZN(n465) );
  XNOR2_X1 U568 ( .A(n465), .B(KEYINPUT25), .ZN(n466) );
  XNOR2_X1 U569 ( .A(n467), .B(n466), .ZN(n555) );
  AND2_X1 U570 ( .A1(n714), .A2(n716), .ZN(n468) );
  NAND2_X1 U571 ( .A1(n619), .A2(n468), .ZN(n528) );
  XNOR2_X1 U572 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n472), .B(n471), .ZN(n478) );
  NAND2_X1 U574 ( .A1(n780), .A2(G224), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U576 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U577 ( .A(n478), .B(n477), .ZN(n482) );
  XNOR2_X1 U578 ( .A(n479), .B(KEYINPUT72), .ZN(n480) );
  INV_X1 U579 ( .A(n643), .ZN(n637) );
  INV_X1 U580 ( .A(G237), .ZN(n484) );
  NAND2_X1 U581 ( .A1(n520), .A2(n484), .ZN(n487) );
  NAND2_X1 U582 ( .A1(n487), .A2(G210), .ZN(n486) );
  INV_X1 U583 ( .A(KEYINPUT92), .ZN(n485) );
  NAND2_X1 U584 ( .A1(n487), .A2(G214), .ZN(n582) );
  NAND2_X1 U585 ( .A1(G237), .A2(G234), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n488), .B(KEYINPUT14), .ZN(n489) );
  XOR2_X1 U587 ( .A(KEYINPUT73), .B(n489), .Z(n702) );
  NAND2_X1 U588 ( .A1(G952), .A2(n780), .ZN(n530) );
  INV_X1 U589 ( .A(n530), .ZN(n490) );
  NAND2_X1 U590 ( .A1(n702), .A2(n490), .ZN(n494) );
  XNOR2_X1 U591 ( .A(KEYINPUT93), .B(G898), .ZN(n767) );
  NAND2_X1 U592 ( .A1(G953), .A2(n767), .ZN(n773) );
  NOR2_X1 U593 ( .A1(n520), .A2(n773), .ZN(n491) );
  NAND2_X1 U594 ( .A1(n491), .A2(n702), .ZN(n492) );
  XNOR2_X1 U595 ( .A(n492), .B(KEYINPUT94), .ZN(n493) );
  NAND2_X1 U596 ( .A1(n494), .A2(n493), .ZN(n495) );
  INV_X1 U597 ( .A(KEYINPUT65), .ZN(n496) );
  XNOR2_X1 U598 ( .A(G122), .B(KEYINPUT7), .ZN(n497) );
  XNOR2_X1 U599 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U600 ( .A(n499), .B(KEYINPUT102), .Z(n501) );
  XNOR2_X1 U601 ( .A(n501), .B(n500), .ZN(n504) );
  NAND2_X1 U602 ( .A1(n502), .A2(G217), .ZN(n503) );
  XNOR2_X1 U603 ( .A(n504), .B(n503), .ZN(n507) );
  INV_X1 U604 ( .A(n505), .ZN(n506) );
  NAND2_X1 U605 ( .A1(n690), .A2(n520), .ZN(n508) );
  XNOR2_X1 U606 ( .A(n508), .B(G478), .ZN(n570) );
  INV_X1 U607 ( .A(n570), .ZN(n523) );
  NAND2_X1 U608 ( .A1(n509), .A2(G214), .ZN(n513) );
  INV_X1 U609 ( .A(n510), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n512), .B(n511), .ZN(n778) );
  XNOR2_X1 U611 ( .A(n513), .B(n778), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U613 ( .A(n516), .B(KEYINPUT12), .Z(n517) );
  XNOR2_X1 U614 ( .A(n517), .B(KEYINPUT11), .ZN(n518) );
  XNOR2_X1 U615 ( .A(n519), .B(n518), .ZN(n662) );
  NAND2_X1 U616 ( .A1(n662), .A2(n520), .ZN(n522) );
  XNOR2_X1 U617 ( .A(KEYINPUT13), .B(G475), .ZN(n521) );
  XNOR2_X1 U618 ( .A(n522), .B(n521), .ZN(n569) );
  AND2_X1 U619 ( .A1(n523), .A2(n569), .ZN(n708) );
  NAND2_X1 U620 ( .A1(n526), .A2(n360), .ZN(n527) );
  OR2_X1 U621 ( .A1(n554), .A2(n528), .ZN(n631) );
  XNOR2_X1 U622 ( .A(n631), .B(G101), .ZN(G3) );
  INV_X1 U623 ( .A(n720), .ZN(n534) );
  NOR2_X1 U624 ( .A1(G900), .A2(n780), .ZN(n529) );
  NAND2_X1 U625 ( .A1(G902), .A2(n529), .ZN(n531) );
  NAND2_X1 U626 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U627 ( .A(n557), .B(KEYINPUT67), .Z(n533) );
  OR2_X1 U628 ( .A1(n534), .A2(n585), .ZN(n536) );
  XOR2_X1 U629 ( .A(KEYINPUT28), .B(KEYINPUT110), .Z(n535) );
  XNOR2_X1 U630 ( .A(n536), .B(n535), .ZN(n537) );
  INV_X1 U631 ( .A(n558), .ZN(n547) );
  XNOR2_X1 U632 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n538) );
  INV_X1 U633 ( .A(n582), .ZN(n706) );
  INV_X1 U634 ( .A(KEYINPUT112), .ZN(n539) );
  XNOR2_X1 U635 ( .A(n540), .B(n539), .ZN(n705) );
  NAND2_X1 U636 ( .A1(n705), .A2(n708), .ZN(n543) );
  INV_X1 U637 ( .A(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U638 ( .A(n541), .B(KEYINPUT41), .ZN(n542) );
  XNOR2_X1 U639 ( .A(n543), .B(n542), .ZN(n727) );
  NAND2_X1 U640 ( .A1(n568), .A2(n727), .ZN(n544) );
  XNOR2_X1 U641 ( .A(n596), .B(G137), .ZN(G39) );
  INV_X1 U642 ( .A(n717), .ZN(n546) );
  OR2_X1 U643 ( .A1(n555), .A2(n546), .ZN(n713) );
  INV_X1 U644 ( .A(n713), .ZN(n548) );
  NAND2_X1 U645 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U646 ( .A1(n720), .A2(n549), .ZN(n550) );
  NOR2_X1 U647 ( .A1(n545), .A2(n550), .ZN(n552) );
  INV_X1 U648 ( .A(KEYINPUT100), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n552), .B(n551), .ZN(n743) );
  OR2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n755) );
  NOR2_X1 U651 ( .A1(n743), .A2(n755), .ZN(n553) );
  XOR2_X1 U652 ( .A(G104), .B(n553), .Z(G6) );
  XNOR2_X1 U653 ( .A(n556), .B(G110), .ZN(G12) );
  NOR2_X1 U654 ( .A1(n558), .A2(n557), .ZN(n559) );
  AND2_X1 U655 ( .A1(n559), .A2(n716), .ZN(n561) );
  NAND2_X1 U656 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U657 ( .A(n586), .ZN(n606) );
  NOR2_X1 U658 ( .A1(n592), .A2(n606), .ZN(n564) );
  INV_X1 U659 ( .A(KEYINPUT109), .ZN(n563) );
  XNOR2_X1 U660 ( .A(n564), .B(n563), .ZN(n566) );
  INV_X1 U661 ( .A(n569), .ZN(n565) );
  AND2_X1 U662 ( .A1(n570), .A2(n565), .ZN(n621) );
  AND2_X1 U663 ( .A1(n566), .A2(n621), .ZN(n751) );
  XNOR2_X1 U664 ( .A(n758), .B(KEYINPUT104), .ZN(n601) );
  AND2_X1 U665 ( .A1(n601), .A2(n755), .ZN(n704) );
  INV_X1 U666 ( .A(n704), .ZN(n571) );
  OR2_X1 U667 ( .A1(KEYINPUT83), .A2(n571), .ZN(n572) );
  NAND2_X1 U668 ( .A1(n752), .A2(n572), .ZN(n574) );
  INV_X1 U669 ( .A(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U670 ( .A1(n574), .A2(n573), .ZN(n577) );
  NOR2_X1 U671 ( .A1(KEYINPUT47), .A2(KEYINPUT83), .ZN(n575) );
  OR2_X1 U672 ( .A1(n704), .A2(n575), .ZN(n576) );
  NAND2_X1 U673 ( .A1(n577), .A2(n576), .ZN(n580) );
  INV_X1 U674 ( .A(n752), .ZN(n578) );
  NAND2_X1 U675 ( .A1(n578), .A2(KEYINPUT47), .ZN(n579) );
  NAND2_X1 U676 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U677 ( .A1(n751), .A2(n581), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n755), .A2(n619), .ZN(n583) );
  NAND2_X1 U679 ( .A1(n583), .A2(n582), .ZN(n584) );
  AND2_X1 U680 ( .A1(n586), .A2(n603), .ZN(n588) );
  XNOR2_X1 U681 ( .A(KEYINPUT36), .B(KEYINPUT114), .ZN(n587) );
  XNOR2_X1 U682 ( .A(n588), .B(n587), .ZN(n589) );
  INV_X1 U683 ( .A(n761), .ZN(n590) );
  AND2_X1 U684 ( .A1(n591), .A2(n590), .ZN(n599) );
  INV_X1 U685 ( .A(KEYINPUT111), .ZN(n593) );
  XNOR2_X1 U686 ( .A(n593), .B(KEYINPUT40), .ZN(n594) );
  NAND2_X1 U687 ( .A1(n787), .A2(n596), .ZN(n598) );
  INV_X1 U688 ( .A(KEYINPUT48), .ZN(n600) );
  OR2_X1 U689 ( .A1(n602), .A2(n601), .ZN(n763) );
  XOR2_X1 U690 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n605) );
  NAND2_X1 U691 ( .A1(n603), .A2(n714), .ZN(n604) );
  XNOR2_X1 U692 ( .A(n605), .B(n604), .ZN(n607) );
  AND2_X1 U693 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U694 ( .A(KEYINPUT108), .ZN(n608) );
  XNOR2_X1 U695 ( .A(n609), .B(n608), .ZN(n788) );
  AND2_X1 U696 ( .A1(n763), .A2(n788), .ZN(n610) );
  INV_X1 U697 ( .A(KEYINPUT86), .ZN(n611) );
  XNOR2_X2 U698 ( .A(n648), .B(n611), .ZN(n779) );
  INV_X1 U699 ( .A(KEYINPUT44), .ZN(n615) );
  INV_X1 U700 ( .A(KEYINPUT34), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X2 U702 ( .A(n623), .B(KEYINPUT35), .ZN(n696) );
  NAND2_X1 U703 ( .A1(n696), .A2(KEYINPUT44), .ZN(n634) );
  NAND2_X1 U704 ( .A1(n720), .A2(n393), .ZN(n723) );
  OR2_X1 U705 ( .A1(n723), .A2(n545), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n757), .A2(n743), .ZN(n630) );
  XNOR2_X1 U708 ( .A(n704), .B(KEYINPUT83), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n632) );
  AND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  INV_X1 U712 ( .A(KEYINPUT87), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n779), .A2(n642), .ZN(n697) );
  INV_X1 U714 ( .A(n637), .ZN(n639) );
  OR2_X1 U715 ( .A1(KEYINPUT85), .A2(n639), .ZN(n638) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n698) );
  NOR2_X1 U717 ( .A1(n639), .A2(n698), .ZN(n640) );
  NOR2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n647) );
  INV_X1 U719 ( .A(n642), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n645), .A2(KEYINPUT85), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n653) );
  BUF_X1 U722 ( .A(n648), .Z(n649) );
  INV_X1 U723 ( .A(n649), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n650), .A2(KEYINPUT2), .ZN(n652) );
  OR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n700) );
  NAND2_X1 U726 ( .A1(n349), .A2(G217), .ZN(n654) );
  XOR2_X1 U727 ( .A(n655), .B(n654), .Z(n658) );
  INV_X1 U728 ( .A(G952), .ZN(n656) );
  INV_X1 U729 ( .A(n692), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(G66) );
  XNOR2_X1 U731 ( .A(G119), .B(KEYINPUT126), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n347), .B(n659), .ZN(G21) );
  NAND2_X1 U733 ( .A1(n689), .A2(G475), .ZN(n664) );
  XNOR2_X1 U734 ( .A(KEYINPUT91), .B(KEYINPUT59), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U736 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U737 ( .A1(n665), .A2(n692), .ZN(n667) );
  XNOR2_X1 U738 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G60) );
  NAND2_X1 U740 ( .A1(n689), .A2(G469), .ZN(n671) );
  XOR2_X1 U741 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n671), .B(n670), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n672), .A2(n692), .ZN(n674) );
  INV_X1 U745 ( .A(KEYINPUT122), .ZN(n673) );
  XNOR2_X1 U746 ( .A(n674), .B(n673), .ZN(G54) );
  NAND2_X1 U747 ( .A1(n689), .A2(G210), .ZN(n680) );
  XOR2_X1 U748 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n677) );
  XNOR2_X1 U749 ( .A(KEYINPUT55), .B(KEYINPUT90), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U751 ( .A(n675), .B(n678), .ZN(n679) );
  XNOR2_X1 U752 ( .A(n680), .B(n679), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(n692), .ZN(n683) );
  INV_X1 U754 ( .A(KEYINPUT56), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n683), .B(n682), .ZN(G51) );
  NAND2_X1 U756 ( .A1(n349), .A2(G472), .ZN(n686) );
  XNOR2_X1 U757 ( .A(n684), .B(KEYINPUT62), .ZN(n685) );
  XNOR2_X1 U758 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n687), .A2(n692), .ZN(n688) );
  XNOR2_X1 U760 ( .A(n688), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U761 ( .A1(n349), .A2(G478), .ZN(n691) );
  XNOR2_X1 U762 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n695) );
  INV_X1 U764 ( .A(KEYINPUT124), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n695), .B(n694), .ZN(G63) );
  XOR2_X1 U766 ( .A(n696), .B(G122), .Z(G24) );
  BUF_X1 U767 ( .A(n697), .Z(n699) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n739) );
  NAND2_X1 U770 ( .A1(G952), .A2(n702), .ZN(n733) );
  NAND2_X1 U771 ( .A1(n705), .A2(n571), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  AND2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n703), .A2(n712), .ZN(n730) );
  NAND2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U777 ( .A(n715), .B(KEYINPUT50), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U779 ( .A(KEYINPUT49), .B(n718), .Z(n719) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n724) );
  NAND2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U783 ( .A(KEYINPUT118), .B(n725), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n726), .B(KEYINPUT51), .ZN(n728) );
  INV_X1 U785 ( .A(n727), .ZN(n735) );
  NOR2_X1 U786 ( .A1(n728), .A2(n735), .ZN(n729) );
  NOR2_X1 U787 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U788 ( .A(n731), .B(KEYINPUT52), .ZN(n732) );
  NOR2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U790 ( .A(n734), .B(KEYINPUT119), .Z(n737) );
  NOR2_X1 U791 ( .A1(n703), .A2(n735), .ZN(n736) );
  NOR2_X1 U792 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n740), .B(KEYINPUT120), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n741), .A2(G953), .ZN(n742) );
  XNOR2_X1 U796 ( .A(n742), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U797 ( .A1(n743), .A2(n758), .ZN(n745) );
  XNOR2_X1 U798 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n745), .B(n744), .ZN(n746) );
  XNOR2_X1 U800 ( .A(G107), .B(n746), .ZN(G9) );
  XOR2_X1 U801 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n749) );
  INV_X1 U802 ( .A(n758), .ZN(n747) );
  NAND2_X1 U803 ( .A1(n752), .A2(n747), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n749), .B(n748), .ZN(n750) );
  XOR2_X1 U805 ( .A(G128), .B(n750), .Z(G30) );
  XOR2_X1 U806 ( .A(G143), .B(n751), .Z(G45) );
  XNOR2_X1 U807 ( .A(G146), .B(KEYINPUT116), .ZN(n754) );
  NAND2_X1 U808 ( .A1(n752), .A2(n410), .ZN(n753) );
  XNOR2_X1 U809 ( .A(n754), .B(n753), .ZN(G48) );
  NOR2_X1 U810 ( .A1(n755), .A2(n757), .ZN(n756) );
  XOR2_X1 U811 ( .A(G113), .B(n756), .Z(G15) );
  NOR2_X1 U812 ( .A1(n758), .A2(n757), .ZN(n760) );
  XNOR2_X1 U813 ( .A(G116), .B(KEYINPUT117), .ZN(n759) );
  XNOR2_X1 U814 ( .A(n760), .B(n759), .ZN(G18) );
  XNOR2_X1 U815 ( .A(G125), .B(n761), .ZN(n762) );
  XNOR2_X1 U816 ( .A(n762), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U817 ( .A(n763), .ZN(n764) );
  XOR2_X1 U818 ( .A(G134), .B(n764), .Z(G36) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n765) );
  XOR2_X1 U820 ( .A(KEYINPUT61), .B(n765), .Z(n766) );
  NOR2_X1 U821 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U822 ( .A(n768), .B(KEYINPUT125), .ZN(n769) );
  NAND2_X1 U823 ( .A1(n770), .A2(n769), .ZN(n776) );
  XNOR2_X1 U824 ( .A(n771), .B(n772), .ZN(n774) );
  NAND2_X1 U825 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U826 ( .A(n776), .B(n775), .Z(G69) );
  XNOR2_X1 U827 ( .A(n778), .B(n777), .ZN(n782) );
  XOR2_X1 U828 ( .A(n782), .B(n779), .Z(n781) );
  NAND2_X1 U829 ( .A1(n781), .A2(n780), .ZN(n786) );
  XNOR2_X1 U830 ( .A(G227), .B(n782), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n783), .A2(G900), .ZN(n784) );
  NAND2_X1 U832 ( .A1(n784), .A2(G953), .ZN(n785) );
  NAND2_X1 U833 ( .A1(n786), .A2(n785), .ZN(G72) );
  XNOR2_X1 U834 ( .A(G131), .B(n787), .ZN(G33) );
  XNOR2_X1 U835 ( .A(G140), .B(n788), .ZN(G42) );
endmodule

