//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G221), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(G214), .B1(G237), .B2(G902), .ZN(new_n193));
  INV_X1    g007(.A(G469), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT0), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT0), .B(G128), .Z(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n195), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n201), .B2(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR3_X1    g018(.A1(new_n201), .A2(KEYINPUT3), .A3(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(G107), .ZN(new_n206));
  OAI211_X1 g020(.A(KEYINPUT79), .B(KEYINPUT3), .C1(new_n201), .C2(G107), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT4), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G101), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(G101), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n201), .A2(KEYINPUT3), .A3(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT80), .B(G101), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n216), .A3(new_n204), .A4(new_n207), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n200), .B(new_n210), .C1(new_n211), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(G104), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n201), .A2(KEYINPUT81), .A3(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G101), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT1), .B1(new_n227), .B2(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G143), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(G128), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n195), .A2(new_n238), .A3(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n226), .A2(new_n240), .A3(KEYINPUT10), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT11), .ZN(new_n242));
  INV_X1    g056(.A(G134), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n243), .B2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G131), .ZN(new_n249));
  INV_X1    g063(.A(G131), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n244), .A2(new_n246), .A3(new_n250), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n197), .B1(new_n231), .B2(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n239), .B1(new_n254), .B2(new_n195), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(new_n217), .A3(new_n225), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT10), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n219), .A2(new_n241), .A3(new_n253), .A4(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G140), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(G227), .ZN(new_n262));
  XOR2_X1   g076(.A(new_n260), .B(new_n262), .Z(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT82), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n219), .A2(new_n241), .A3(new_n258), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n252), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(KEYINPUT82), .A3(new_n263), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n197), .B1(new_n228), .B2(KEYINPUT65), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n195), .B1(new_n271), .B2(new_n233), .ZN(new_n272));
  INV_X1    g086(.A(new_n239), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n217), .A2(new_n225), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n256), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT12), .B1(new_n277), .B2(new_n252), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT12), .ZN(new_n279));
  AOI211_X1 g093(.A(new_n279), .B(new_n253), .C1(new_n276), .C2(new_n256), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n259), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n263), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n270), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT83), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n270), .A2(new_n286), .A3(new_n283), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n194), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n263), .B1(new_n268), .B2(new_n259), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n259), .B(new_n263), .C1(new_n278), .C2(new_n280), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n194), .A3(new_n188), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n194), .A2(new_n188), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n192), .B(new_n193), .C1(new_n288), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT2), .B(G113), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n306), .B1(new_n301), .B2(new_n303), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n304), .B2(new_n299), .ZN(new_n310));
  INV_X1    g124(.A(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT2), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n319), .B(new_n210), .C1(new_n211), .C2(new_n218), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n301), .B2(KEYINPUT5), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n300), .A3(KEYINPUT84), .A4(G116), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n322), .A2(G113), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n304), .A2(KEYINPUT66), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n306), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n325), .B1(new_n328), .B2(new_n323), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n226), .A2(new_n318), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G110), .B(G122), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n320), .A2(new_n330), .A3(new_n332), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n274), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n199), .A2(new_n195), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(G125), .A3(new_n198), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G224), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G953), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT6), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n345), .A3(new_n333), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n336), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n317), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT67), .B1(new_n315), .B2(new_n316), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n322), .A2(G113), .A3(new_n324), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n304), .A2(new_n323), .ZN(new_n351));
  OAI22_X1  g165(.A1(new_n348), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n226), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n329), .A2(new_n318), .A3(new_n275), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n332), .B(KEYINPUT8), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n353), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n335), .A2(new_n357), .ZN(new_n358));
  OR3_X1    g172(.A1(new_n240), .A2(KEYINPUT86), .A3(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n338), .A2(KEYINPUT86), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n340), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT7), .B1(new_n342), .B2(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n356), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n226), .B2(new_n352), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n355), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n362), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n338), .A2(new_n340), .A3(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n358), .A2(new_n363), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n347), .A2(new_n370), .A3(new_n188), .ZN(new_n371));
  OAI21_X1  g185(.A(G210), .B1(G237), .B2(G902), .ZN(new_n372));
  XOR2_X1   g186(.A(new_n372), .B(KEYINPUT87), .Z(new_n373));
  AOI21_X1  g187(.A(new_n298), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n373), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n335), .A2(new_n369), .A3(new_n357), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(new_n366), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n377), .B2(new_n363), .ZN(new_n378));
  INV_X1    g192(.A(new_n373), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n347), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n374), .B1(new_n381), .B2(new_n298), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n261), .A3(G214), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n227), .ZN(new_n386));
  NOR2_X1   g200(.A1(G237), .A2(G953), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G143), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT89), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n388), .ZN(new_n393));
  AOI21_X1  g207(.A(G143), .B1(new_n387), .B2(G214), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT18), .B(G131), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G140), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G125), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n337), .A2(G140), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G146), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n230), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n386), .A2(KEYINPUT89), .A3(new_n388), .A4(new_n389), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n392), .A2(new_n395), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n250), .B1(new_n386), .B2(new_n388), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n408), .A2(KEYINPUT18), .B1(new_n402), .B2(new_n400), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n409), .A2(KEYINPUT90), .A3(new_n392), .A4(new_n404), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G131), .B1(new_n393), .B2(new_n394), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n386), .A2(new_n250), .A3(new_n388), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n408), .A2(KEYINPUT17), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT16), .ZN(new_n418));
  OR3_X1    g232(.A1(new_n337), .A2(KEYINPUT16), .A3(G140), .ZN(new_n419));
  AOI21_X1  g233(.A(G146), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(new_n419), .A3(G146), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G113), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(new_n201), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n383), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n407), .A2(new_n410), .B1(new_n417), .B2(new_n424), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT92), .A3(new_n428), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n412), .A2(new_n414), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n399), .A2(KEYINPUT19), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n401), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n422), .B1(new_n437), .B2(G146), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n411), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n428), .B1(new_n441), .B2(KEYINPUT91), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n439), .B1(new_n407), .B2(new_n410), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n430), .A2(new_n432), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(G475), .A2(G902), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT20), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT92), .B1(new_n431), .B2(new_n428), .ZN(new_n450));
  AND4_X1   g264(.A1(KEYINPUT92), .A2(new_n411), .A3(new_n425), .A4(new_n428), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n429), .B1(new_n443), .B2(new_n444), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n411), .A2(new_n440), .A3(new_n444), .ZN(new_n453));
  OAI22_X1  g267(.A1(new_n450), .A2(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n302), .B2(G122), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT94), .A3(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n302), .A2(G122), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n462), .A2(G107), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G107), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n197), .B2(G143), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n227), .A2(KEYINPUT95), .A3(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n197), .A2(G143), .ZN(new_n471));
  AOI21_X1  g285(.A(G134), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n462), .A2(KEYINPUT14), .A3(G107), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(G134), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n227), .A2(G128), .ZN(new_n477));
  AOI211_X1 g291(.A(new_n243), .B(new_n477), .C1(new_n468), .C2(new_n469), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT13), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n471), .A2(new_n479), .A3(G134), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n478), .A2(new_n472), .A3(new_n481), .ZN(new_n482));
  AND4_X1   g296(.A1(new_n479), .A2(new_n470), .A3(G134), .A4(new_n471), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n466), .B(new_n476), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n187), .A2(G217), .A3(new_n261), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT96), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n473), .A2(new_n475), .ZN(new_n487));
  OAI22_X1  g301(.A1(new_n487), .A2(new_n474), .B1(new_n465), .B2(new_n464), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n486), .B1(new_n484), .B2(new_n488), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n188), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n431), .A2(new_n428), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n430), .B2(new_n432), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT93), .B1(new_n498), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n450), .A2(new_n451), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n500), .B(new_n188), .C1(new_n501), .C2(new_n497), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n502), .A3(G475), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n261), .A2(G952), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(G234), .B2(G237), .ZN(new_n505));
  NAND2_X1  g319(.A1(G234), .A2(G237), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(G902), .A3(G953), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT97), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g323(.A(KEYINPUT21), .B(G898), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n457), .A2(new_n496), .A3(new_n503), .A4(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n297), .A2(new_n382), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n245), .A2(KEYINPUT64), .A3(G134), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT64), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n245), .B2(G134), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n243), .A2(G137), .ZN(new_n520));
  OAI211_X1 g334(.A(G131), .B(new_n517), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n251), .B(new_n521), .C1(new_n272), .C2(new_n273), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n252), .A2(new_n200), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n328), .A2(new_n299), .B1(new_n310), .B2(new_n317), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n524), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n530), .B2(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n521), .A2(new_n251), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n237), .B2(new_n239), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n339), .A2(new_n198), .B1(new_n249), .B2(new_n251), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n319), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n525), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n531), .B2(new_n537), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n529), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n387), .A2(G210), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT68), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(KEYINPUT30), .C1(new_n533), .C2(new_n534), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n548), .A2(KEYINPUT30), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(KEYINPUT30), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n522), .A2(new_n523), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n319), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n525), .A2(new_n546), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT69), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n525), .A2(new_n557), .A3(new_n546), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT31), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n524), .B1(new_n549), .B2(new_n552), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n525), .A2(new_n557), .A3(new_n546), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .A3(new_n556), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n542), .A2(new_n547), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n566), .A2(KEYINPUT73), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT73), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n527), .B(KEYINPUT72), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n531), .A2(new_n537), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT71), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n571), .B1(new_n573), .B2(new_n539), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT31), .B1(new_n564), .B2(new_n556), .ZN(new_n575));
  AND4_X1   g389(.A1(KEYINPUT31), .A2(new_n554), .A3(new_n556), .A4(new_n558), .ZN(new_n576));
  OAI22_X1  g390(.A1(new_n574), .A2(new_n546), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n577), .B2(new_n567), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n516), .B1(new_n569), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n542), .A2(new_n547), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n565), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n568), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT29), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n554), .A2(new_n525), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n547), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n584), .B(new_n586), .C1(new_n542), .C2(new_n547), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n535), .A2(new_n525), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n526), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n571), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n547), .A2(new_n584), .ZN(new_n591));
  AOI21_X1  g405(.A(G902), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G472), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n579), .A2(new_n583), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n300), .A2(G128), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n197), .A2(G119), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT24), .B(G110), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n418), .A2(G146), .A3(new_n419), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n600), .B1(new_n601), .B2(new_n420), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n603), .B1(new_n300), .B2(G128), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT23), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT23), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n607), .A3(new_n596), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G110), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT75), .B1(new_n602), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT75), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n423), .A2(new_n612), .A3(new_n609), .A4(new_n600), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n605), .A2(new_n607), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT76), .ZN(new_n616));
  INV_X1    g430(.A(G110), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n596), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT76), .B1(new_n608), .B2(G110), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n598), .A2(new_n599), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n422), .A3(new_n402), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT22), .B(G137), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n614), .A2(new_n622), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n625), .B1(new_n614), .B2(new_n622), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n614), .A2(new_n622), .ZN(new_n630));
  INV_X1    g444(.A(new_n625), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n614), .A2(new_n622), .A3(new_n625), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n188), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT25), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G217), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(G234), .B2(new_n188), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(G902), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT77), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n639), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n629), .B2(new_n636), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT77), .ZN(new_n646));
  INV_X1    g460(.A(new_n642), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n515), .A2(new_n595), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(new_n216), .Z(G3));
  OAI21_X1  g467(.A(G472), .B1(new_n566), .B2(G902), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n569), .B2(new_n578), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n192), .B1(new_n288), .B2(new_n296), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n649), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n491), .A2(KEYINPUT99), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n484), .A2(new_n488), .ZN(new_n660));
  INV_X1    g474(.A(new_n486), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n484), .A2(new_n488), .A3(new_n486), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT33), .B1(new_n489), .B2(new_n490), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(KEYINPUT100), .B(KEYINPUT33), .C1(new_n489), .C2(new_n490), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n667), .A2(new_n672), .A3(G478), .A4(new_n188), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n492), .A2(new_n493), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n457), .A2(new_n503), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n193), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n375), .B2(new_n380), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n512), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n657), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT34), .B(G104), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G6));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n503), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n499), .A2(new_n502), .A3(KEYINPUT102), .A4(G475), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n454), .A2(new_n455), .A3(new_n447), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n455), .B1(new_n454), .B2(new_n447), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT101), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n449), .A2(new_n689), .A3(new_n456), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n684), .A2(new_n685), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n495), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n657), .A2(new_n692), .A3(new_n679), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT35), .B(G107), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  OAI21_X1  g509(.A(KEYINPUT73), .B1(new_n566), .B2(new_n568), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n577), .A2(new_n570), .A3(new_n567), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n630), .B(KEYINPUT103), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n631), .A2(KEYINPUT36), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n645), .B1(new_n701), .B2(new_n641), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n515), .A2(new_n698), .A3(new_n654), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n617), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G12));
  NAND2_X1  g521(.A1(new_n684), .A2(new_n685), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n688), .A2(new_n690), .ZN(new_n709));
  INV_X1    g523(.A(G900), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n505), .B1(new_n509), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n495), .A2(new_n708), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  AOI211_X1 g527(.A(G469), .B(G902), .C1(new_n290), .C2(new_n291), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n294), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n270), .A2(new_n286), .A3(new_n283), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n286), .B1(new_n270), .B2(new_n283), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n191), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n677), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n713), .A2(new_n595), .A3(new_n721), .A4(new_n703), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT105), .B(G128), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G30));
  XNOR2_X1  g538(.A(new_n711), .B(KEYINPUT39), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT40), .B1(new_n656), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n371), .A2(new_n373), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n379), .B1(new_n378), .B2(new_n347), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n298), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n374), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n731), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT88), .B1(new_n375), .B2(new_n380), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n733), .B1(new_n734), .B2(new_n374), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n656), .A2(new_n725), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT40), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n703), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(G472), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n559), .B1(new_n588), .B2(new_n546), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n188), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT107), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n579), .A2(new_n583), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n496), .B1(new_n457), .B2(new_n503), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n193), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n737), .A2(new_n740), .A3(new_n745), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  NAND2_X1  g563(.A1(new_n457), .A2(new_n503), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n673), .A2(new_n674), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n711), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n595), .A2(new_n721), .A3(new_n703), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  NOR3_X1   g569(.A1(new_n566), .A2(new_n516), .A3(new_n568), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n698), .B2(new_n516), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n649), .B1(new_n757), .B2(new_n594), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n194), .B1(new_n292), .B2(new_n188), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n714), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n192), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n752), .A2(new_n761), .A3(new_n678), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n513), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT41), .B(G113), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G15));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n678), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n758), .A2(new_n692), .A3(new_n513), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G116), .ZN(G18));
  AOI21_X1  g582(.A(new_n702), .B1(new_n757), .B2(new_n594), .ZN(new_n769));
  INV_X1    g583(.A(new_n514), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n766), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G119), .ZN(G21));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n654), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n645), .A2(new_n647), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n581), .B1(new_n546), .B2(new_n590), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n567), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT108), .B(G472), .C1(new_n566), .C2(G902), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n761), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n679), .A3(new_n746), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G122), .ZN(G24));
  AND4_X1   g596(.A1(new_n703), .A2(new_n774), .A3(new_n777), .A4(new_n778), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n753), .A3(new_n766), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  NOR2_X1   g599(.A1(new_n191), .A2(new_n676), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n734), .A2(new_n374), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n293), .B(new_n295), .C1(new_n284), .C2(new_n194), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n675), .A3(new_n712), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n516), .B1(new_n566), .B2(new_n568), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n594), .A2(new_n583), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n792), .A2(KEYINPUT42), .A3(new_n775), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT109), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n729), .A2(new_n789), .A3(new_n730), .A4(new_n786), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n752), .A3(new_n711), .ZN(new_n796));
  INV_X1    g610(.A(new_n775), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n593), .A2(G472), .B1(new_n582), .B2(KEYINPUT32), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n791), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n799), .A3(new_n800), .A4(KEYINPUT42), .ZN(new_n801));
  INV_X1    g615(.A(new_n795), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n595), .A2(new_n802), .A3(new_n650), .A4(new_n753), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT42), .ZN(new_n804));
  AOI22_X1  g618(.A1(new_n794), .A2(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(KEYINPUT110), .B(G131), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G33));
  NAND3_X1  g621(.A1(new_n758), .A2(new_n713), .A3(new_n802), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  NOR3_X1   g623(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT45), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  OAI21_X1  g625(.A(G469), .B1(new_n284), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(KEYINPUT46), .B(new_n295), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT111), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n285), .A2(new_n811), .A3(new_n287), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n270), .A2(new_n283), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n194), .B1(new_n816), .B2(KEYINPUT45), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n294), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT46), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n814), .A2(new_n293), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT112), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n818), .A2(KEYINPUT46), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n814), .A2(new_n820), .A3(new_n824), .A4(new_n293), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n725), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n826), .A2(new_n192), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT43), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n829), .A2(new_n751), .A3(new_n457), .A4(new_n503), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n499), .A2(new_n502), .A3(G475), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n686), .A2(new_n687), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT113), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n457), .A2(new_n503), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n751), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n830), .B1(new_n836), .B2(KEYINPUT43), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n655), .A3(new_n703), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT44), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n382), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n676), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n838), .B2(new_n839), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n828), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n245), .ZN(G39));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n826), .A2(new_n846), .A3(new_n192), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n826), .B2(new_n192), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n595), .A2(new_n650), .A3(new_n676), .A4(new_n841), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n753), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  NAND4_X1  g666(.A1(new_n729), .A2(new_n760), .A3(new_n730), .A4(new_n786), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n382), .A2(KEYINPUT117), .A3(new_n760), .A4(new_n786), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n579), .A2(new_n583), .A3(new_n744), .ZN(new_n858));
  INV_X1    g672(.A(new_n505), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n649), .A2(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n675), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n504), .B(KEYINPUT119), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n859), .B(new_n830), .C1(KEYINPUT43), .C2(new_n836), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(new_n779), .ZN(new_n866));
  INV_X1    g680(.A(new_n766), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n862), .B(new_n863), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n864), .A2(new_n799), .A3(new_n857), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT48), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n869), .A2(KEYINPUT48), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n505), .A2(new_n837), .A3(new_n783), .A4(new_n857), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n732), .A2(new_n735), .A3(new_n676), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n864), .A2(KEYINPUT50), .A3(new_n780), .A4(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n837), .A2(new_n780), .A3(new_n505), .A4(new_n874), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT50), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n873), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n750), .ZN(new_n880));
  INV_X1    g694(.A(new_n751), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n857), .A2(new_n858), .A3(new_n880), .A4(new_n860), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n751), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n760), .A2(new_n191), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n847), .B2(new_n848), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n866), .A2(new_n676), .A3(new_n841), .ZN(new_n890));
  AOI211_X1 g704(.A(KEYINPUT51), .B(new_n887), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n889), .A2(new_n890), .ZN(new_n893));
  INV_X1    g707(.A(new_n887), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n872), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n382), .A2(new_n193), .A3(new_n496), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT114), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n734), .A2(new_n495), .A3(new_n676), .A4(new_n374), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT114), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n691), .A3(new_n904), .A4(new_n712), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n769), .A2(new_n902), .A3(new_n719), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n808), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n457), .A2(new_n503), .A3(new_n495), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n512), .B1(new_n752), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n657), .A2(new_n193), .A3(new_n841), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n796), .A2(new_n783), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n651), .A3(new_n704), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n899), .B1(new_n913), .B2(KEYINPUT116), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n722), .A2(new_n784), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AND4_X1   g731(.A1(new_n677), .A2(new_n746), .A3(new_n712), .A4(new_n789), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(new_n745), .A3(new_n192), .A4(new_n702), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(KEYINPUT52), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n722), .A2(KEYINPUT115), .A3(new_n784), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n917), .A2(new_n754), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n722), .A2(new_n919), .A3(new_n754), .A4(new_n784), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT52), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n767), .A2(new_n771), .A3(new_n763), .A4(new_n781), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n805), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT116), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n907), .B2(new_n912), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n914), .A2(new_n926), .A3(new_n928), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n913), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n923), .B(KEYINPUT52), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n899), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n927), .A2(new_n805), .A3(new_n907), .A4(new_n912), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n899), .A3(new_n926), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT53), .B1(new_n932), .B2(new_n933), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT54), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT120), .B(new_n872), .C1(new_n891), .C2(new_n895), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n898), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  OR2_X1    g758(.A1(G952), .A2(G953), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n760), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT49), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n858), .A2(new_n775), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n786), .B1(new_n947), .B2(KEYINPUT49), .ZN(new_n950));
  OR4_X1    g764(.A1(new_n736), .A2(new_n949), .A3(new_n836), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G75));
  NOR2_X1   g766(.A1(new_n261), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n188), .B1(new_n931), .B2(new_n934), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT56), .B1(new_n955), .B2(new_n373), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n336), .A2(new_n346), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(new_n344), .Z(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT55), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n956), .A2(new_n957), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n958), .B1(new_n963), .B2(new_n965), .ZN(G51));
  INV_X1    g780(.A(new_n912), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n906), .A2(new_n808), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT116), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n928), .A3(KEYINPUT53), .A4(new_n930), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n922), .A2(new_n925), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n923), .B(new_n924), .ZN(new_n973));
  AOI21_X1  g787(.A(KEYINPUT53), .B1(new_n937), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(KEYINPUT54), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(KEYINPUT122), .A3(new_n936), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n931), .A2(new_n934), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(new_n978), .A3(KEYINPUT54), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n294), .B(KEYINPUT57), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n292), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n955), .A2(new_n815), .A3(new_n817), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n953), .B1(new_n982), .B2(new_n983), .ZN(G54));
  AND2_X1   g798(.A1(KEYINPUT58), .A2(G475), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(KEYINPUT123), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n955), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n446), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n446), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n989), .A2(new_n990), .A3(new_n953), .ZN(G60));
  NAND2_X1  g805(.A1(G478), .A2(G902), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT59), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n941), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n667), .A2(new_n672), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n953), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n995), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n976), .A2(new_n997), .A3(new_n979), .A4(new_n993), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G63));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT60), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n977), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n626), .B2(new_n627), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n701), .B(KEYINPUT124), .Z(new_n1004));
  NAND3_X1  g818(.A1(new_n977), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n954), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1003), .A2(KEYINPUT61), .A3(new_n954), .A4(new_n1005), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G66));
  OAI21_X1  g824(.A(G953), .B1(new_n511), .B2(new_n342), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n910), .A2(new_n651), .A3(new_n704), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n927), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1011), .B1(new_n1013), .B2(G953), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n960), .B1(G898), .B2(new_n261), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1014), .B(new_n1015), .ZN(G69));
  XOR2_X1   g830(.A(new_n553), .B(new_n437), .Z(new_n1017));
  NAND2_X1  g831(.A1(G900), .A2(G953), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n799), .A2(new_n677), .A3(new_n746), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n808), .B1(new_n828), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n844), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n917), .A2(new_n754), .A3(new_n921), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n805), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n851), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1017), .B(new_n1018), .C1(new_n1024), .C2(G953), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n917), .A2(new_n748), .A3(new_n754), .A4(new_n921), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT62), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n752), .A2(new_n908), .ZN(new_n1029));
  AND3_X1   g843(.A1(new_n758), .A2(new_n738), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n844), .B1(new_n842), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1028), .A2(new_n1031), .A3(new_n851), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1032), .A2(new_n261), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1025), .B1(new_n1033), .B2(new_n1017), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(G72));
  INV_X1    g850(.A(KEYINPUT126), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1013), .ZN(new_n1038));
  OR2_X1    g852(.A1(new_n1024), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g853(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1037), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1037), .B(new_n1042), .C1(new_n1024), .C2(new_n1038), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(new_n547), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1043), .A2(new_n1045), .A3(new_n585), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n586), .A2(new_n559), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n938), .A2(new_n939), .A3(new_n1042), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT127), .ZN(new_n1049));
  XNOR2_X1  g863(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1042), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1051), .A2(new_n546), .A3(new_n585), .ZN(new_n1052));
  NAND3_X1  g866(.A1(new_n1050), .A2(new_n1052), .A3(new_n954), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1046), .A2(new_n1053), .ZN(G57));
endmodule


