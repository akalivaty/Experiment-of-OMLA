//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1192, new_n1193, new_n1194,
    new_n1196, new_n1197, new_n1198, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n207), .B1(new_n201), .B2(new_n203), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n206), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n203), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n214), .B(new_n227), .C1(new_n231), .C2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(G97), .B(G107), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G58), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  AOI21_X1  g0049(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G226), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n251), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n222), .A3(new_n253), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n250), .B1(new_n256), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g0067(.A(G1), .B(G13), .C1(new_n257), .C2(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n270), .A2(G238), .B1(G274), .B2(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT13), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n263), .A2(new_n274), .A3(new_n271), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT14), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(new_n277), .A3(G169), .ZN(new_n278));
  INV_X1    g0078(.A(new_n275), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n263), .B2(new_n271), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT14), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n278), .B(new_n283), .C1(new_n284), .C2(new_n276), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n286), .A2(new_n228), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(G1), .B2(new_n229), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n223), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n223), .A2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n229), .A2(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n291), .B1(new_n292), .B2(new_n206), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n287), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(KEYINPUT11), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(KEYINPUT11), .ZN(new_n300));
  INV_X1    g0100(.A(G1), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n301), .A2(G13), .A3(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n223), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT12), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n290), .A2(new_n299), .A3(new_n300), .A4(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n285), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n281), .B2(G190), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n276), .A2(KEYINPUT71), .A3(G200), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT71), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n281), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT18), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT8), .B(G58), .Z(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n303), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n316), .B2(new_n288), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n221), .A2(new_n223), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n202), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n293), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT7), .B1(new_n261), .B2(new_n229), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n223), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n252), .B2(G20), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT73), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n322), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n287), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n223), .B1(new_n327), .B2(new_n328), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n318), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n266), .A2(G274), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n269), .B2(new_n222), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n258), .A2(new_n260), .A3(G226), .A4(G1698), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n339), .B1(G33), .B2(G87), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n252), .A2(KEYINPUT75), .A3(G223), .A4(new_n253), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n252), .A2(KEYINPUT74), .A3(G226), .A4(G1698), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n258), .A2(new_n260), .A3(G223), .A4(new_n253), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT75), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n340), .A2(new_n341), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  AOI211_X1 g0146(.A(new_n284), .B(new_n337), .C1(new_n346), .C2(new_n250), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n341), .A3(new_n342), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n338), .A2(new_n339), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G87), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n250), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n337), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n282), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n315), .B1(new_n335), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n322), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT73), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n327), .B2(KEYINPUT73), .ZN(new_n359));
  OAI211_X1 g0159(.A(KEYINPUT16), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(new_n297), .A3(new_n334), .ZN(new_n361));
  INV_X1    g0161(.A(new_n318), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n352), .A2(G179), .A3(new_n353), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n337), .B1(new_n346), .B2(new_n250), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n282), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(KEYINPUT18), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n352), .A2(new_n353), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G200), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n352), .A2(G190), .A3(new_n353), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n369), .A2(new_n361), .A3(new_n362), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT76), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n375), .B(new_n337), .C1(new_n346), .C2(new_n250), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n311), .B1(new_n352), .B2(new_n353), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n335), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n356), .A2(new_n367), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  MUX2_X1   g0182(.A(G222), .B(G223), .S(G1698), .Z(new_n383));
  OAI21_X1  g0183(.A(new_n250), .B1(new_n383), .B2(new_n261), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n206), .B2(new_n261), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n336), .B1(new_n269), .B2(new_n255), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n284), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(G169), .B2(new_n387), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n229), .B1(new_n205), .B2(new_n208), .ZN(new_n390));
  INV_X1    g0190(.A(new_n316), .ZN(new_n391));
  INV_X1    g0191(.A(G150), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n391), .A2(new_n292), .B1(new_n392), .B2(new_n294), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n297), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  MUX2_X1   g0194(.A(new_n302), .B(new_n288), .S(G50), .Z(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n387), .A2(new_n311), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n399), .B1(G190), .B2(new_n387), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT70), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n397), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(KEYINPUT70), .A2(KEYINPUT9), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n401), .A2(new_n402), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n396), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n400), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT10), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT10), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n409), .B(new_n400), .C1(new_n403), .C2(new_n406), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n398), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n314), .A2(new_n382), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT69), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n316), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(new_n292), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n287), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n303), .A2(new_n206), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n288), .B2(new_n206), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n336), .B1(new_n269), .B2(new_n216), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n252), .A2(G238), .A3(G1698), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n423));
  INV_X1    g0223(.A(G107), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n422), .B(new_n423), .C1(new_n424), .C2(new_n252), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(KEYINPUT67), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n268), .B1(new_n425), .B2(KEYINPUT67), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n420), .B1(new_n429), .B2(new_n282), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT68), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n429), .B2(G179), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(KEYINPUT68), .A3(new_n284), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n420), .B1(new_n429), .B2(new_n375), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n428), .A2(new_n311), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n413), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n433), .A2(new_n434), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n430), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(KEYINPUT69), .C1(new_n437), .C2(new_n436), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n412), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n254), .B2(new_n216), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n445), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n250), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n301), .B(G45), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n268), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G257), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n451), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n264), .A2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT79), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(G274), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n450), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G169), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n462), .B1(new_n449), .B2(new_n250), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G179), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT6), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n244), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n424), .A2(G97), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(G20), .B1(G77), .B2(new_n293), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n424), .B1(new_n327), .B2(new_n328), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(KEYINPUT77), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(KEYINPUT77), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n297), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n302), .A2(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n301), .A2(G33), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n302), .A2(new_n479), .A3(new_n228), .A4(new_n286), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n478), .B1(new_n481), .B2(G97), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n465), .A2(new_n467), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT78), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n470), .A2(new_n468), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n468), .B2(new_n244), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n486), .A2(new_n229), .B1(new_n206), .B2(new_n294), .ZN(new_n487));
  INV_X1    g0287(.A(new_n473), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n287), .B1(new_n490), .B2(new_n475), .ZN(new_n491));
  INV_X1    g0291(.A(new_n482), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n482), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n466), .A2(new_n311), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(G190), .B2(new_n466), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n483), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n259), .A2(G33), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n501));
  OAI21_X1  g0301(.A(G303), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n258), .A2(new_n260), .A3(G257), .A4(new_n253), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n258), .A2(new_n260), .A3(G264), .A4(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n505), .A2(new_n250), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n268), .B(G270), .C1(new_n451), .C2(new_n452), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n461), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(G169), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n302), .A2(new_n479), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT80), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(G116), .A4(new_n287), .ZN(new_n512));
  INV_X1    g0312(.A(G116), .ZN(new_n513));
  OAI21_X1  g0313(.A(KEYINPUT80), .B1(new_n480), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n303), .A2(new_n513), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n286), .A2(new_n228), .B1(G20), .B2(new_n513), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n448), .B(new_n229), .C1(G33), .C2(new_n217), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(KEYINPUT20), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT20), .B1(new_n517), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n499), .B1(new_n509), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n512), .A2(new_n514), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n524), .B(new_n516), .C1(new_n520), .C2(new_n519), .ZN(new_n525));
  INV_X1    g0325(.A(new_n508), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n505), .A2(new_n250), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT21), .A4(G169), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n506), .A2(new_n508), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n525), .A2(new_n530), .A3(G179), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n424), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n302), .B2(G107), .ZN(new_n535));
  AOI22_X1  g0335(.A1(G107), .A2(new_n481), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT82), .ZN(new_n537));
  INV_X1    g0337(.A(G87), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n539), .A2(new_n258), .A3(new_n260), .A4(new_n229), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n252), .A2(KEYINPUT22), .A3(new_n229), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n229), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n424), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT24), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n542), .A2(new_n543), .A3(new_n549), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n537), .B1(new_n554), .B2(new_n297), .ZN(new_n555));
  AOI211_X1 g0355(.A(KEYINPUT82), .B(new_n287), .C1(new_n551), .C2(new_n553), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n536), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n258), .A2(new_n260), .A3(G257), .A4(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n258), .A2(new_n260), .A3(G250), .A4(new_n253), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(G264), .A2(new_n454), .B1(new_n561), .B2(new_n250), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n461), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(G179), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n282), .B2(new_n563), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n532), .B1(new_n557), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n252), .A2(G238), .A3(new_n253), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n252), .A2(G244), .A3(G1698), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n544), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n250), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n301), .A2(G45), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G250), .ZN(new_n572));
  INV_X1    g0372(.A(G274), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n250), .A2(new_n572), .B1(new_n573), .B2(new_n571), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G200), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT19), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n229), .B1(new_n251), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n538), .A2(new_n217), .A3(new_n424), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n258), .A2(new_n260), .A3(new_n229), .A4(G68), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n578), .B1(new_n292), .B2(new_n217), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n297), .B1(new_n415), .B2(new_n303), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n481), .A2(G87), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n574), .B1(new_n569), .B2(new_n250), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G190), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n577), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n284), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n585), .B1(new_n415), .B2(new_n480), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(G169), .C2(new_n587), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n311), .B1(new_n562), .B2(new_n461), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n561), .A2(new_n250), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n268), .B(G264), .C1(new_n451), .C2(new_n452), .ZN(new_n596));
  AND4_X1   g0396(.A1(G190), .A2(new_n595), .A3(new_n461), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n598), .B(new_n536), .C1(new_n555), .C2(new_n556), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n525), .B1(G190), .B2(new_n530), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n311), .B2(new_n530), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n593), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n443), .A2(new_n498), .A3(new_n566), .A4(new_n602), .ZN(G372));
  INV_X1    g0403(.A(new_n592), .ZN(new_n604));
  AOI211_X1 g0404(.A(new_n375), .B(new_n574), .C1(new_n569), .C2(new_n250), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(G200), .B2(new_n576), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n585), .A2(KEYINPUT83), .A3(new_n586), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT83), .B1(new_n585), .B2(new_n586), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(G169), .B1(new_n570), .B2(new_n575), .ZN(new_n610));
  AOI211_X1 g0410(.A(G179), .B(new_n574), .C1(new_n569), .C2(new_n250), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n606), .A2(new_n609), .B1(new_n612), .B2(new_n591), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n599), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n566), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n604), .B1(new_n615), .B2(new_n498), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n483), .B2(new_n593), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n465), .A2(new_n467), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n613), .A2(new_n493), .A3(new_n619), .A4(new_n494), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n443), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n363), .A2(new_n625), .A3(new_n366), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n363), .B2(new_n366), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n315), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT84), .B1(new_n335), .B2(new_n355), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n363), .A2(new_n625), .A3(new_n366), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n435), .B1(new_n285), .B2(new_n306), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n374), .A2(new_n381), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n313), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n408), .A2(new_n410), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n398), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n624), .A2(new_n638), .ZN(G369));
  INV_X1    g0439(.A(G13), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(G20), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n301), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT27), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G213), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(G343), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n557), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n648), .A2(new_n599), .B1(new_n557), .B2(new_n565), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n557), .A2(new_n565), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n647), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n532), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n601), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n525), .A2(new_n647), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  MUX2_X1   g0457(.A(new_n655), .B(new_n654), .S(new_n657), .Z(new_n658));
  INV_X1    g0458(.A(G330), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT86), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(KEYINPUT86), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n653), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n654), .A2(new_n647), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n651), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n663), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n212), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n580), .A2(G116), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n232), .B2(new_n671), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT29), .ZN(new_n676));
  INV_X1    g0476(.A(new_n647), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n623), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n498), .A2(new_n602), .A3(new_n566), .A4(new_n677), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT87), .B1(new_n528), .B2(new_n284), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n526), .A2(new_n681), .A3(G179), .A4(new_n527), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n587), .A2(new_n562), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n680), .A2(new_n466), .A3(new_n682), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND4_X1   g0486(.A1(new_n450), .A2(new_n463), .A3(new_n562), .A4(new_n587), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(KEYINPUT30), .A3(new_n682), .A4(new_n680), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n530), .A2(G179), .A3(new_n587), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n464), .A3(new_n563), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n686), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n647), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT31), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n647), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n679), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n477), .A2(new_n482), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n619), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n589), .A2(new_n592), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT26), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n701), .B1(KEYINPUT26), .B2(new_n620), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n647), .B1(new_n616), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n678), .B(new_n697), .C1(new_n676), .C2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n675), .B1(new_n705), .B2(G1), .ZN(G364));
  NAND2_X1  g0506(.A1(new_n661), .A2(new_n662), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n658), .A2(new_n659), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT88), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n301), .B1(new_n641), .B2(G45), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n670), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n707), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT89), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n229), .A2(G190), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n311), .A2(G179), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(G283), .A2(new_n719), .B1(new_n722), .B2(G329), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  INV_X1    g0524(.A(G303), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n229), .A2(new_n375), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n717), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n284), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G322), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n725), .A2(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n716), .A2(new_n728), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(new_n252), .B(new_n731), .C1(G311), .C2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n229), .B1(new_n720), .B2(G190), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n724), .B(new_n734), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT92), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n375), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G326), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n739), .A2(G190), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(KEYINPUT33), .B(G317), .Z(new_n744));
  OAI21_X1  g0544(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n729), .A2(new_n221), .B1(new_n732), .B2(new_n206), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT91), .ZN(new_n747));
  INV_X1    g0547(.A(new_n740), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n747), .B1(new_n295), .B2(new_n748), .C1(new_n223), .C2(new_n743), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n718), .A2(new_n424), .ZN(new_n750));
  INV_X1    g0550(.A(new_n727), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n261), .B(new_n750), .C1(G87), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n736), .A2(new_n217), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G159), .ZN(new_n755));
  OAI21_X1  g0555(.A(KEYINPUT32), .B1(new_n721), .B2(new_n755), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n721), .A2(KEYINPUT32), .A3(new_n755), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n752), .A2(new_n754), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n737), .A2(new_n745), .B1(new_n749), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n228), .B1(G20), .B2(new_n282), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n760), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n252), .A2(new_n212), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(KEYINPUT90), .B2(G355), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(KEYINPUT90), .B2(G355), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(G116), .B2(new_n212), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n248), .A2(G45), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n669), .A2(new_n252), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(new_n265), .B2(new_n233), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n761), .B(new_n712), .C1(new_n766), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(new_n658), .B2(new_n764), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n714), .A2(new_n715), .A3(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n435), .A2(new_n677), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n677), .A2(new_n420), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n441), .B1(new_n438), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT97), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n647), .B1(new_n616), .B2(new_n622), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT98), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n783), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n784), .A2(KEYINPUT98), .A3(new_n785), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n712), .B1(new_n791), .B2(new_n697), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(new_n697), .B2(new_n791), .ZN(new_n793));
  INV_X1    g0593(.A(new_n729), .ZN(new_n794));
  XNOR2_X1  g0594(.A(KEYINPUT95), .B(G143), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n794), .A2(new_n795), .B1(new_n733), .B2(G159), .ZN(new_n796));
  INV_X1    g0596(.A(G137), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n796), .B1(new_n748), .B2(new_n797), .C1(new_n392), .C2(new_n743), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT34), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n252), .B1(new_n727), .B2(new_n295), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n718), .A2(new_n223), .B1(new_n721), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n736), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n804), .C1(G58), .C2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n800), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n727), .A2(new_n424), .B1(new_n732), .B2(new_n513), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n729), .A2(new_n735), .B1(new_n721), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n261), .B1(new_n718), .B2(new_n538), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n808), .A2(new_n810), .A3(new_n811), .A4(new_n753), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n812), .B1(new_n813), .B2(new_n743), .C1(new_n725), .C2(new_n748), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT96), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(KEYINPUT96), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n816), .A2(new_n760), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n712), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n760), .A2(new_n762), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n206), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n821), .C1(new_n787), .C2(new_n763), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n793), .A2(new_n822), .ZN(G384));
  NOR3_X1   g0623(.A1(new_n232), .A2(new_n206), .A3(new_n319), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n201), .A2(new_n223), .ZN(new_n825));
  OAI211_X1 g0625(.A(G1), .B(new_n640), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(G116), .B(new_n231), .C1(new_n471), .C2(KEYINPUT35), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(KEYINPUT35), .B2(new_n471), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(KEYINPUT36), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(KEYINPUT36), .B2(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n306), .A2(new_n647), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n307), .A2(new_n313), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n285), .A2(new_n306), .A3(new_n647), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n783), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT102), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n679), .A2(new_n694), .A3(new_n838), .A4(new_n695), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n364), .B(new_n645), .C1(new_n282), .C2(new_n365), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n363), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n371), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n360), .A2(new_n297), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n362), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n842), .A2(new_n848), .B1(new_n335), .B2(new_n378), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n845), .B1(new_n849), .B2(new_n844), .ZN(new_n850));
  INV_X1    g0650(.A(new_n645), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(KEYINPUT38), .C1(new_n382), .C2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n356), .A2(new_n367), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n634), .ZN(new_n857));
  INV_X1    g0657(.A(new_n852), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n859), .A2(KEYINPUT99), .A3(KEYINPUT38), .A4(new_n850), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n363), .A2(new_n851), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n632), .B2(new_n634), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n371), .B(new_n863), .C1(new_n626), .C2(new_n627), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT37), .B1(new_n335), .B2(new_n378), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n865), .A2(KEYINPUT37), .B1(new_n843), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n862), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT40), .B1(new_n841), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT40), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n859), .B2(new_n850), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n852), .B1(new_n856), .B2(new_n634), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n848), .A2(new_n842), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n371), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(KEYINPUT37), .B1(new_n866), .B2(new_n843), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n874), .A2(new_n877), .A3(new_n862), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n836), .A2(new_n840), .A3(new_n872), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n871), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(G330), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n659), .B1(new_n837), .B2(new_n839), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n443), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT103), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n881), .A2(new_n443), .A3(new_n840), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n780), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n785), .B2(new_n787), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n879), .A3(new_n834), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n632), .B2(new_n851), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT39), .B1(new_n873), .B2(new_n878), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT39), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n861), .A2(new_n868), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n861), .A2(new_n868), .A3(new_n895), .A4(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n285), .A2(new_n306), .A3(new_n677), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n893), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n678), .B1(new_n676), .B2(new_n703), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT101), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n905), .A2(new_n443), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n906), .B1(new_n905), .B2(new_n443), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n638), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n904), .B(new_n911), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n888), .A2(new_n912), .B1(new_n301), .B2(new_n641), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n913), .A2(KEYINPUT104), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n888), .A2(new_n912), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n913), .B2(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n830), .B1(new_n914), .B2(new_n916), .ZN(G367));
  NAND3_X1  g0717(.A1(new_n493), .A2(new_n494), .A3(new_n647), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n493), .A2(new_n494), .A3(new_n619), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n498), .A2(new_n918), .B1(new_n920), .B2(new_n647), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n665), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n699), .B1(new_n921), .B2(new_n650), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n677), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n609), .A2(new_n677), .ZN(new_n929));
  MUX2_X1   g0729(.A(new_n613), .B(new_n604), .S(new_n929), .Z(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT43), .B1(new_n930), .B2(KEYINPUT105), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT105), .B2(new_n930), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT106), .Z(new_n935));
  XNOR2_X1  g0735(.A(new_n932), .B(new_n935), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n653), .B(new_n921), .C1(new_n661), .C2(new_n662), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n670), .B(KEYINPUT41), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n667), .A2(new_n921), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n663), .A2(KEYINPUT107), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT44), .B1(new_n667), .B2(new_n921), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n667), .A2(KEYINPUT44), .A3(new_n921), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n663), .A2(KEYINPUT107), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n707), .A2(new_n652), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n951), .A2(new_n663), .ZN(new_n952));
  INV_X1    g0752(.A(new_n664), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n950), .A2(new_n705), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n940), .B1(new_n955), .B2(new_n705), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n938), .B1(new_n956), .B2(new_n711), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n241), .A2(new_n773), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n765), .B1(new_n212), .B2(new_n415), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(new_n819), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n727), .A2(new_n221), .B1(new_n718), .B2(new_n206), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n252), .B1(new_n736), .B2(new_n223), .C1(new_n797), .C2(new_n721), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(G150), .C2(new_n794), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n742), .A2(G159), .B1(new_n201), .B2(new_n733), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n740), .A2(new_n795), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n964), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n751), .A2(G116), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n729), .A2(new_n725), .B1(new_n718), .B2(new_n217), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(G317), .B2(new_n722), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n261), .B1(new_n732), .B2(new_n813), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G107), .B2(new_n805), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n971), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n735), .A2(new_n743), .B1(new_n748), .B2(new_n809), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT47), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n760), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n978), .A2(new_n979), .ZN(new_n982));
  INV_X1    g0782(.A(new_n764), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n961), .B1(new_n981), .B2(new_n982), .C1(new_n930), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n957), .A2(new_n984), .ZN(G387));
  OR3_X1    g0785(.A1(new_n391), .A2(KEYINPUT50), .A3(G50), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n672), .B(new_n265), .C1(new_n223), .C2(new_n206), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT109), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT50), .B1(new_n391), .B2(G50), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n987), .A2(new_n988), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n772), .B1(new_n991), .B2(new_n992), .C1(new_n238), .C2(new_n265), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(G107), .B2(new_n212), .C1(new_n672), .C2(new_n767), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n819), .B1(new_n994), .B2(new_n765), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n652), .B2(new_n983), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n729), .A2(new_n295), .B1(new_n732), .B2(new_n223), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n727), .A2(new_n206), .B1(new_n721), .B2(new_n392), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n252), .B1(new_n718), .B2(new_n217), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n736), .A2(new_n415), .ZN(new_n1000));
  NOR4_X1   g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n1001), .B1(new_n755), .B2(new_n748), .C1(new_n391), .C2(new_n743), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G317), .A2(new_n794), .B1(new_n733), .B2(G303), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n748), .B2(new_n730), .C1(new_n809), .C2(new_n743), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n813), .B2(new_n736), .C1(new_n735), .C2(new_n727), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT110), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT49), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n261), .B1(new_n718), .B2(new_n513), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G326), .B2(new_n722), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT49), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1002), .B1(new_n1009), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n996), .B1(new_n1014), .B2(new_n760), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(new_n954), .B2(new_n711), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n954), .A2(new_n705), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n670), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n954), .A2(new_n705), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1016), .B1(new_n1018), .B2(new_n1019), .ZN(G393));
  NAND3_X1  g0820(.A1(new_n1017), .A2(new_n948), .A3(new_n949), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1021), .A2(new_n955), .A3(new_n670), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n740), .A2(G317), .B1(G311), .B2(new_n794), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT52), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n727), .A2(new_n813), .B1(new_n721), .B2(new_n730), .ZN(new_n1025));
  OR4_X1    g0825(.A1(new_n252), .A2(new_n1024), .A3(new_n750), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G294), .A2(new_n733), .B1(new_n805), .B2(G116), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n743), .B2(new_n725), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT112), .Z(new_n1029));
  OAI22_X1  g0829(.A1(new_n748), .A2(new_n392), .B1(new_n755), .B2(new_n729), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT51), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G68), .A2(new_n751), .B1(new_n722), .B2(new_n795), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT111), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n742), .A2(new_n201), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n736), .A2(new_n206), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n252), .B1(new_n718), .B2(new_n538), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n316), .C2(new_n733), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1026), .A2(new_n1029), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n760), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n245), .A2(new_n773), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n765), .B1(new_n217), .B2(new_n212), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n712), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n921), .B2(new_n764), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n950), .B2(new_n711), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1022), .A2(new_n1047), .ZN(G390));
  INV_X1    g0848(.A(new_n820), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n712), .B1(new_n1049), .B2(new_n316), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n729), .A2(new_n513), .B1(new_n718), .B2(new_n223), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n732), .A2(new_n217), .B1(new_n721), .B2(new_n735), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n261), .B1(new_n727), .B2(new_n538), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1037), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(new_n424), .B2(new_n743), .C1(new_n813), .C2(new_n748), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n727), .A2(new_n392), .ZN(new_n1056));
  XOR2_X1   g0856(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G159), .B2(new_n805), .ZN(new_n1059));
  XOR2_X1   g0859(.A(KEYINPUT54), .B(G143), .Z(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT116), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n733), .ZN(new_n1062));
  INV_X1    g0862(.A(G125), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n729), .A2(new_n803), .B1(new_n721), .B2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n261), .B(new_n1064), .C1(new_n201), .C2(new_n719), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1059), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(G128), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1067), .A2(new_n748), .B1(new_n743), .B2(new_n797), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1055), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1050), .B1(new_n1069), .B2(new_n760), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n901), .B2(new_n763), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n902), .B1(new_n890), .B2(new_n835), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n899), .A2(new_n1072), .A3(new_n900), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n703), .A2(new_n782), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n780), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n834), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n902), .A3(new_n869), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n787), .A2(new_n696), .A3(G330), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n835), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1073), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n836), .A2(new_n840), .A3(G330), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1083));
  OAI21_X1  g0883(.A(KEYINPUT113), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n1082), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1088), .B2(new_n710), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n638), .B(new_n884), .C1(new_n907), .C2(new_n908), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n784), .B1(new_n883), .B2(KEYINPUT114), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1092), .B(new_n659), .C1(new_n837), .C2(new_n839), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n835), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1079), .A2(new_n1075), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1078), .A2(new_n835), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1082), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n891), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1090), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1084), .A2(new_n1087), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1084), .A2(new_n1100), .A3(new_n1087), .A4(KEYINPUT115), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1100), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n671), .B1(new_n1088), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(G378));
  INV_X1    g0909(.A(KEYINPUT57), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1090), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n411), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n396), .A3(new_n851), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n411), .B1(new_n397), .B2(new_n645), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n881), .B2(G330), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n881), .A2(G330), .A3(new_n1119), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n904), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n904), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n659), .B(new_n1118), .C1(new_n871), .C2(new_n880), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1123), .A2(new_n1126), .A3(KEYINPUT119), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT119), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1121), .A2(new_n904), .A3(new_n1128), .A4(new_n1122), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1110), .B1(new_n1111), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT120), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(KEYINPUT120), .B(new_n1110), .C1(new_n1111), .C2(new_n1130), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1111), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1110), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n671), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1133), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1127), .A2(new_n711), .A3(new_n1129), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n712), .B1(new_n1049), .B2(new_n201), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n252), .A2(G41), .ZN(new_n1141));
  AOI211_X1 g0941(.A(G50), .B(new_n1141), .C1(new_n257), .C2(new_n264), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT118), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1141), .B1(new_n223), .B2(new_n736), .C1(new_n206), .C2(new_n727), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n729), .A2(new_n424), .B1(new_n721), .B2(new_n813), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n718), .A2(new_n221), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n732), .A2(new_n415), .ZN(new_n1147));
  NOR4_X1   g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n217), .B2(new_n743), .C1(new_n513), .C2(new_n748), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT58), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G128), .A2(new_n794), .B1(new_n733), .B2(G137), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n392), .B2(new_n736), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n751), .B2(new_n1061), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n1063), .B2(new_n748), .C1(new_n803), .C2(new_n743), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n719), .A2(G159), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G33), .B(G41), .C1(new_n722), .C2(G124), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(KEYINPUT59), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1151), .B1(new_n1150), .B2(new_n1149), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1140), .B1(new_n1161), .B2(new_n760), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1119), .B2(new_n763), .ZN(new_n1163));
  AND2_X1   g0963(.A1(new_n1139), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1138), .A2(new_n1164), .ZN(G375));
  INV_X1    g0965(.A(KEYINPUT121), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n710), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(KEYINPUT121), .A3(new_n711), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n819), .B1(new_n223), .B2(new_n820), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n727), .A2(new_n217), .B1(new_n732), .B2(new_n424), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n729), .A2(new_n813), .B1(new_n721), .B2(new_n725), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n261), .B1(new_n718), .B2(new_n206), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1000), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n513), .B2(new_n743), .C1(new_n735), .C2(new_n748), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n748), .A2(new_n803), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n261), .B(new_n1146), .C1(G50), .C2(new_n805), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1061), .A2(new_n742), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G137), .A2(new_n794), .B1(new_n722), .B2(G128), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G159), .A2(new_n751), .B1(new_n733), .B2(G150), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1176), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(KEYINPUT122), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(KEYINPUT122), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n760), .ZN(new_n1186));
  OAI221_X1 g0986(.A(new_n1171), .B1(new_n1184), .B2(new_n1186), .C1(new_n834), .C2(new_n763), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1169), .A2(new_n1170), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1168), .A2(new_n1090), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1189), .A2(new_n939), .A3(new_n1106), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(G381));
  OR2_X1    g0991(.A1(G393), .A2(G396), .ZN(new_n1192));
  OR4_X1    g0992(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1138), .A2(new_n1108), .A3(new_n1164), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1193), .A2(new_n1194), .A3(G381), .ZN(G407));
  NAND2_X1  g0995(.A1(new_n646), .A2(G213), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT123), .Z(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G407), .B(G213), .C1(new_n1194), .C2(new_n1198), .ZN(G409));
  INV_X1    g0999(.A(KEYINPUT60), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1189), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1201), .A2(new_n670), .A3(new_n1106), .A4(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1203), .A2(new_n1188), .A3(G384), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G384), .B1(new_n1203), .B2(new_n1188), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1138), .A2(G378), .A3(new_n1164), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1111), .A2(new_n1130), .A3(new_n940), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1163), .B1(new_n1209), .B2(new_n710), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1108), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT124), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT124), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n1108), .C1(new_n1208), .C2(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1198), .B(new_n1206), .C1(new_n1207), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT62), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1198), .B1(new_n1207), .B2(new_n1215), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1197), .A2(G2897), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1206), .B(new_n1219), .Z(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1138), .A2(G378), .A3(new_n1164), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(new_n1198), .A4(new_n1206), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1217), .A2(new_n1221), .A3(new_n1222), .A4(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G387), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n957), .A2(new_n984), .A3(G390), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(G393), .A2(G396), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1192), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1229), .A2(new_n1192), .A3(new_n1232), .A4(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  XOR2_X1   g1036(.A(new_n1236), .B(KEYINPUT125), .Z(new_n1237));
  NAND2_X1  g1037(.A1(new_n1227), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1216), .A2(new_n1240), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1224), .A2(KEYINPUT63), .A3(new_n1198), .A4(new_n1206), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1236), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1239), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1238), .A2(new_n1244), .ZN(G405));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1206), .A2(new_n1246), .A3(KEYINPUT127), .ZN(new_n1247));
  OAI21_X1  g1047(.A(KEYINPUT127), .B1(new_n1206), .B2(new_n1246), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(new_n1236), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G375), .A2(new_n1108), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1206), .A2(new_n1246), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1223), .A3(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1250), .B(new_n1253), .ZN(G402));
endmodule


