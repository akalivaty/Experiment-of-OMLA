//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .A3(G107), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT78), .A2(G104), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT78), .A2(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT79), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(new_n193), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n197), .B1(new_n198), .B2(G107), .ZN(new_n199));
  NOR4_X1   g013(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT79), .A4(new_n191), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n195), .B(new_n196), .C1(new_n199), .C2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT4), .ZN(new_n202));
  OR2_X1    g016(.A1(KEYINPUT78), .A2(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(KEYINPUT78), .A2(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(G107), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(KEYINPUT79), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n196), .B1(new_n206), .B2(new_n195), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n195), .B1(new_n199), .B2(new_n200), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G101), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n212), .A3(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n218), .ZN(new_n222));
  OR2_X1    g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n219), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n211), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n188), .B1(new_n208), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n209), .A2(G101), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(KEYINPUT4), .A3(new_n201), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT80), .A3(new_n226), .A4(new_n211), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n194), .B1(G104), .B2(new_n191), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n201), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n201), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n217), .A2(G146), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(G128), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n222), .ZN(new_n242));
  INV_X1    g056(.A(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n214), .A2(new_n216), .A3(new_n218), .A4(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT10), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n241), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n245), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n201), .A2(new_n235), .A3(new_n251), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n238), .A2(new_n248), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G131), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n259), .A3(new_n262), .A4(new_n257), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n232), .A2(new_n253), .A3(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G110), .B(G140), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G227), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n267), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n265), .B1(new_n232), .B2(new_n253), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n275));
  INV_X1    g089(.A(new_n252), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n246), .B1(new_n236), .B2(new_n237), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(KEYINPUT82), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT82), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n246), .C1(new_n236), .C2(new_n237), .ZN(new_n280));
  AOI211_X1 g094(.A(new_n275), .B(new_n265), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(KEYINPUT82), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n280), .A3(new_n252), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n283), .B2(new_n264), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n266), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n274), .B1(new_n285), .B2(new_n270), .ZN(new_n286));
  OAI21_X1  g100(.A(G469), .B1(new_n286), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT83), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT83), .B(G469), .C1(new_n286), .C2(G902), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n283), .A2(new_n264), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n275), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(KEYINPUT12), .A3(new_n264), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n272), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n232), .A2(new_n253), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n264), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n271), .B1(new_n298), .B2(new_n266), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n291), .B(new_n292), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n289), .A2(new_n290), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G221), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT77), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n304), .B2(new_n292), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n246), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n225), .A2(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n268), .A2(G224), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT85), .Z(new_n316));
  NAND2_X1  g130(.A1(new_n201), .A2(new_n235), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT81), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G116), .ZN(new_n320));
  OAI21_X1  g134(.A(G113), .B1(new_n320), .B2(KEYINPUT5), .ZN(new_n321));
  INV_X1    g135(.A(G116), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT68), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G116), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n325), .A3(G119), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(new_n320), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n327), .B2(KEYINPUT5), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT2), .B(G113), .Z(new_n329));
  AND3_X1   g143(.A1(new_n329), .A2(new_n326), .A3(new_n320), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n201), .A2(new_n233), .A3(new_n235), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n318), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n329), .B1(new_n326), .B2(new_n320), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n230), .A2(new_n336), .A3(new_n211), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n337), .A3(KEYINPUT84), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G122), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n333), .A2(new_n337), .A3(new_n342), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT6), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n342), .B1(new_n338), .B2(new_n339), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(KEYINPUT6), .A3(new_n341), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n316), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n313), .B1(G224), .B2(new_n268), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n311), .A2(KEYINPUT87), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n242), .A2(new_n245), .ZN(new_n353));
  OR3_X1    g167(.A1(new_n353), .A2(KEYINPUT87), .A3(G125), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n312), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT7), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n356), .A2(KEYINPUT88), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(KEYINPUT88), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n314), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n351), .A2(KEYINPUT7), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n360), .A2(new_n345), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n317), .B1(new_n330), .B2(new_n328), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n333), .A2(KEYINPUT86), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n342), .B(KEYINPUT8), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(KEYINPUT86), .C2(new_n333), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n309), .B1(new_n350), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n315), .B(KEYINPUT85), .ZN(new_n369));
  INV_X1    g183(.A(new_n349), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n348), .A2(new_n341), .B1(KEYINPUT6), .B2(new_n345), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n308), .A3(new_n366), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT89), .B(new_n309), .C1(new_n350), .C2(new_n367), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n304), .A2(G217), .A3(new_n268), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT94), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n243), .A2(G143), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n243), .A2(G143), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n383), .A2(G134), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n323), .A2(new_n325), .A3(G122), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n322), .A2(G122), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n191), .A3(new_n387), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n243), .B2(G143), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n217), .A2(KEYINPUT13), .A3(G128), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n382), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G134), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT93), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(KEYINPUT93), .A3(G134), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT95), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n386), .A2(new_n403), .A3(new_n387), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n323), .A2(new_n325), .A3(KEYINPUT14), .A4(G122), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G107), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n402), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n386), .A2(new_n403), .A3(new_n387), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n408), .A2(KEYINPUT95), .A3(G107), .A4(new_n405), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n388), .A2(G107), .ZN(new_n411));
  OR3_X1    g225(.A1(new_n383), .A2(G134), .A3(new_n384), .ZN(new_n412));
  OAI21_X1  g226(.A(G134), .B1(new_n383), .B2(new_n384), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n381), .A2(new_n401), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n391), .A2(new_n400), .A3(KEYINPUT94), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n380), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n401), .A2(new_n381), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n414), .ZN(new_n419));
  AND4_X1   g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .A4(new_n380), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n292), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT96), .ZN(new_n422));
  INV_X1    g236(.A(G478), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT15), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n419), .A3(new_n416), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n379), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n415), .A2(new_n416), .A3(new_n380), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n292), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n422), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n421), .A2(new_n424), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT97), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n431), .B2(new_n433), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n268), .ZN(new_n439));
  XOR2_X1   g253(.A(new_n439), .B(KEYINPUT98), .Z(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(G898), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n445));
  INV_X1    g259(.A(G237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n268), .A3(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n217), .ZN(new_n448));
  NOR2_X1   g262(.A1(G237), .A2(G953), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G143), .A3(G214), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT17), .A3(G131), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT16), .ZN(new_n453));
  INV_X1    g267(.A(G140), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n310), .A2(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n455), .B1(new_n458), .B2(new_n453), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n212), .ZN(new_n460));
  OAI211_X1 g274(.A(G146), .B(new_n455), .C1(new_n458), .C2(new_n453), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n452), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n451), .A2(G131), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT17), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n448), .A2(new_n262), .A3(new_n450), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n458), .A2(KEYINPUT90), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(KEYINPUT90), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G146), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n458), .A2(G146), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT18), .A2(G131), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n451), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n189), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n467), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(KEYINPUT91), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT91), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n462), .A2(new_n466), .B1(new_n473), .B2(new_n475), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n482), .A2(new_n478), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n445), .B(new_n292), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(KEYINPUT91), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n481), .A3(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT92), .B1(new_n489), .B2(G902), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n490), .A3(G475), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n468), .A2(KEYINPUT19), .A3(new_n469), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n492), .B1(KEYINPUT19), .B2(new_n458), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G146), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n461), .B(KEYINPUT75), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n463), .A2(new_n465), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n476), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n478), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n480), .B2(new_n483), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  INV_X1    g316(.A(G475), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .A4(new_n292), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n487), .A2(new_n488), .B1(new_n498), .B2(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n292), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT20), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n491), .A2(new_n508), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n437), .A2(new_n444), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n377), .A2(new_n378), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n187), .B1(new_n307), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G217), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(G234), .B2(new_n292), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n319), .A2(G128), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n243), .A2(KEYINPUT23), .A3(G119), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n319), .A2(G128), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(KEYINPUT23), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(G110), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n243), .A2(G119), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT24), .B(G110), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n471), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n495), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n460), .A2(new_n461), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n518), .A2(G110), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n527), .C1(new_n521), .C2(new_n522), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT22), .B(G137), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n268), .A2(G221), .A3(G234), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n528), .A3(new_n532), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT25), .B1(new_n536), .B2(new_n292), .ZN(new_n537));
  AND4_X1   g351(.A1(KEYINPUT25), .A2(new_n534), .A3(new_n292), .A4(new_n535), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n514), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n514), .A2(G902), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n536), .B(KEYINPUT76), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n258), .A2(G134), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n255), .A2(G137), .ZN(new_n547));
  OAI21_X1  g361(.A(G131), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n263), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT66), .B1(new_n246), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT65), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n225), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT65), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n264), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n263), .A2(new_n548), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT66), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n353), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n550), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT67), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(KEYINPUT70), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT70), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n549), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n353), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n226), .A2(new_n264), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT69), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT69), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n226), .B2(new_n264), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(KEYINPUT30), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT67), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n558), .A2(new_n572), .A3(new_n559), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n561), .A2(new_n336), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n566), .B(new_n335), .C1(new_n568), .C2(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n449), .A2(G210), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n576), .B(KEYINPUT27), .Z(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT26), .B(G101), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n577), .B(new_n578), .Z(new_n579));
  NAND3_X1  g393(.A1(new_n574), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT31), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n574), .A2(KEYINPUT31), .A3(new_n575), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n558), .A2(new_n336), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n575), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n567), .A2(new_n335), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n246), .B1(new_n562), .B2(new_n564), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n585), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT71), .B(new_n585), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n579), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT72), .ZN(new_n599));
  OR3_X1    g413(.A1(new_n599), .A2(G472), .A3(G902), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(G472), .B2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(KEYINPUT73), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n596), .B1(new_n582), .B2(new_n583), .ZN(new_n605));
  INV_X1    g419(.A(new_n602), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n605), .A2(new_n606), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT29), .B1(new_n595), .B2(new_n579), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n574), .A2(new_n575), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n579), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n566), .B1(new_n568), .B2(new_n570), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(new_n336), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n575), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n594), .B1(new_n617), .B2(KEYINPUT28), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n579), .A2(KEYINPUT29), .ZN(new_n619));
  AOI21_X1  g433(.A(G902), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n611), .A2(KEYINPUT32), .B1(new_n621), .B2(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n545), .B1(new_n610), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n431), .A2(new_n433), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT97), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n509), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n444), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n306), .A4(new_n301), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n512), .A2(new_n623), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G101), .ZN(G3));
  INV_X1    g448(.A(new_n307), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n603), .A2(new_n607), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n598), .A2(new_n637), .A3(new_n292), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT100), .B1(new_n605), .B2(G902), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(G472), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n545), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n368), .A2(new_n373), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n378), .A3(new_n629), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n422), .A2(new_n423), .A3(new_n430), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n425), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT33), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n428), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n426), .A2(new_n648), .A3(new_n427), .A4(KEYINPUT33), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(G478), .A3(new_n292), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n509), .A2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n643), .A2(new_n645), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT34), .B(G104), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G6));
  AND2_X1   g471(.A1(new_n491), .A2(new_n508), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n437), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n645), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n635), .A2(new_n642), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n529), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n541), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n539), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n641), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n512), .A2(new_n632), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND3_X1  g486(.A1(new_n644), .A2(new_n378), .A3(new_n667), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n441), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n440), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n437), .A2(new_n658), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n610), .A2(new_n622), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n301), .A3(new_n680), .A4(new_n306), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  XOR2_X1   g496(.A(new_n676), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n635), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n375), .A2(new_n376), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  INV_X1    g502(.A(new_n378), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n658), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n437), .A2(new_n690), .A3(new_n668), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  INV_X1    g506(.A(new_n579), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n574), .B2(new_n575), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n292), .B1(new_n617), .B2(new_n579), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT102), .Z(new_n697));
  INV_X1    g511(.A(KEYINPUT32), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n605), .A2(new_n698), .A3(new_n606), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n610), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n688), .A2(new_n692), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n685), .A2(new_n686), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  INV_X1    g519(.A(new_n654), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n677), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n673), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n301), .A3(new_n680), .A4(new_n306), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n294), .A2(new_n295), .ZN(new_n711));
  INV_X1    g525(.A(new_n272), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n299), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(G902), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n306), .A3(new_n300), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n644), .A2(new_n378), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n654), .A2(new_n444), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n623), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  INV_X1    g535(.A(new_n715), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n623), .A2(new_n660), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND4_X1  g538(.A1(new_n628), .A2(new_n378), .A3(new_n644), .A4(new_n667), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n714), .A2(new_n306), .A3(new_n300), .A4(new_n629), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n680), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND3_X1  g543(.A1(new_n644), .A2(new_n437), .A3(new_n690), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n584), .B1(new_n579), .B2(new_n618), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n602), .B(KEYINPUT104), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(G472), .B1(new_n605), .B2(G902), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n544), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n654), .A2(new_n676), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT105), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n734), .A2(new_n735), .A3(new_n667), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n717), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NAND2_X1  g557(.A1(new_n687), .A2(new_n378), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n287), .A2(new_n745), .A3(new_n300), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n745), .B1(new_n287), .B2(new_n300), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n306), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n744), .B1(new_n748), .B2(KEYINPUT107), .ZN(new_n749));
  INV_X1    g563(.A(new_n274), .ZN(new_n750));
  INV_X1    g564(.A(new_n266), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n294), .B2(new_n295), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n750), .B1(new_n752), .B2(new_n271), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n291), .B1(new_n753), .B2(new_n292), .ZN(new_n754));
  INV_X1    g568(.A(new_n300), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT106), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n287), .A2(new_n745), .A3(new_n300), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n305), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n749), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT32), .B1(new_n598), .B2(new_n602), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT108), .B1(new_n762), .B2(new_n699), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n611), .A2(KEYINPUT32), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n698), .B1(new_n605), .B2(new_n606), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n621), .A2(G472), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n763), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n544), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n740), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT42), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n740), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(KEYINPUT42), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n749), .A2(new_n774), .A3(new_n623), .A4(new_n760), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n262), .ZN(G33));
  INV_X1    g591(.A(new_n678), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n749), .A2(new_n623), .A3(new_n778), .A4(new_n760), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  NAND2_X1  g594(.A1(G469), .A2(G902), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n286), .B2(KEYINPUT45), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n753), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n781), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n755), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT46), .B(new_n781), .C1(new_n782), .C2(new_n784), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n305), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n744), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n789), .A2(new_n683), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n658), .A2(new_n653), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(KEYINPUT43), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(KEYINPUT43), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n641), .B2(new_n667), .ZN(new_n797));
  AOI211_X1 g611(.A(KEYINPUT109), .B(new_n668), .C1(new_n636), .C2(new_n640), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT44), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n791), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n789), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n707), .A2(new_n544), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n378), .A3(new_n687), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT111), .B1(new_n809), .B2(new_n680), .ZN(new_n810));
  INV_X1    g624(.A(new_n680), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n790), .A2(new_n811), .A3(new_n812), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n807), .B(new_n814), .C1(new_n789), .C2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n377), .A2(new_n378), .A3(new_n718), .ZN(new_n819));
  INV_X1    g633(.A(new_n625), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n509), .A3(new_n444), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n375), .A2(new_n821), .A3(new_n376), .A4(new_n378), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n822), .A2(KEYINPUT114), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n635), .B(new_n642), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n633), .A2(new_n670), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n730), .B1(new_n700), .B2(new_n610), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n667), .A2(new_n676), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n306), .B(new_n829), .C1(new_n746), .C2(new_n747), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT115), .B1(new_n758), .B2(new_n829), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n681), .A2(new_n742), .A3(new_n709), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT52), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n790), .B1(new_n758), .B2(new_n759), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n740), .A2(new_n741), .ZN(new_n838));
  AOI211_X1 g652(.A(KEYINPUT107), .B(new_n305), .C1(new_n756), .C2(new_n757), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n727), .A2(new_n680), .B1(new_n731), .B2(new_n736), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n676), .B1(new_n539), .B2(new_n666), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n820), .A2(new_n658), .A3(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n689), .B(new_n843), .C1(new_n375), .C2(new_n376), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n301), .A3(new_n680), .A4(new_n306), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n841), .A2(new_n719), .A3(new_n845), .A4(new_n723), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n840), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n835), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n830), .A2(new_n831), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n758), .A2(KEYINPUT115), .A3(new_n829), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n828), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n848), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n827), .A2(new_n836), .A3(new_n847), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n772), .A2(new_n775), .A3(new_n779), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n818), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n835), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n848), .B2(new_n852), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n772), .A2(new_n775), .A3(new_n779), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n719), .A2(new_n728), .A3(new_n723), .A4(new_n737), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n845), .C1(new_n838), .C2(new_n761), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n633), .A2(new_n670), .A3(new_n826), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n742), .A2(new_n681), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n818), .B1(new_n865), .B2(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n859), .A2(new_n860), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n856), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT116), .B1(new_n868), .B2(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n865), .B2(KEYINPUT52), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n856), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT116), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n856), .A2(new_n867), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n869), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n793), .A2(new_n794), .A3(new_n440), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n744), .A2(new_n715), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n770), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n881));
  NOR2_X1   g695(.A1(KEYINPUT120), .A2(KEYINPUT48), .ZN(new_n882));
  OR3_X1    g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(new_n881), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n701), .A2(new_n545), .A3(new_n440), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n706), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n268), .A2(G952), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n878), .A2(new_n736), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n887), .B1(new_n888), .B2(new_n717), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n883), .A2(new_n884), .A3(new_n886), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n879), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n509), .A3(new_n653), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n879), .A2(new_n741), .A3(new_n878), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT119), .Z(new_n894));
  OAI21_X1  g708(.A(new_n807), .B1(new_n789), .B2(new_n815), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n714), .A2(new_n300), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n306), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n888), .A2(new_n790), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n892), .B(new_n894), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n715), .A2(new_n378), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n888), .A2(new_n688), .A3(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n888), .A2(KEYINPUT117), .A3(new_n688), .A4(new_n900), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(KEYINPUT118), .A3(new_n904), .A4(new_n905), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n908), .B(new_n909), .C1(new_n904), .C2(new_n901), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n899), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT51), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n890), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n912), .B2(new_n911), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n877), .A2(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n545), .A2(new_n792), .A3(new_n305), .A4(new_n689), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT112), .Z(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(KEYINPUT49), .B2(new_n896), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(KEYINPUT49), .B2(new_n896), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n688), .A3(new_n702), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT113), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n921), .ZN(G75));
  AOI21_X1  g736(.A(new_n292), .B1(new_n856), .B2(new_n867), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G210), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n347), .A2(new_n349), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT121), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n369), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n268), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n926), .A2(new_n930), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G51));
  XOR2_X1   g750(.A(new_n781), .B(KEYINPUT57), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n875), .B1(new_n856), .B2(new_n867), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n713), .B(KEYINPUT122), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n782), .A2(new_n784), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n923), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n932), .B1(new_n942), .B2(new_n944), .ZN(G54));
  AND2_X1   g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n923), .A2(new_n501), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n501), .B1(new_n923), .B2(new_n946), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n932), .ZN(G60));
  NAND2_X1  g763(.A1(new_n650), .A2(new_n651), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(G478), .A2(G902), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT59), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n877), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n951), .B(new_n953), .C1(new_n938), .C2(new_n939), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n933), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n954), .A2(new_n956), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT60), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n868), .A2(new_n665), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n959), .B1(new_n856), .B2(new_n867), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n961), .B(new_n933), .C1(new_n543), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(KEYINPUT123), .A3(new_n933), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n964), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n962), .A2(new_n543), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n932), .B1(new_n962), .B2(new_n665), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n966), .B(new_n967), .C1(KEYINPUT123), .C2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n965), .A2(new_n969), .ZN(G66));
  NAND2_X1  g784(.A1(new_n827), .A2(new_n861), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n268), .ZN(new_n972));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n442), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(KEYINPUT124), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(KEYINPUT124), .B2(new_n972), .ZN(new_n976));
  INV_X1    g790(.A(G898), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n928), .B1(new_n977), .B2(G953), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G69));
  NAND2_X1  g793(.A1(G227), .A2(G900), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n803), .A2(new_n848), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n803), .A2(new_n983), .A3(new_n848), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n730), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n789), .A2(new_n770), .A3(new_n683), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n816), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n855), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(KEYINPUT127), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n803), .A2(new_n983), .A3(new_n848), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n983), .B1(new_n803), .B2(new_n848), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n989), .B(KEYINPUT127), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n268), .B1(new_n990), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n674), .A2(G953), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT125), .Z(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n573), .A2(new_n571), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n572), .B1(new_n558), .B2(new_n559), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(new_n493), .ZN(new_n1002));
  OAI211_X1 g816(.A(G953), .B(new_n980), .C1(new_n998), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n980), .A2(G953), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n704), .A2(new_n848), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT62), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n820), .A2(new_n509), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n790), .B(new_n623), .C1(new_n706), .C2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n803), .B(new_n816), .C1(new_n684), .C2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1002), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  INV_X1    g825(.A(new_n997), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n993), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1012), .B1(new_n1016), .B2(new_n268), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1004), .B(new_n1011), .C1(new_n1017), .C2(new_n1002), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1003), .A2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(G472), .A2(G902), .ZN(new_n1020));
  XOR2_X1   g834(.A(new_n1020), .B(KEYINPUT63), .Z(new_n1021));
  INV_X1    g835(.A(new_n580), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n613), .A2(new_n579), .ZN(new_n1023));
  OAI211_X1 g837(.A(new_n872), .B(new_n1021), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1021), .ZN(new_n1025));
  INV_X1    g839(.A(new_n971), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n1010), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n694), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n933), .B(new_n1024), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n613), .A2(new_n693), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1015), .A2(new_n1026), .A3(new_n993), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1021), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1029), .A2(new_n1032), .ZN(G57));
endmodule


