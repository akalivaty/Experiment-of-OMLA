

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X2 U552 ( .A(n599), .Z(n517) );
  XNOR2_X1 U553 ( .A(KEYINPUT69), .B(n543), .ZN(n599) );
  INV_X1 U554 ( .A(KEYINPUT103), .ZN(n709) );
  XNOR2_X1 U555 ( .A(n730), .B(KEYINPUT104), .ZN(n734) );
  NAND2_X1 U556 ( .A1(n890), .A2(G137), .ZN(n524) );
  XNOR2_X2 U557 ( .A(KEYINPUT70), .B(n551), .ZN(n589) );
  AND2_X1 U558 ( .A1(n695), .A2(n694), .ZN(n518) );
  AND2_X1 U559 ( .A1(n731), .A2(G8), .ZN(n519) );
  NOR2_X1 U560 ( .A1(n742), .A2(n745), .ZN(n520) );
  INV_X1 U561 ( .A(n992), .ZN(n696) );
  NAND2_X1 U562 ( .A1(n696), .A2(n695), .ZN(n687) );
  NOR2_X1 U563 ( .A1(n698), .A2(n697), .ZN(n699) );
  INV_X1 U564 ( .A(n736), .ZN(n718) );
  XNOR2_X1 U565 ( .A(n710), .B(n709), .ZN(n716) );
  OR2_X1 U566 ( .A1(n735), .A2(n742), .ZN(n730) );
  XNOR2_X1 U567 ( .A(n748), .B(KEYINPUT32), .ZN(n749) );
  NOR2_X1 U568 ( .A1(n732), .A2(n519), .ZN(n733) );
  INV_X1 U569 ( .A(KEYINPUT107), .ZN(n753) );
  XNOR2_X1 U570 ( .A(n754), .B(n753), .ZN(n801) );
  INV_X1 U571 ( .A(KEYINPUT79), .ZN(n583) );
  NAND2_X1 U572 ( .A1(n685), .A2(n775), .ZN(n736) );
  XNOR2_X1 U573 ( .A(n583), .B(KEYINPUT12), .ZN(n584) );
  XNOR2_X1 U574 ( .A(n585), .B(n584), .ZN(n587) );
  INV_X1 U575 ( .A(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n643) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n530), .ZN(n895) );
  AND2_X1 U578 ( .A1(n533), .A2(n532), .ZN(G160) );
  NOR2_X2 U579 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U580 ( .A(n522), .B(n521), .ZN(n890) );
  INV_X1 U581 ( .A(G2105), .ZN(n530) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U583 ( .A1(G113), .A2(n894), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U585 ( .A(n525), .B(KEYINPUT67), .ZN(n529) );
  XOR2_X1 U586 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n527) );
  AND2_X1 U587 ( .A1(n530), .A2(G2104), .ZN(n891) );
  NAND2_X1 U588 ( .A1(G101), .A2(n891), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n527), .B(n526), .ZN(n528) );
  AND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U591 ( .A1(G125), .A2(n895), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n531), .Z(n532) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U594 ( .A1(G135), .A2(n890), .ZN(n535) );
  NAND2_X1 U595 ( .A1(G111), .A2(n894), .ZN(n534) );
  NAND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n895), .A2(G123), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT18), .B(n536), .Z(n537) );
  NOR2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n540) );
  NAND2_X1 U600 ( .A1(n891), .A2(G99), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n943) );
  XNOR2_X1 U602 ( .A(G2096), .B(n943), .ZN(n541) );
  OR2_X1 U603 ( .A1(G2100), .A2(n541), .ZN(G156) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  NAND2_X1 U606 ( .A1(G90), .A2(n643), .ZN(n545) );
  INV_X1 U607 ( .A(G651), .ZN(n549) );
  XOR2_X1 U608 ( .A(G543), .B(KEYINPUT0), .Z(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT68), .B(n542), .ZN(n655) );
  OR2_X1 U610 ( .A1(n549), .A2(n655), .ZN(n543) );
  NAND2_X1 U611 ( .A1(G77), .A2(n517), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT9), .ZN(n548) );
  NOR2_X2 U614 ( .A1(G651), .A2(n655), .ZN(n649) );
  NAND2_X1 U615 ( .A1(G52), .A2(n649), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n554) );
  NOR2_X1 U617 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT1), .B(n550), .Z(n551) );
  NAND2_X1 U619 ( .A1(n589), .A2(G64), .ZN(n552) );
  XOR2_X1 U620 ( .A(KEYINPUT72), .B(n552), .Z(n553) );
  NOR2_X1 U621 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U622 ( .A1(G138), .A2(n890), .ZN(n556) );
  NAND2_X1 U623 ( .A1(G102), .A2(n891), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G114), .A2(n894), .ZN(n558) );
  NAND2_X1 U626 ( .A1(G126), .A2(n895), .ZN(n557) );
  NAND2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(G164) );
  NAND2_X1 U629 ( .A1(n649), .A2(G53), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT74), .B(n561), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G65), .A2(n589), .ZN(n562) );
  XOR2_X1 U632 ( .A(KEYINPUT73), .B(n562), .Z(n563) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(KEYINPUT75), .B(n565), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G91), .A2(n643), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G78), .A2(n517), .ZN(n566) );
  AND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G299) );
  NAND2_X1 U639 ( .A1(G89), .A2(n643), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT4), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT82), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G76), .A2(n517), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT5), .ZN(n579) );
  NAND2_X1 U645 ( .A1(n649), .A2(G51), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G63), .A2(n589), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT6), .B(n577), .Z(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U650 ( .A(n580), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U651 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n581), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U654 ( .A(G223), .ZN(n837) );
  NAND2_X1 U655 ( .A1(n837), .A2(G567), .ZN(n582) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  XOR2_X1 U657 ( .A(G860), .B(KEYINPUT80), .Z(n610) );
  NAND2_X1 U658 ( .A1(G81), .A2(n643), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G68), .A2(n517), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U661 ( .A(KEYINPUT13), .B(n588), .Z(n594) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n591) );
  NAND2_X1 U663 ( .A1(G56), .A2(n589), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n591), .B(n590), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT77), .B(n592), .Z(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n649), .A2(G43), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n992) );
  OR2_X1 U669 ( .A1(n610), .A2(n992), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(n649), .A2(G54), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G66), .A2(n589), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n603) );
  NAND2_X1 U674 ( .A1(G92), .A2(n643), .ZN(n601) );
  NAND2_X1 U675 ( .A1(G79), .A2(n517), .ZN(n600) );
  NAND2_X1 U676 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U678 ( .A(n604), .B(KEYINPUT15), .ZN(n997) );
  NOR2_X1 U679 ( .A1(n694), .A2(G868), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT81), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(G284) );
  NOR2_X1 U683 ( .A1(G868), .A2(G299), .ZN(n609) );
  INV_X1 U684 ( .A(G868), .ZN(n666) );
  NOR2_X1 U685 ( .A1(G286), .A2(n666), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n609), .A2(n608), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n611), .A2(n694), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G559), .A2(n666), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n694), .A2(n613), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT83), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n992), .A2(G868), .ZN(n615) );
  NOR2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G93), .A2(n643), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G67), .A2(n589), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n517), .A2(G80), .ZN(n619) );
  XOR2_X1 U699 ( .A(KEYINPUT84), .B(n619), .Z(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n649), .A2(G55), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n665) );
  NAND2_X1 U703 ( .A1(G559), .A2(n694), .ZN(n624) );
  XNOR2_X1 U704 ( .A(n992), .B(n624), .ZN(n663) );
  NOR2_X1 U705 ( .A1(G860), .A2(n663), .ZN(n625) );
  XOR2_X1 U706 ( .A(n665), .B(n625), .Z(G145) );
  NAND2_X1 U707 ( .A1(G86), .A2(n643), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G61), .A2(n589), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n517), .A2(G73), .ZN(n628) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n628), .Z(n629) );
  NOR2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n649), .A2(G48), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U715 ( .A1(n649), .A2(G50), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT87), .B(n633), .Z(n635) );
  NAND2_X1 U717 ( .A1(G62), .A2(n589), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U719 ( .A(KEYINPUT88), .B(n636), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G88), .A2(n643), .ZN(n638) );
  NAND2_X1 U721 ( .A1(G75), .A2(n517), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U723 ( .A1(n640), .A2(n639), .ZN(G166) );
  NAND2_X1 U724 ( .A1(G72), .A2(n517), .ZN(n642) );
  NAND2_X1 U725 ( .A1(G47), .A2(n649), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G85), .A2(n643), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G60), .A2(n589), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U730 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT71), .ZN(G290) );
  NAND2_X1 U732 ( .A1(n649), .A2(G49), .ZN(n650) );
  XOR2_X1 U733 ( .A(KEYINPUT85), .B(n650), .Z(n652) );
  NAND2_X1 U734 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U736 ( .A(KEYINPUT86), .B(n653), .ZN(n654) );
  NOR2_X1 U737 ( .A1(n589), .A2(n654), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(G288) );
  XNOR2_X1 U740 ( .A(G305), .B(KEYINPUT19), .ZN(n659) );
  INV_X1 U741 ( .A(G299), .ZN(n985) );
  XNOR2_X1 U742 ( .A(G166), .B(n985), .ZN(n658) );
  XNOR2_X1 U743 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U745 ( .A(n661), .B(n665), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(G288), .ZN(n907) );
  XOR2_X1 U747 ( .A(n663), .B(n907), .Z(n664) );
  NAND2_X1 U748 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2084), .A2(G2078), .ZN(n669) );
  XNOR2_X1 U752 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT89), .B(n670), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(KEYINPUT90), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n673) );
  XNOR2_X1 U757 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G2072), .A2(n675), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U760 ( .A(KEYINPUT76), .B(G132), .Z(G219) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U762 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U763 ( .A1(G108), .A2(n677), .ZN(n841) );
  NAND2_X1 U764 ( .A1(n841), .A2(G567), .ZN(n683) );
  NOR2_X1 U765 ( .A1(G219), .A2(G220), .ZN(n678) );
  XNOR2_X1 U766 ( .A(KEYINPUT22), .B(n678), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n679), .A2(G96), .ZN(n680) );
  NOR2_X1 U768 ( .A1(G218), .A2(n680), .ZN(n681) );
  XOR2_X1 U769 ( .A(KEYINPUT92), .B(n681), .Z(n842) );
  NAND2_X1 U770 ( .A1(G2106), .A2(n842), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n843) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U773 ( .A1(n843), .A2(n684), .ZN(n840) );
  NAND2_X1 U774 ( .A1(n840), .A2(G36), .ZN(G176) );
  XNOR2_X1 U775 ( .A(KEYINPUT93), .B(G166), .ZN(G303) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n774) );
  INV_X1 U777 ( .A(n774), .ZN(n685) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NAND2_X1 U779 ( .A1(G8), .A2(n736), .ZN(n811) );
  NAND2_X1 U780 ( .A1(n718), .A2(G1996), .ZN(n686) );
  XOR2_X1 U781 ( .A(n686), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U782 ( .A1(G1341), .A2(n736), .ZN(n695) );
  NOR2_X1 U783 ( .A1(n698), .A2(n687), .ZN(n692) );
  NAND2_X1 U784 ( .A1(n718), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U785 ( .A(n688), .B(KEYINPUT27), .ZN(n711) );
  XOR2_X1 U786 ( .A(G1956), .B(KEYINPUT100), .Z(n1009) );
  NOR2_X1 U787 ( .A1(n718), .A2(n1009), .ZN(n712) );
  INV_X1 U788 ( .A(n712), .ZN(n689) );
  NAND2_X1 U789 ( .A1(n985), .A2(n689), .ZN(n690) );
  OR2_X1 U790 ( .A1(n711), .A2(n690), .ZN(n704) );
  INV_X1 U791 ( .A(n704), .ZN(n691) );
  NOR2_X1 U792 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U793 ( .A1(n997), .A2(n693), .ZN(n708) );
  INV_X1 U794 ( .A(n997), .ZN(n694) );
  NAND2_X1 U795 ( .A1(n518), .A2(n696), .ZN(n697) );
  XNOR2_X1 U796 ( .A(n699), .B(KEYINPUT101), .ZN(n706) );
  AND2_X1 U797 ( .A1(n718), .A2(G2067), .ZN(n700) );
  XOR2_X1 U798 ( .A(n700), .B(KEYINPUT102), .Z(n702) );
  NAND2_X1 U799 ( .A1(n736), .A2(G1348), .ZN(n701) );
  NAND2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n703) );
  AND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n712), .ZN(n713) );
  OR2_X1 U805 ( .A1(n985), .A2(n713), .ZN(n714) );
  XNOR2_X1 U806 ( .A(KEYINPUT28), .B(n714), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U808 ( .A(n717), .B(KEYINPUT29), .ZN(n722) );
  XOR2_X1 U809 ( .A(G2078), .B(KEYINPUT25), .Z(n965) );
  NOR2_X1 U810 ( .A1(n965), .A2(n736), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n718), .A2(G1961), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n723) );
  NOR2_X1 U813 ( .A1(G301), .A2(n723), .ZN(n721) );
  NOR2_X1 U814 ( .A1(n722), .A2(n721), .ZN(n735) );
  AND2_X1 U815 ( .A1(G301), .A2(n723), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n811), .ZN(n732) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n736), .ZN(n731) );
  NOR2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n724) );
  NAND2_X1 U819 ( .A1(G8), .A2(n724), .ZN(n725) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n725), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G168), .A2(n726), .ZN(n727) );
  NOR2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n729), .B(KEYINPUT31), .ZN(n742) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n752) );
  INV_X1 U825 ( .A(n735), .ZN(n743) );
  INV_X1 U826 ( .A(G8), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n811), .ZN(n738) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n739), .A2(G303), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n745) );
  NAND2_X1 U832 ( .A1(n743), .A2(n520), .ZN(n747) );
  AND2_X1 U833 ( .A1(G286), .A2(G8), .ZN(n744) );
  OR2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n750) );
  XOR2_X1 U836 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n748) );
  XNOR2_X1 U837 ( .A(n750), .B(n749), .ZN(n751) );
  NAND2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n754) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U841 ( .A1(n981), .A2(n755), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n801), .A2(n756), .ZN(n757) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NAND2_X1 U844 ( .A1(n757), .A2(n983), .ZN(n758) );
  NOR2_X2 U845 ( .A1(n811), .A2(n758), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT64), .ZN(n760) );
  NOR2_X1 U847 ( .A1(KEYINPUT33), .A2(n760), .ZN(n763) );
  NAND2_X1 U848 ( .A1(n981), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n761), .A2(n811), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n799) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n978) );
  NAND2_X1 U852 ( .A1(G140), .A2(n890), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G104), .A2(n891), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U855 ( .A(KEYINPUT34), .B(n766), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G116), .A2(n894), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G128), .A2(n895), .ZN(n767) );
  NAND2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U859 ( .A(n769), .B(KEYINPUT35), .Z(n770) );
  NOR2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U861 ( .A(KEYINPUT36), .B(n772), .Z(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT94), .B(n773), .Z(n887) );
  XNOR2_X1 U863 ( .A(G2067), .B(KEYINPUT37), .ZN(n828) );
  NOR2_X1 U864 ( .A1(n887), .A2(n828), .ZN(n934) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n830) );
  NAND2_X1 U866 ( .A1(n934), .A2(n830), .ZN(n776) );
  XOR2_X1 U867 ( .A(KEYINPUT95), .B(n776), .Z(n826) );
  INV_X1 U868 ( .A(n826), .ZN(n796) );
  NAND2_X1 U869 ( .A1(G107), .A2(n894), .ZN(n778) );
  NAND2_X1 U870 ( .A1(G119), .A2(n895), .ZN(n777) );
  NAND2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U872 ( .A(KEYINPUT96), .B(n779), .Z(n783) );
  NAND2_X1 U873 ( .A1(G131), .A2(n890), .ZN(n781) );
  NAND2_X1 U874 ( .A1(G95), .A2(n891), .ZN(n780) );
  AND2_X1 U875 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n783), .A2(n782), .ZN(n877) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n877), .ZN(n784) );
  XNOR2_X1 U878 ( .A(n784), .B(KEYINPUT97), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G141), .A2(n890), .ZN(n785) );
  XNOR2_X1 U880 ( .A(n785), .B(KEYINPUT98), .ZN(n792) );
  NAND2_X1 U881 ( .A1(G117), .A2(n894), .ZN(n787) );
  NAND2_X1 U882 ( .A1(G129), .A2(n895), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n891), .A2(G105), .ZN(n788) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n886) );
  AND2_X1 U888 ( .A1(G1996), .A2(n886), .ZN(n793) );
  NOR2_X1 U889 ( .A1(n794), .A2(n793), .ZN(n940) );
  INV_X1 U890 ( .A(n830), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n940), .A2(n795), .ZN(n822) );
  NOR2_X1 U892 ( .A1(n796), .A2(n822), .ZN(n817) );
  AND2_X1 U893 ( .A1(n978), .A2(n817), .ZN(n797) );
  XNOR2_X1 U894 ( .A(G1986), .B(G290), .ZN(n994) );
  NAND2_X1 U895 ( .A1(n994), .A2(n830), .ZN(n800) );
  AND2_X1 U896 ( .A1(n797), .A2(n800), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n835) );
  INV_X1 U898 ( .A(n800), .ZN(n819) );
  INV_X1 U899 ( .A(n801), .ZN(n809) );
  NOR2_X1 U900 ( .A1(G2090), .A2(G303), .ZN(n802) );
  NAND2_X1 U901 ( .A1(G8), .A2(n802), .ZN(n803) );
  XOR2_X1 U902 ( .A(KEYINPUT108), .B(n803), .Z(n807) );
  NOR2_X1 U903 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XNOR2_X1 U904 ( .A(n804), .B(KEYINPUT24), .ZN(n805) );
  XNOR2_X1 U905 ( .A(n805), .B(KEYINPUT99), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n806), .A2(n811), .ZN(n810) );
  OR2_X1 U907 ( .A1(n807), .A2(n810), .ZN(n808) );
  NOR2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n815) );
  INV_X1 U909 ( .A(n810), .ZN(n813) );
  INV_X1 U910 ( .A(n811), .ZN(n812) );
  AND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n833) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n886), .ZN(n937) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n877), .ZN(n942) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n942), .A2(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U920 ( .A(KEYINPUT109), .B(n823), .Z(n824) );
  NOR2_X1 U921 ( .A1(n937), .A2(n824), .ZN(n825) );
  XNOR2_X1 U922 ( .A(KEYINPUT39), .B(n825), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n887), .A2(n828), .ZN(n933) );
  NAND2_X1 U925 ( .A1(n829), .A2(n933), .ZN(n831) );
  AND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(G188) );
  NOR2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G325) );
  XOR2_X1 U936 ( .A(KEYINPUT112), .B(G325), .Z(G261) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  INV_X1 U941 ( .A(n843), .ZN(G319) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2084), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2078), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n846), .B(G2100), .Z(n848) );
  XNOR2_X1 U946 ( .A(G2090), .B(G2072), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT113), .B(G2678), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(G227) );
  XNOR2_X1 U952 ( .A(G1976), .B(G2474), .ZN(n862) );
  XOR2_X1 U953 ( .A(G1956), .B(G1961), .Z(n854) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1971), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U956 ( .A(G1981), .B(G1966), .Z(n856) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U960 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U963 ( .A1(G124), .A2(n895), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n894), .A2(G112), .ZN(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G136), .A2(n890), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G100), .A2(n891), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G118), .A2(n894), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G130), .A2(n895), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G142), .A2(n890), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G106), .A2(n891), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(n874), .B(KEYINPUT45), .Z(n875) );
  NOR2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n885) );
  XOR2_X1 U980 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n943), .B(n881), .ZN(n883) );
  XNOR2_X1 U984 ( .A(G164), .B(G162), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U986 ( .A(n885), .B(n884), .Z(n889) );
  XOR2_X1 U987 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n903) );
  NAND2_X1 U989 ( .A1(G139), .A2(n890), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G103), .A2(n891), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G115), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G127), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U997 ( .A(KEYINPUT115), .B(n901), .ZN(n928) );
  XNOR2_X1 U998 ( .A(n928), .B(G160), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n992), .B(KEYINPUT118), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(G171), .B(n694), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n907), .B(G286), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  XNOR2_X1 U1007 ( .A(G2427), .B(KEYINPUT110), .ZN(n920) );
  XOR2_X1 U1008 ( .A(G2430), .B(G2446), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G2435), .B(G2438), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1011 ( .A(G2454), .B(KEYINPUT111), .Z(n914) );
  XNOR2_X1 U1012 ( .A(G1348), .B(G1341), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(n916), .B(n915), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G2451), .B(G2443), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n920), .B(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n921), .A2(G14), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n927), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n922), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(G395), .A2(G397), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1025 ( .A(G225), .ZN(G308) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(n927), .ZN(G401) );
  XNOR2_X1 U1028 ( .A(G164), .B(G2078), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(G2072), .B(KEYINPUT119), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(n932), .B(KEYINPUT50), .ZN(n950) );
  INV_X1 U1033 ( .A(n933), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n948) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n938), .Z(n939) );
  NAND2_X1 U1038 ( .A1(n940), .A2(n939), .ZN(n946) );
  XOR2_X1 U1039 ( .A(G160), .B(G2084), .Z(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1046 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n974), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n953), .A2(G29), .ZN(n1036) );
  XOR2_X1 U1049 ( .A(G34), .B(KEYINPUT122), .Z(n955) );
  XNOR2_X1 U1050 ( .A(G2084), .B(KEYINPUT54), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n955), .B(n954), .ZN(n972) );
  XNOR2_X1 U1052 ( .A(G2090), .B(G35), .ZN(n970) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G1991), .B(G25), .Z(n958) );
  NAND2_X1 U1057 ( .A1(n958), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(n959), .B(KEYINPUT120), .ZN(n962) );
  XOR2_X1 U1059 ( .A(G2067), .B(G26), .Z(n960) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(n960), .ZN(n961) );
  NOR2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G27), .B(n965), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1069 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n977), .ZN(n1034) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XNOR2_X1 U1073 ( .A(G168), .B(G1966), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(n980), .B(KEYINPUT57), .ZN(n1004) );
  INV_X1 U1076 ( .A(n981), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT125), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(n985), .B(G1956), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT124), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G303), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT126), .B(n991), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(G1341), .B(n992), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G1348), .B(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G301), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT123), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1032) );
  INV_X1 U1095 ( .A(G16), .ZN(n1030) );
  XNOR2_X1 U1096 ( .A(KEYINPUT127), .B(G1981), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G6), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .Z(n1008) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1008), .ZN(n1011) );
  XOR2_X1 U1100 ( .A(n1009), .B(G20), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G19), .B(G1341), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1016), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G21), .B(G1966), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1028), .ZN(n1029) );
  NAND2_X1 U1118 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1037), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

