//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202));
  AOI22_X1  g001(.A1(new_n202), .A2(KEYINPUT69), .B1(G211gat), .B2(G218gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n203), .B1(KEYINPUT69), .B2(new_n202), .ZN(new_n204));
  XNOR2_X1  g003(.A(G197gat), .B(G204gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT70), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n206), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n215), .A2(new_n216), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(G190gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G183gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n213), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n224), .A2(G183gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n222), .A2(G190gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n218), .A2(new_n220), .ZN(new_n231));
  AND2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n232), .B1(KEYINPUT23), .B2(new_n214), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT25), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G226gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n239), .A2(KEYINPUT26), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n239), .B(new_n241), .C1(new_n232), .C2(KEYINPUT26), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(new_n243), .B2(new_n214), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n222), .A2(new_n224), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n222), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT27), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(G183gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(new_n224), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n246), .B1(new_n250), .B2(KEYINPUT28), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n247), .A2(new_n249), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT28), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n224), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n235), .A2(new_n236), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n259), .B1(new_n235), .B2(new_n255), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n212), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n235), .A2(new_n236), .A3(new_n255), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n251), .A2(new_n254), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n245), .B1(new_n227), .B2(new_n234), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n211), .B(new_n262), .C1(new_n264), .C2(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(G64gat), .B(G92gat), .Z(new_n267));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n273));
  INV_X1    g072(.A(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n261), .A2(new_n265), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT73), .B1(new_n275), .B2(new_n273), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(KEYINPUT73), .A3(new_n273), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT76), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT66), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n286), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n284), .A2(G127gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(new_n287), .B2(KEYINPUT1), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(G120gat), .ZN(new_n296));
  INV_X1    g095(.A(G120gat), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(G113gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n299), .B(new_n286), .C1(new_n291), .C2(new_n289), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302));
  INV_X1    g101(.A(G155gat), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G148gat), .ZN(new_n309));
  INV_X1    g108(.A(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G141gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT74), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(new_n308), .A3(G148gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G141gat), .B(G148gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT2), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT4), .B1(new_n301), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n281), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n301), .A2(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n322), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT76), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n315), .B2(new_n320), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n301), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n334), .A3(new_n320), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT75), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n315), .A2(new_n320), .A3(new_n339), .A4(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n333), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n325), .A2(new_n330), .A3(new_n331), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(new_n341), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n344), .A2(new_n328), .A3(new_n332), .A4(new_n329), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n293), .A2(new_n321), .A3(new_n300), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n331), .B1(new_n347), .B2(new_n333), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(G57gat), .B(G85gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n353), .B1(new_n343), .B2(new_n349), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n349), .ZN(new_n359));
  INV_X1    g158(.A(new_n353), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n280), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G78gat), .B(G106gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n211), .B1(new_n341), .B2(new_n257), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n206), .A2(new_n210), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n209), .B1(new_n204), .B2(new_n205), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n257), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n322), .B1(new_n372), .B2(new_n334), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n368), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G22gat), .ZN(new_n375));
  AND2_X1   g174(.A1(new_n207), .A2(new_n208), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n204), .A2(new_n376), .A3(new_n205), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n204), .B2(new_n205), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT29), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n321), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n338), .B2(new_n340), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n380), .B(new_n367), .C1(new_n211), .C2(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n374), .A2(new_n375), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n374), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n366), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n382), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G22gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n374), .A2(new_n375), .A3(new_n382), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n366), .B(KEYINPUT77), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n383), .A2(new_n384), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT78), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n363), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT34), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n235), .A2(new_n255), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n301), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n235), .A2(new_n255), .A3(new_n300), .A4(new_n293), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G227gat), .ZN(new_n402));
  INV_X1    g201(.A(G233gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n397), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT34), .B(new_n404), .C1(new_n399), .C2(new_n400), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n399), .A2(new_n404), .A3(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT67), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(G71gat), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n413), .A2(KEYINPUT67), .ZN(new_n416));
  INV_X1    g215(.A(G71gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(KEYINPUT67), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G99gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n419), .A3(G99gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n410), .A2(new_n412), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n409), .B(KEYINPUT32), .C1(new_n411), .C2(new_n424), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT68), .B(new_n408), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n401), .A2(new_n405), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT34), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n401), .A2(new_n397), .A3(new_n405), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT68), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT68), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n406), .B2(new_n407), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n412), .A3(new_n425), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(new_n435), .A3(new_n427), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT36), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT36), .B1(new_n429), .B2(new_n437), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AND4_X1   g241(.A1(KEYINPUT78), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT78), .B1(new_n393), .B2(new_n389), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n385), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n325), .A2(new_n330), .A3(new_n344), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT39), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n333), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n353), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT39), .B1(new_n347), .B2(new_n333), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n447), .B2(new_n333), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n446), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n454), .A2(KEYINPUT40), .A3(new_n353), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n359), .A2(new_n360), .ZN(new_n456));
  INV_X1    g255(.A(new_n275), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT30), .ZN(new_n458));
  INV_X1    g257(.A(new_n279), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n458), .B(new_n272), .C1(new_n459), .C2(new_n277), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n453), .A2(new_n455), .A3(new_n456), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n456), .A2(new_n355), .A3(new_n354), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n361), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n261), .B2(new_n265), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT79), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT38), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n266), .A2(KEYINPUT37), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n261), .A2(new_n265), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n261), .A2(new_n265), .A3(KEYINPUT81), .A4(new_n472), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n271), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n275), .B1(new_n471), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n475), .A2(new_n476), .A3(new_n271), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(new_n469), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n464), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n396), .B(new_n442), .C1(new_n462), .C2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n392), .A2(new_n438), .A3(new_n394), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT35), .B1(new_n484), .B2(new_n363), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n460), .B1(new_n463), .B2(new_n361), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n445), .A2(new_n486), .A3(new_n487), .A4(new_n438), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT82), .ZN(new_n492));
  INV_X1    g291(.A(G29gat), .ZN(new_n493));
  INV_X1    g292(.A(G36gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT82), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n495), .A2(KEYINPUT14), .A3(new_n496), .ZN(new_n497));
  OAI22_X1  g296(.A1(new_n496), .A2(KEYINPUT14), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT15), .B(new_n491), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(KEYINPUT14), .A3(new_n496), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  INV_X1    g302(.A(G43gat), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(G50gat), .ZN(new_n505));
  INV_X1    g304(.A(G50gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(G43gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT83), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n497), .A2(new_n498), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(KEYINPUT83), .A3(new_n501), .A4(new_n508), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT84), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT84), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n516), .A3(new_n513), .ZN(new_n517));
  OR2_X1    g316(.A1(KEYINPUT89), .A2(G85gat), .ZN(new_n518));
  INV_X1    g317(.A(G92gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(KEYINPUT89), .A2(G85gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT8), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n525));
  AND2_X1   g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G106gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n421), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT90), .A3(new_n522), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G85gat), .A2(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT88), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT88), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(G85gat), .A3(G92gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT7), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n524), .A2(new_n532), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n528), .A2(new_n531), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n523), .A3(new_n521), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n541), .B1(new_n542), .B2(new_n537), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n543), .A3(KEYINPUT91), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n543), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n515), .A2(new_n517), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(G232gat), .A2(G233gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT41), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n511), .A2(new_n516), .A3(new_n513), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n516), .B1(new_n511), .B2(new_n513), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT17), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n547), .A2(new_n544), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n514), .A2(KEYINPUT17), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n548), .B(new_n550), .C1(new_n553), .C2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n557), .A2(KEYINPUT92), .ZN(new_n558));
  XNOR2_X1  g357(.A(G190gat), .B(G218gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n560), .B1(new_n557), .B2(KEYINPUT92), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n557), .A2(KEYINPUT92), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n559), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n560), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n574), .A2(new_n567), .A3(new_n566), .A4(new_n558), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n417), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G57gat), .A2(G64gat), .ZN(new_n580));
  OR2_X1    g379(.A1(G57gat), .A2(G64gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n417), .A2(new_n578), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT86), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n583), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n586), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(G127gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(G15gat), .B(G22gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT16), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(G1gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(G1gat), .B2(new_n594), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G8gat), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n585), .A2(KEYINPUT87), .A3(new_n587), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT87), .B1(new_n585), .B2(new_n587), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n593), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G155gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n603), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n576), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n547), .A2(new_n601), .A3(KEYINPUT10), .A4(new_n544), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n582), .B(new_n586), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n541), .A2(KEYINPUT94), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n545), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n613), .A2(new_n540), .A3(new_n543), .A4(new_n614), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n612), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT95), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n622), .A2(new_n625), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G229gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT85), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n515), .A2(new_n598), .A3(new_n517), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n597), .B(G8gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n555), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n636), .B(new_n637), .C1(new_n553), .C2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT18), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n638), .B1(new_n551), .B2(new_n552), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n637), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n636), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT17), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n515), .A2(new_n648), .A3(new_n517), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n598), .B1(new_n514), .B2(KEYINPUT17), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n651), .A2(KEYINPUT18), .A3(new_n636), .A4(new_n637), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n642), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G113gat), .B(G141gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G197gat), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT11), .B(G169gat), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT12), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n640), .A2(new_n641), .B1(new_n644), .B2(new_n646), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n658), .A3(new_n652), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n611), .A2(new_n634), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n490), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n464), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n280), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT97), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT97), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(G8gat), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT16), .B(G8gat), .Z(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n676), .B2(new_n677), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n678), .B(new_n680), .C1(new_n682), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g482(.A(new_n438), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n670), .A2(G15gat), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n670), .B2(new_n442), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n670), .A2(new_n445), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n466), .A2(new_n467), .ZN(new_n691));
  AOI211_X1 g490(.A(KEYINPUT79), .B(new_n465), .C1(new_n261), .C2(new_n265), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT38), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n457), .B1(new_n693), .B2(new_n480), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT38), .B1(new_n477), .B2(new_n466), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n361), .A3(new_n463), .A4(new_n695), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n696), .A2(new_n461), .A3(new_n445), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n684), .A2(KEYINPUT36), .ZN(new_n698));
  INV_X1    g497(.A(new_n441), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n698), .B(new_n699), .C1(new_n445), .C2(new_n486), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT100), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n392), .A2(new_n438), .A3(new_n394), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n487), .B1(new_n702), .B2(new_n486), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n484), .A2(new_n363), .A3(KEYINPUT35), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT101), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n485), .A2(new_n488), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n696), .A2(new_n461), .A3(new_n445), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n396), .A4(new_n442), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n701), .A2(new_n705), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n576), .A2(KEYINPUT44), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n570), .A2(new_n575), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n490), .A2(new_n713), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n711), .A2(new_n712), .B1(new_n714), .B2(KEYINPUT44), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n610), .A2(new_n664), .A3(new_n634), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT99), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n493), .B1(new_n719), .B2(new_n672), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n490), .A2(new_n713), .A3(new_n716), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n493), .A3(new_n672), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT98), .B(KEYINPUT45), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT102), .ZN(G1328gat));
  NAND3_X1  g525(.A1(new_n721), .A2(new_n494), .A3(new_n460), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT46), .Z(new_n728));
  NOR3_X1   g527(.A1(new_n715), .A2(new_n280), .A3(new_n718), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(KEYINPUT103), .ZN(new_n730));
  OAI21_X1  g529(.A(G36gat), .B1(new_n729), .B2(KEYINPUT103), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(G1329gat));
  NAND3_X1  g531(.A1(new_n721), .A2(new_n504), .A3(new_n438), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n715), .A2(new_n442), .A3(new_n718), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT47), .B(new_n733), .C1(new_n734), .C2(new_n504), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n734), .B2(new_n504), .ZN(new_n737));
  INV_X1    g536(.A(new_n442), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n711), .A2(new_n712), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n714), .A2(KEYINPUT44), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n738), .B(new_n717), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(KEYINPUT104), .A3(G43gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(new_n742), .A3(new_n733), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n735), .B1(new_n746), .B2(new_n747), .ZN(G1330gat));
  AOI21_X1  g547(.A(new_n506), .B1(new_n719), .B2(new_n395), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n395), .A2(new_n506), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT106), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n721), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g552(.A(new_n634), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n611), .A2(new_n754), .A3(new_n663), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT107), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n464), .B(KEYINPUT108), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n711), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g558(.A(new_n280), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n711), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n761), .B(new_n762), .Z(G1333gat));
  NAND4_X1  g562(.A1(new_n756), .A2(G71gat), .A3(new_n738), .A4(new_n711), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n438), .B(KEYINPUT109), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n756), .A2(new_n711), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n764), .B1(new_n766), .B2(G71gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g567(.A1(new_n756), .A2(new_n395), .A3(new_n711), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT110), .B(G78gat), .Z(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n610), .A2(new_n663), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT111), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n576), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n711), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(KEYINPUT51), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n634), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n518), .A2(new_n520), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n672), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n773), .A2(new_n754), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n715), .A2(new_n782), .A3(new_n464), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n780), .B2(new_n783), .ZN(G1336gat));
  NAND2_X1  g583(.A1(new_n460), .A2(new_n519), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n778), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n715), .A2(new_n782), .A3(new_n280), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n519), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(G92gat), .B1(new_n787), .B2(KEYINPUT112), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(KEYINPUT112), .B2(new_n787), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(G1337gat));
  AOI21_X1  g592(.A(G99gat), .B1(new_n779), .B2(new_n438), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n715), .A2(new_n782), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n442), .A2(new_n421), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(G1338gat));
  NAND2_X1  g596(.A1(new_n395), .A2(new_n529), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n715), .A2(new_n782), .A3(new_n445), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n778), .A2(new_n798), .B1(new_n799), .B2(new_n529), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n576), .A2(new_n610), .A3(new_n754), .A4(new_n664), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n612), .A2(new_n619), .A3(new_n624), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n622), .A2(new_n805), .A3(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n624), .B1(new_n612), .B2(new_n619), .ZN(new_n807));
  XOR2_X1   g606(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n808));
  AOI21_X1  g607(.A(new_n630), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n633), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n806), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n804), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n809), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n816), .A2(KEYINPUT114), .A3(new_n633), .A4(new_n810), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n813), .A2(new_n817), .A3(new_n663), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n551), .A2(new_n638), .A3(new_n552), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n649), .B2(new_n650), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n821), .A2(new_n636), .B1(new_n644), .B2(new_n646), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n819), .B1(new_n822), .B2(new_n657), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n636), .B1(new_n651), .B2(new_n637), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n644), .A2(new_n646), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n819), .B(new_n657), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n634), .B(new_n662), .C1(new_n823), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n576), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n657), .B1(new_n824), .B2(new_n825), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n642), .A2(new_n647), .A3(new_n652), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n832), .A2(new_n826), .B1(new_n833), .B2(new_n658), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n713), .A2(new_n813), .A3(new_n817), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n608), .A2(new_n609), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n803), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n757), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n702), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n460), .ZN(new_n842));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n663), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n672), .A2(new_n280), .ZN(new_n844));
  NOR4_X1   g643(.A1(new_n838), .A2(new_n395), .A3(new_n684), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n664), .A2(new_n295), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(G1340gat));
  NAND2_X1  g646(.A1(new_n634), .A2(new_n297), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT116), .Z(new_n849));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n845), .ZN(new_n851));
  OAI21_X1  g650(.A(G120gat), .B1(new_n851), .B2(new_n754), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n842), .A2(new_n854), .A3(new_n610), .ZN(new_n855));
  OAI21_X1  g654(.A(G127gat), .B1(new_n851), .B2(new_n837), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NOR2_X1   g656(.A1(new_n576), .A2(new_n460), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT117), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n841), .A2(G134gat), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n851), .B2(new_n576), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(KEYINPUT56), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(G1343gat));
  NOR2_X1   g663(.A1(new_n738), .A2(new_n445), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n840), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n460), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n663), .A2(new_n308), .ZN(new_n868));
  XOR2_X1   g667(.A(new_n868), .B(KEYINPUT118), .Z(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n738), .A2(new_n844), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n838), .B2(new_n445), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n834), .A2(new_n570), .A3(new_n575), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n813), .A2(new_n817), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n810), .A2(new_n633), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n653), .A2(new_n659), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n658), .B1(new_n661), .B2(new_n652), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n879), .B(new_n816), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n882), .A2(new_n828), .B1(new_n570), .B2(new_n575), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n837), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n802), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n445), .A2(new_n874), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n873), .B1(new_n875), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n308), .B1(new_n888), .B2(new_n663), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n871), .A2(KEYINPUT58), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT58), .B1(new_n871), .B2(new_n889), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n310), .A2(KEYINPUT59), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n888), .B2(new_n634), .ZN(new_n895));
  INV_X1    g694(.A(new_n886), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n811), .A2(new_n812), .ZN(new_n897));
  AND4_X1   g696(.A1(new_n575), .A2(new_n834), .A3(new_n897), .A4(new_n570), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n837), .B1(new_n898), .B2(new_n883), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n445), .B1(new_n899), .B2(new_n802), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n838), .A2(new_n896), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n872), .A2(new_n634), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n310), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT120), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n899), .A2(new_n802), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n395), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n713), .B1(new_n818), .B2(new_n828), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n837), .B1(new_n909), .B2(new_n878), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n896), .B1(new_n910), .B2(new_n802), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n903), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G148gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT59), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n895), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n867), .A2(new_n310), .A3(new_n634), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT121), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n875), .A2(new_n887), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n872), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n893), .B1(new_n921), .B2(new_n754), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n914), .B1(new_n913), .B2(KEYINPUT59), .ZN(new_n923));
  AOI211_X1 g722(.A(KEYINPUT120), .B(new_n905), .C1(new_n912), .C2(G148gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n917), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n919), .A2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n921), .B2(new_n837), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n867), .A2(new_n303), .A3(new_n610), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1346gat));
  AOI21_X1  g730(.A(new_n304), .B1(new_n888), .B2(new_n713), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n866), .A2(G162gat), .A3(new_n859), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(G1347gat));
  NOR2_X1   g733(.A1(new_n838), .A2(new_n672), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n484), .A2(new_n280), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(G169gat), .B1(new_n937), .B2(new_n663), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n757), .A2(new_n280), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n765), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT122), .Z(new_n941));
  NOR2_X1   g740(.A1(new_n838), .A2(new_n395), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n943), .A2(new_n237), .A3(new_n664), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n938), .A2(new_n944), .ZN(G1348gat));
  INV_X1    g744(.A(new_n943), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n946), .A2(G176gat), .A3(new_n634), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n634), .A3(new_n936), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT123), .A3(new_n238), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT123), .B1(new_n948), .B2(new_n238), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT124), .ZN(G1349gat));
  NAND3_X1  g751(.A1(new_n937), .A2(new_n252), .A3(new_n610), .ZN(new_n953));
  OAI21_X1  g752(.A(G183gat), .B1(new_n943), .B2(new_n837), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n937), .A2(new_n224), .A3(new_n713), .ZN(new_n957));
  OAI21_X1  g756(.A(G190gat), .B1(new_n943), .B2(new_n576), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1351gat));
  NOR3_X1   g760(.A1(new_n738), .A2(new_n280), .A3(new_n445), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n935), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n663), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n901), .B(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n442), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(G197gat), .A3(new_n663), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(G1352gat));
  NOR3_X1   g769(.A1(new_n963), .A2(G204gat), .A3(new_n754), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n966), .A2(new_n634), .A3(new_n968), .ZN(new_n973));
  INV_X1    g772(.A(G204gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n901), .A2(new_n610), .A3(new_n968), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G211gat), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  NOR3_X1   g777(.A1(new_n963), .A2(G211gat), .A3(new_n837), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT126), .Z(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1354gat));
  AOI21_X1  g780(.A(G218gat), .B1(new_n964), .B2(new_n713), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n966), .A2(new_n968), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n713), .A2(G218gat), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT127), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n982), .B1(new_n983), .B2(new_n985), .ZN(G1355gat));
endmodule


