

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U550 ( .A(n693), .B(n692), .ZN(n706) );
  NOR2_X2 U551 ( .A1(G1966), .A2(n777), .ZN(n738) );
  NOR2_X2 U552 ( .A1(n558), .A2(n557), .ZN(G160) );
  BUF_X1 U553 ( .A(n621), .Z(n622) );
  XNOR2_X2 U554 ( .A(n517), .B(n516), .ZN(n625) );
  XOR2_X1 U555 ( .A(KEYINPUT31), .B(n704), .Z(n513) );
  NOR2_X1 U556 ( .A1(n777), .A2(n761), .ZN(n514) );
  XOR2_X1 U557 ( .A(n698), .B(n697), .Z(n515) );
  XNOR2_X1 U558 ( .A(KEYINPUT93), .B(KEYINPUT30), .ZN(n697) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n712) );
  AND2_X1 U560 ( .A1(G160), .A2(G40), .ZN(n783) );
  INV_X1 U561 ( .A(KEYINPUT68), .ZN(n516) );
  NAND2_X1 U562 ( .A1(n625), .A2(G114), .ZN(n518) );
  AND2_X1 U563 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XNOR2_X1 U565 ( .A(n518), .B(KEYINPUT86), .ZN(n526) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n519), .Z(n621) );
  AND2_X1 U568 ( .A1(n621), .A2(G138), .ZN(n524) );
  INV_X1 U569 ( .A(G2104), .ZN(n520) );
  AND2_X2 U570 ( .A1(n520), .A2(G2105), .ZN(n872) );
  NAND2_X1 U571 ( .A1(G126), .A2(n872), .ZN(n522) );
  NOR2_X1 U572 ( .A1(G2105), .A2(n520), .ZN(n549) );
  BUF_X1 U573 ( .A(n549), .Z(n867) );
  NAND2_X1 U574 ( .A1(G102), .A2(n867), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U576 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT65), .B(n527), .Z(n647) );
  NAND2_X1 U579 ( .A1(G85), .A2(n647), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n641) );
  INV_X1 U581 ( .A(G651), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n641), .A2(n530), .ZN(n651) );
  NAND2_X1 U583 ( .A1(G72), .A2(n651), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n537) );
  NOR2_X1 U585 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n531), .Z(n532) );
  XNOR2_X1 U587 ( .A(KEYINPUT70), .B(n532), .ZN(n648) );
  NAND2_X1 U588 ( .A1(G60), .A2(n648), .ZN(n535) );
  NOR2_X1 U589 ( .A1(G651), .A2(n641), .ZN(n533) );
  XNOR2_X1 U590 ( .A(KEYINPUT66), .B(n533), .ZN(n656) );
  NAND2_X1 U591 ( .A1(G47), .A2(n656), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U593 ( .A1(n537), .A2(n536), .ZN(G290) );
  XOR2_X1 U594 ( .A(G2438), .B(G2454), .Z(n539) );
  XNOR2_X1 U595 ( .A(G2435), .B(G2430), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U597 ( .A(n540), .B(G2427), .Z(n542) );
  XNOR2_X1 U598 ( .A(G1341), .B(G1348), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n542), .B(n541), .ZN(n546) );
  XOR2_X1 U600 ( .A(G2443), .B(G2446), .Z(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT102), .B(G2451), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(n546), .B(n545), .Z(n547) );
  AND2_X1 U604 ( .A1(G14), .A2(n547), .ZN(G401) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U606 ( .A1(G125), .A2(n872), .ZN(n548) );
  XNOR2_X1 U607 ( .A(n548), .B(KEYINPUT67), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G101), .A2(n549), .ZN(n550) );
  XNOR2_X1 U609 ( .A(KEYINPUT23), .B(n550), .ZN(n551) );
  NOR2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n621), .A2(G137), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n558) );
  AND2_X1 U613 ( .A1(G113), .A2(n625), .ZN(n556) );
  INV_X1 U614 ( .A(KEYINPUT69), .ZN(n555) );
  XNOR2_X1 U615 ( .A(n556), .B(n555), .ZN(n557) );
  INV_X1 U616 ( .A(G108), .ZN(G238) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  NAND2_X1 U618 ( .A1(n656), .A2(G52), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n559), .B(KEYINPUT71), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G90), .A2(n647), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G77), .A2(n651), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U623 ( .A(n562), .B(KEYINPUT9), .ZN(n564) );
  NAND2_X1 U624 ( .A1(G64), .A2(n648), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U626 ( .A1(n566), .A2(n565), .ZN(G171) );
  INV_X1 U627 ( .A(G171), .ZN(G301) );
  NAND2_X1 U628 ( .A1(G88), .A2(n647), .ZN(n568) );
  NAND2_X1 U629 ( .A1(G75), .A2(n651), .ZN(n567) );
  NAND2_X1 U630 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT78), .B(n569), .Z(n573) );
  NAND2_X1 U632 ( .A1(n648), .A2(G62), .ZN(n571) );
  NAND2_X1 U633 ( .A1(n656), .A2(G50), .ZN(n570) );
  AND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n573), .A2(n572), .ZN(G303) );
  NAND2_X1 U636 ( .A1(n647), .A2(G89), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT4), .ZN(n576) );
  NAND2_X1 U638 ( .A1(G76), .A2(n651), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U640 ( .A(n577), .B(KEYINPUT5), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G63), .A2(n648), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G51), .A2(n656), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT6), .B(n580), .Z(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U646 ( .A(n583), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U647 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U648 ( .A1(G7), .A2(G661), .ZN(n584) );
  XOR2_X1 U649 ( .A(n584), .B(KEYINPUT10), .Z(n833) );
  AND2_X1 U650 ( .A1(G567), .A2(n833), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U652 ( .A1(n647), .A2(G81), .ZN(n586) );
  XNOR2_X1 U653 ( .A(n586), .B(KEYINPUT12), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G68), .A2(n651), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT13), .B(n589), .Z(n593) );
  NAND2_X1 U657 ( .A1(n648), .A2(G56), .ZN(n590) );
  XNOR2_X1 U658 ( .A(n590), .B(KEYINPUT14), .ZN(n591) );
  XNOR2_X1 U659 ( .A(n591), .B(KEYINPUT73), .ZN(n592) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G43), .A2(n656), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n724) );
  INV_X1 U663 ( .A(n724), .ZN(n957) );
  NAND2_X1 U664 ( .A1(n957), .A2(G860), .ZN(G153) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U666 ( .A1(G92), .A2(n647), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G79), .A2(n651), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G66), .A2(n648), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G54), .A2(n656), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(KEYINPUT15), .B(n602), .Z(n948) );
  OR2_X1 U674 ( .A1(n948), .A2(G868), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G65), .A2(n648), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G53), .A2(n656), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G91), .A2(n647), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G78), .A2(n651), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n715) );
  INV_X1 U683 ( .A(n715), .ZN(G299) );
  INV_X1 U684 ( .A(G868), .ZN(n670) );
  NOR2_X1 U685 ( .A1(G286), .A2(n670), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT74), .ZN(n613) );
  NOR2_X1 U687 ( .A1(G299), .A2(G868), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U689 ( .A(G860), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n614), .A2(G559), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n615), .A2(n948), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n724), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G868), .A2(n948), .ZN(n617) );
  NOR2_X1 U695 ( .A1(G559), .A2(n617), .ZN(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U697 ( .A1(n872), .A2(G123), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G135), .A2(n622), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G99), .A2(n867), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G111), .A2(n625), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n923) );
  XOR2_X1 U705 ( .A(n923), .B(G2096), .Z(n630) );
  INV_X1 U706 ( .A(G2100), .ZN(n894) );
  NAND2_X1 U707 ( .A1(n630), .A2(n894), .ZN(G156) );
  NAND2_X1 U708 ( .A1(n647), .A2(G93), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n631), .B(KEYINPUT76), .ZN(n633) );
  NAND2_X1 U710 ( .A1(G80), .A2(n651), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G67), .A2(n648), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G55), .A2(n656), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  OR2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n671) );
  NAND2_X1 U716 ( .A1(n948), .A2(G559), .ZN(n668) );
  XNOR2_X1 U717 ( .A(KEYINPUT75), .B(n957), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n668), .B(n638), .ZN(n639) );
  NOR2_X1 U719 ( .A1(G860), .A2(n639), .ZN(n640) );
  XOR2_X1 U720 ( .A(n671), .B(n640), .Z(G145) );
  NAND2_X1 U721 ( .A1(G87), .A2(n641), .ZN(n643) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n642) );
  NAND2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n648), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(G49), .A2(n656), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U727 ( .A1(G86), .A2(n647), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G61), .A2(n648), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G73), .A2(n651), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n653), .B(KEYINPUT77), .ZN(n654) );
  NOR2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G48), .A2(n656), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(G305) );
  XOR2_X1 U736 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n659) );
  XNOR2_X1 U737 ( .A(G288), .B(n659), .ZN(n660) );
  XOR2_X1 U738 ( .A(n660), .B(KEYINPUT81), .Z(n662) );
  XOR2_X1 U739 ( .A(G303), .B(KEYINPUT79), .Z(n661) );
  XNOR2_X1 U740 ( .A(n662), .B(n661), .ZN(n665) );
  XOR2_X1 U741 ( .A(n671), .B(n724), .Z(n663) );
  XNOR2_X1 U742 ( .A(n663), .B(G305), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(n667) );
  XOR2_X1 U744 ( .A(G290), .B(G299), .Z(n666) );
  XNOR2_X1 U745 ( .A(n667), .B(n666), .ZN(n884) );
  XNOR2_X1 U746 ( .A(n884), .B(n668), .ZN(n669) );
  NOR2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U748 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U749 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U754 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT22), .B(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G96), .ZN(n680) );
  NOR2_X1 U760 ( .A1(G218), .A2(n680), .ZN(n681) );
  XOR2_X1 U761 ( .A(KEYINPUT82), .B(n681), .Z(n839) );
  NAND2_X1 U762 ( .A1(n839), .A2(G2106), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n682), .B(KEYINPUT83), .ZN(n688) );
  NAND2_X1 U764 ( .A1(G120), .A2(G69), .ZN(n683) );
  XNOR2_X1 U765 ( .A(KEYINPUT84), .B(n683), .ZN(n684) );
  NOR2_X1 U766 ( .A1(G238), .A2(n684), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G57), .A2(n685), .ZN(n686) );
  XOR2_X1 U768 ( .A(KEYINPUT85), .B(n686), .Z(n840) );
  AND2_X1 U769 ( .A1(G567), .A2(n840), .ZN(n687) );
  NOR2_X1 U770 ( .A1(n688), .A2(n687), .ZN(G319) );
  INV_X1 U771 ( .A(G319), .ZN(n690) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U773 ( .A1(n690), .A2(n689), .ZN(n838) );
  NAND2_X1 U774 ( .A1(n838), .A2(G36), .ZN(G176) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n784) );
  AND2_X1 U776 ( .A1(n783), .A2(n784), .ZN(n693) );
  INV_X1 U777 ( .A(KEYINPUT64), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n706), .A2(G2084), .ZN(n694) );
  NAND2_X1 U779 ( .A1(G8), .A2(n694), .ZN(n741) );
  NAND2_X1 U780 ( .A1(n706), .A2(G8), .ZN(n777) );
  NOR2_X1 U781 ( .A1(n738), .A2(n694), .ZN(n695) );
  XNOR2_X1 U782 ( .A(n695), .B(KEYINPUT92), .ZN(n696) );
  NAND2_X1 U783 ( .A1(n696), .A2(G8), .ZN(n698) );
  NOR2_X1 U784 ( .A1(G168), .A2(n515), .ZN(n703) );
  XOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .Z(n1001) );
  INV_X1 U786 ( .A(n706), .ZN(n719) );
  NAND2_X1 U787 ( .A1(n1001), .A2(n719), .ZN(n700) );
  NAND2_X1 U788 ( .A1(n706), .A2(G1961), .ZN(n699) );
  NAND2_X1 U789 ( .A1(n700), .A2(n699), .ZN(n705) );
  NAND2_X1 U790 ( .A1(G301), .A2(n705), .ZN(n701) );
  XOR2_X1 U791 ( .A(KEYINPUT94), .B(n701), .Z(n702) );
  NOR2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U793 ( .A1(G301), .A2(n705), .ZN(n736) );
  INV_X1 U794 ( .A(G2072), .ZN(n998) );
  NOR2_X1 U795 ( .A1(n706), .A2(n998), .ZN(n708) );
  XOR2_X1 U796 ( .A(KEYINPUT27), .B(KEYINPUT89), .Z(n707) );
  XNOR2_X1 U797 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n706), .A2(G1956), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U800 ( .A(KEYINPUT90), .B(n711), .Z(n714) );
  NOR2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n713) );
  XNOR2_X1 U802 ( .A(n713), .B(n712), .ZN(n733) );
  NAND2_X1 U803 ( .A1(n715), .A2(n714), .ZN(n731) );
  NAND2_X1 U804 ( .A1(G2067), .A2(n719), .ZN(n717) );
  NAND2_X1 U805 ( .A1(n706), .A2(G1348), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U807 ( .A(KEYINPUT91), .B(n718), .ZN(n727) );
  OR2_X1 U808 ( .A1(n948), .A2(n727), .ZN(n726) );
  NAND2_X1 U809 ( .A1(n719), .A2(G1996), .ZN(n720) );
  XNOR2_X1 U810 ( .A(n720), .B(KEYINPUT26), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n706), .A2(G1341), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n727), .A2(n948), .ZN(n728) );
  AND2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U819 ( .A(KEYINPUT29), .B(n734), .Z(n735) );
  NAND2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n513), .A2(n737), .ZN(n743) );
  XNOR2_X1 U822 ( .A(KEYINPUT95), .B(n743), .ZN(n739) );
  NOR2_X1 U823 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n741), .A2(n740), .ZN(n756) );
  AND2_X1 U825 ( .A1(G286), .A2(G8), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n743), .A2(n742), .ZN(n752) );
  INV_X1 U827 ( .A(G8), .ZN(n750) );
  NOR2_X1 U828 ( .A1(n706), .A2(G2090), .ZN(n745) );
  XNOR2_X1 U829 ( .A(n745), .B(KEYINPUT96), .ZN(n747) );
  NOR2_X1 U830 ( .A1(n777), .A2(G1971), .ZN(n746) );
  NOR2_X1 U831 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U833 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U834 ( .A1(n752), .A2(n751), .ZN(n754) );
  XOR2_X1 U835 ( .A(KEYINPUT97), .B(KEYINPUT32), .Z(n753) );
  XNOR2_X1 U836 ( .A(n754), .B(n753), .ZN(n755) );
  NAND2_X1 U837 ( .A1(n756), .A2(n755), .ZN(n776) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U840 ( .A1(n952), .A2(n757), .ZN(n758) );
  NAND2_X1 U841 ( .A1(n776), .A2(n758), .ZN(n759) );
  XNOR2_X1 U842 ( .A(n759), .B(KEYINPUT98), .ZN(n766) );
  NAND2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n760) );
  XOR2_X1 U844 ( .A(KEYINPUT99), .B(n760), .Z(n945) );
  INV_X1 U845 ( .A(n945), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n952), .A2(KEYINPUT33), .ZN(n762) );
  NOR2_X1 U847 ( .A1(n762), .A2(n777), .ZN(n764) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n958) );
  INV_X1 U849 ( .A(n958), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n770) );
  AND2_X1 U851 ( .A1(n514), .A2(n770), .ZN(n765) );
  AND2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n782) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n767) );
  NAND2_X1 U854 ( .A1(G8), .A2(n767), .ZN(n774) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n768) );
  XOR2_X1 U856 ( .A(n768), .B(KEYINPUT24), .Z(n769) );
  OR2_X1 U857 ( .A1(n777), .A2(n769), .ZN(n772) );
  NAND2_X1 U858 ( .A1(n770), .A2(KEYINPUT33), .ZN(n771) );
  NAND2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n778) );
  INV_X1 U860 ( .A(n778), .ZN(n773) );
  AND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U862 ( .A1(n776), .A2(n775), .ZN(n780) );
  OR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  AND2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n812) );
  INV_X1 U866 ( .A(n783), .ZN(n785) );
  NOR2_X1 U867 ( .A1(n785), .A2(n784), .ZN(n828) );
  NAND2_X1 U868 ( .A1(G119), .A2(n872), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G131), .A2(n622), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U871 ( .A1(n867), .A2(G95), .ZN(n788) );
  XOR2_X1 U872 ( .A(KEYINPUT88), .B(n788), .Z(n789) );
  NOR2_X1 U873 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U874 ( .A1(G107), .A2(n625), .ZN(n791) );
  NAND2_X1 U875 ( .A1(n792), .A2(n791), .ZN(n855) );
  NAND2_X1 U876 ( .A1(G1991), .A2(n855), .ZN(n801) );
  NAND2_X1 U877 ( .A1(G129), .A2(n872), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G141), .A2(n622), .ZN(n793) );
  NAND2_X1 U879 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U880 ( .A1(n867), .A2(G105), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G117), .A2(n625), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n879) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n879), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n921) );
  NAND2_X1 U887 ( .A1(n828), .A2(n921), .ZN(n817) );
  XNOR2_X1 U888 ( .A(KEYINPUT37), .B(G2067), .ZN(n826) );
  NAND2_X1 U889 ( .A1(G104), .A2(n867), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G140), .A2(n622), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U892 ( .A(KEYINPUT34), .B(n804), .ZN(n809) );
  NAND2_X1 U893 ( .A1(G128), .A2(n872), .ZN(n806) );
  NAND2_X1 U894 ( .A1(G116), .A2(n625), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U896 ( .A(KEYINPUT35), .B(n807), .Z(n808) );
  NOR2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U898 ( .A(KEYINPUT36), .B(n810), .ZN(n864) );
  NOR2_X1 U899 ( .A1(n826), .A2(n864), .ZN(n934) );
  NAND2_X1 U900 ( .A1(n828), .A2(n934), .ZN(n825) );
  NAND2_X1 U901 ( .A1(n817), .A2(n825), .ZN(n811) );
  NOR2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U903 ( .A(n813), .B(KEYINPUT100), .ZN(n816) );
  XNOR2_X1 U904 ( .A(G1986), .B(G290), .ZN(n944) );
  NAND2_X1 U905 ( .A1(n828), .A2(n944), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT87), .B(n814), .Z(n815) );
  NAND2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n879), .ZN(n926) );
  INV_X1 U909 ( .A(n817), .ZN(n820) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n855), .ZN(n922) );
  NOR2_X1 U912 ( .A1(n818), .A2(n922), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n926), .A2(n821), .ZN(n822) );
  XOR2_X1 U915 ( .A(n822), .B(KEYINPUT101), .Z(n823) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n823), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n826), .A2(n864), .ZN(n936) );
  NAND2_X1 U919 ( .A1(n827), .A2(n936), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U922 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U924 ( .A(n833), .ZN(G223) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U926 ( .A(G661), .ZN(n834) );
  NOR2_X1 U927 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U928 ( .A(n836), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n838), .A2(n837), .ZN(G188) );
  XOR2_X1 U931 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  XNOR2_X1 U932 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  NOR2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  NAND2_X1 U937 ( .A1(n872), .A2(G124), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G100), .A2(n867), .ZN(n842) );
  NAND2_X1 U940 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U941 ( .A1(G136), .A2(n622), .ZN(n845) );
  NAND2_X1 U942 ( .A1(G112), .A2(n625), .ZN(n844) );
  NAND2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G162) );
  NAND2_X1 U945 ( .A1(G130), .A2(n872), .ZN(n849) );
  NAND2_X1 U946 ( .A1(G118), .A2(n625), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n854) );
  NAND2_X1 U948 ( .A1(G106), .A2(n867), .ZN(n851) );
  NAND2_X1 U949 ( .A1(G142), .A2(n622), .ZN(n850) );
  NAND2_X1 U950 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n852), .B(KEYINPUT45), .Z(n853) );
  NOR2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U954 ( .A(G162), .B(n857), .ZN(n866) );
  XOR2_X1 U955 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n859) );
  XNOR2_X1 U956 ( .A(G160), .B(KEYINPUT110), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U958 ( .A(n860), .B(KEYINPUT109), .Z(n862) );
  XOR2_X1 U959 ( .A(n923), .B(KEYINPUT46), .Z(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U961 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(n882) );
  NAND2_X1 U963 ( .A1(n867), .A2(G103), .ZN(n868) );
  XOR2_X1 U964 ( .A(KEYINPUT111), .B(n868), .Z(n870) );
  NAND2_X1 U965 ( .A1(n622), .A2(G139), .ZN(n869) );
  NAND2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT112), .B(n871), .ZN(n878) );
  NAND2_X1 U968 ( .A1(G127), .A2(n872), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G115), .A2(n625), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U971 ( .A(KEYINPUT113), .B(n875), .ZN(n876) );
  XNOR2_X1 U972 ( .A(KEYINPUT47), .B(n876), .ZN(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n916) );
  XNOR2_X1 U974 ( .A(n916), .B(n879), .ZN(n880) );
  XOR2_X1 U975 ( .A(G164), .B(n880), .Z(n881) );
  XNOR2_X1 U976 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U977 ( .A1(G37), .A2(n883), .ZN(G395) );
  XOR2_X1 U978 ( .A(n884), .B(G286), .Z(n886) );
  XOR2_X1 U979 ( .A(G301), .B(n948), .Z(n885) );
  XNOR2_X1 U980 ( .A(n886), .B(n885), .ZN(n887) );
  NOR2_X1 U981 ( .A1(G37), .A2(n887), .ZN(n888) );
  XOR2_X1 U982 ( .A(KEYINPUT115), .B(n888), .Z(G397) );
  XOR2_X1 U983 ( .A(G2096), .B(KEYINPUT43), .Z(n890) );
  XOR2_X1 U984 ( .A(n998), .B(G2678), .Z(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U986 ( .A(n891), .B(KEYINPUT106), .Z(n893) );
  XNOR2_X1 U987 ( .A(G2067), .B(G2090), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n898) );
  XNOR2_X1 U989 ( .A(KEYINPUT42), .B(n894), .ZN(n896) );
  XNOR2_X1 U990 ( .A(G2084), .B(G2078), .ZN(n895) );
  XNOR2_X1 U991 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(G227) );
  XOR2_X1 U993 ( .A(G2474), .B(G1956), .Z(n900) );
  XNOR2_X1 U994 ( .A(G1996), .B(G1991), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n901), .B(KEYINPUT107), .Z(n903) );
  XNOR2_X1 U997 ( .A(G1966), .B(G1981), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U999 ( .A(G1976), .B(G1971), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1986), .B(G1961), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1002 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT41), .B(KEYINPUT108), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(G229) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n910), .B(KEYINPUT116), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n911), .ZN(n912) );
  NOR2_X1 U1008 ( .A1(G401), .A2(n912), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .Z(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G303), .ZN(G166) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1015 ( .A(G164), .B(G2078), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n916), .B(KEYINPUT119), .ZN(n917) );
  XOR2_X1 U1017 ( .A(n917), .B(G2072), .Z(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT50), .ZN(n939) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n932) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT117), .B(n927), .Z(n928) );
  XNOR2_X1 U1026 ( .A(n928), .B(KEYINPUT51), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(KEYINPUT118), .ZN(n937) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT52), .B(n940), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n1013) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n1013), .ZN(n942) );
  NAND2_X1 U1036 ( .A1(n942), .A2(G29), .ZN(n1022) );
  INV_X1 U1037 ( .A(G16), .ZN(n992) );
  XOR2_X1 U1038 ( .A(n992), .B(KEYINPUT56), .Z(n967) );
  XOR2_X1 U1039 ( .A(G1961), .B(G171), .Z(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n956) );
  XOR2_X1 U1042 ( .A(G1971), .B(G303), .Z(n947) );
  XNOR2_X1 U1043 ( .A(n947), .B(KEYINPUT124), .ZN(n954) );
  XOR2_X1 U1044 ( .A(G299), .B(G1956), .Z(n950) );
  XNOR2_X1 U1045 ( .A(n948), .B(G1348), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n965) );
  XOR2_X1 U1050 ( .A(n957), .B(G1341), .Z(n963) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G168), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT123), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(KEYINPUT57), .B(n961), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n994) );
  XNOR2_X1 U1058 ( .A(KEYINPUT125), .B(G1961), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(n968), .B(G5), .ZN(n980) );
  XNOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n969), .B(G4), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(G1981), .B(G6), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(G20), .B(G1956), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1068 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G21), .ZN(n977) );
  NOR2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(KEYINPUT126), .B(n981), .ZN(n989) );
  XOR2_X1 U1073 ( .A(G1986), .B(G24), .Z(n985) );
  XNOR2_X1 U1074 ( .A(G1971), .B(G22), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT127), .B(n986), .Z(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n1020) );
  XNOR2_X1 U1084 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n995), .B(G34), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G2084), .B(n996), .ZN(n1012) );
  XNOR2_X1 U1087 ( .A(G2090), .B(G35), .ZN(n1010) );
  XOR2_X1 U1088 ( .A(G1991), .B(G25), .Z(n997) );
  NAND2_X1 U1089 ( .A1(n997), .A2(G28), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G2067), .B(G26), .ZN(n1000) );
  XOR2_X1 U1091 ( .A(G33), .B(n998), .Z(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1996), .B(G32), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G27), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT53), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(n1014), .B(n1013), .ZN(n1016) );
  INV_X1 U1102 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

