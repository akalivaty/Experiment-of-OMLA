//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT67), .Z(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT68), .B(new_n466), .C1(new_n464), .C2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT3), .B1(new_n464), .B2(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(G137), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n464), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n469), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n466), .B1(new_n471), .B2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n464), .B2(KEYINPUT69), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(G2105), .B1(new_n484), .B2(new_n470), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n476), .B1(new_n484), .B2(new_n470), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  AND2_X1   g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n475), .A2(new_n476), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n475), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n476), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n494), .A2(new_n497), .A3(new_n501), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT70), .B1(new_n507), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n507), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n522), .A2(G89), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(G51), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n528), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n512), .A2(new_n513), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n516), .B1(new_n541), .B2(new_n542), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G52), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n520), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n523), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n545), .A2(new_n549), .ZN(G171));
  AOI22_X1  g125(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n516), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n522), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n553));
  AND2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  AOI21_X1  g134(.A(new_n509), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n560));
  NOR3_X1   g135(.A1(new_n507), .A2(KEYINPUT70), .A3(G543), .ZN(new_n561));
  OAI211_X1 g136(.A(G65), .B(new_n513), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT76), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  NOR2_X1   g145(.A1(KEYINPUT6), .A2(G651), .ZN(new_n571));
  AND2_X1   g146(.A1(KEYINPUT6), .A2(G651), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(G543), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n518), .A2(new_n575), .A3(G543), .A4(new_n570), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n522), .A2(G91), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n568), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  INV_X1    g155(.A(G166), .ZN(G303));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n516), .B1(new_n539), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT77), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n522), .A2(G87), .B1(new_n520), .B2(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(new_n522), .A2(G86), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT79), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n539), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n512), .A2(KEYINPUT78), .A3(G61), .A4(new_n513), .ZN(new_n593));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n520), .A2(G48), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n522), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n516), .ZN(G290));
  NAND2_X1  g176(.A1(new_n522), .A2(G92), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT10), .Z(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n539), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n520), .A2(KEYINPUT80), .ZN(new_n607));
  INV_X1    g182(.A(G54), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n519), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n606), .A2(G651), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(new_n613), .B2(G171), .ZN(G321));
  MUX2_X1   g191(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g193(.A(new_n612), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g200(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n626));
  NOR3_X1   g201(.A1(new_n466), .A2(new_n464), .A3(G2105), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n487), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n485), .A2(G135), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n633), .A2(KEYINPUT82), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(KEYINPUT82), .B2(new_n633), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n631), .A2(new_n632), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(G2096), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n630), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT83), .Z(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n644), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2451), .B(G2454), .Z(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(new_n657), .A3(G14), .ZN(G401));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n662), .B2(new_n659), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(KEYINPUT86), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(KEYINPUT86), .B2(new_n665), .ZN(new_n667));
  INV_X1    g242(.A(new_n659), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n664), .A3(new_n661), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n660), .A2(new_n664), .A3(new_n662), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  AOI211_X1 g259(.A(new_n681), .B(new_n684), .C1(new_n676), .C2(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n691), .ZN(G229));
  MUX2_X1   g267(.A(G24), .B(G290), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1986), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(KEYINPUT91), .B2(KEYINPUT36), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT90), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n487), .A2(G119), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n485), .A2(G131), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n476), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT89), .Z(new_n704));
  OAI21_X1  g279(.A(new_n695), .B1(new_n697), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n697), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G23), .ZN(new_n708));
  INV_X1    g283(.A(G288), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(new_n707), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(G6), .A2(G16), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G305), .B2(new_n707), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n707), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n707), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n710), .A2(new_n711), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n712), .A2(new_n716), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n714), .A2(new_n715), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n722), .A2(KEYINPUT34), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(KEYINPUT34), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n706), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n727), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G19), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(new_n554), .B2(G16), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT92), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G32), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G105), .B2(new_n478), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n485), .A2(G141), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n487), .A2(G129), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n736), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT27), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1996), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n735), .A2(G26), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n485), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n487), .A2(G128), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n734), .A2(new_n747), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n735), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n735), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT29), .B(G2090), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n707), .A2(G21), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G168), .B2(new_n707), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G1966), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n619), .B2(G16), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n768), .B(new_n771), .C1(G1348), .C2(new_n773), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n773), .A2(G1348), .B1(new_n770), .B2(G1966), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT24), .B(G34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(new_n735), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT97), .Z(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n480), .B2(new_n735), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT99), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G28), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n735), .B1(new_n785), .B2(G28), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n784), .B1(new_n786), .B2(new_n787), .C1(new_n637), .C2(new_n735), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G2072), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n735), .A2(G33), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n465), .A2(new_n467), .A3(G127), .ZN(new_n792));
  INV_X1    g367(.A(G115), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(new_n464), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G2105), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT25), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n485), .B2(G139), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(G29), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n789), .B1(new_n790), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n775), .A2(new_n782), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(G171), .A2(new_n707), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G5), .B2(new_n707), .ZN(new_n805));
  INV_X1    g380(.A(G1961), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NOR2_X1   g383(.A1(G164), .A2(new_n735), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G27), .B2(new_n735), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n801), .A2(new_n790), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n811), .B2(new_n810), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n774), .A2(new_n803), .A3(new_n807), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n707), .A2(G20), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT23), .Z(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G299), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT101), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT100), .B(G1956), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NOR3_X1   g397(.A1(new_n764), .A2(new_n815), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n730), .A2(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  NAND2_X1  g400(.A1(new_n619), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(new_n516), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n522), .A2(G93), .B1(new_n520), .B2(G55), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n554), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT39), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT102), .B(G860), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT103), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n831), .A2(new_n835), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(G145));
  XOR2_X1   g415(.A(new_n757), .B(KEYINPUT105), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n800), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n702), .B(new_n628), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n485), .A2(new_n493), .B1(new_n503), .B2(new_n502), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n495), .B1(new_n484), .B2(new_n470), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n500), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n497), .A2(KEYINPUT104), .A3(new_n501), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n743), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n487), .A2(G130), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n476), .A2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G142), .B2(new_n485), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n851), .B(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n844), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n844), .A2(new_n857), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(new_n637), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G162), .ZN(new_n863));
  AOI21_X1  g438(.A(G37), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT106), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n860), .A2(KEYINPUT106), .A3(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g444(.A1(new_n619), .A2(G299), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n612), .A2(new_n568), .A3(new_n577), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n870), .A2(KEYINPUT41), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n873), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n832), .B(new_n622), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n870), .A2(new_n871), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(KEYINPUT108), .C1(new_n879), .C2(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(G166), .B(KEYINPUT109), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(G288), .B(G290), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(KEYINPUT42), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n887), .ZN(new_n891));
  OR3_X1    g466(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT42), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n883), .A3(new_n880), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G868), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n831), .A2(G868), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(G295));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n901), .A3(new_n899), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n613), .B1(new_n893), .B2(new_n895), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT110), .B1(new_n903), .B2(new_n898), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(G331));
  XNOR2_X1  g480(.A(G168), .B(G171), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n832), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(new_n881), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n878), .A2(new_n907), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n888), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n876), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n907), .A2(KEYINPUT41), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n888), .B(new_n913), .C1(new_n914), .C2(new_n881), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n908), .A2(new_n888), .A3(new_n909), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n912), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n919), .B2(new_n910), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n915), .A2(new_n912), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n922), .B2(new_n910), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n911), .A2(new_n912), .A3(new_n918), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n917), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(new_n925), .ZN(G397));
  NAND2_X1  g501(.A1(G303), .A2(G8), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n927), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G8), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n469), .A2(new_n477), .A3(G40), .A4(new_n479), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n505), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n934), .B2(KEYINPUT50), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n500), .B1(new_n475), .B2(new_n496), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n504), .B(new_n494), .C1(new_n937), .C2(KEYINPUT104), .ZN(new_n938));
  INV_X1    g513(.A(new_n849), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n936), .B(new_n933), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G2090), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n935), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n935), .A2(new_n940), .A3(KEYINPUT112), .A4(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(KEYINPUT45), .B(new_n933), .C1(new_n938), .C2(new_n939), .ZN(new_n947));
  INV_X1    g522(.A(new_n932), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n934), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n719), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(KEYINPUT111), .A3(new_n719), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n946), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n931), .B1(new_n956), .B2(KEYINPUT113), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n951), .A2(KEYINPUT111), .A3(new_n719), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT111), .B1(new_n951), .B2(new_n719), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n958), .B1(new_n961), .B2(new_n946), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n930), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT115), .B(G8), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n850), .A2(new_n933), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n948), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n709), .A2(G1976), .ZN(new_n968));
  INV_X1    g543(.A(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT52), .B1(G288), .B2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n971), .B1(KEYINPUT52), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n596), .A2(new_n587), .A3(new_n597), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(new_n976), .A3(G1981), .ZN(new_n977));
  INV_X1    g552(.A(G1981), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n589), .A2(new_n978), .A3(new_n596), .A4(new_n597), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n976), .B1(new_n975), .B2(G1981), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n974), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(G1981), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT116), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(KEYINPUT49), .A3(new_n979), .A4(new_n977), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(new_n967), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT45), .B1(new_n850), .B2(new_n933), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n948), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n935), .A2(new_n940), .A3(new_n780), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n964), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(G286), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n973), .A2(new_n986), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT63), .B1(new_n963), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n967), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n986), .A2(new_n969), .A3(new_n709), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n979), .B(KEYINPUT117), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n954), .A2(new_n955), .ZN(new_n1003));
  INV_X1    g578(.A(new_n946), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(KEYINPUT113), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n962), .A2(new_n1005), .A3(G8), .A4(new_n930), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n936), .B1(new_n850), .B2(new_n933), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n505), .A2(new_n936), .A3(new_n933), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n948), .A2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1007), .A2(new_n1009), .A3(G2090), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n719), .B2(new_n951), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n929), .B1(new_n1011), .B2(new_n964), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT63), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1006), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n973), .A2(new_n986), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1002), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1956), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n947), .A2(new_n950), .A3(new_n948), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n577), .B(new_n1024), .C1(new_n566), .C2(new_n567), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1019), .A2(new_n1021), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n935), .A2(new_n940), .ZN(new_n1031));
  INV_X1    g606(.A(G1348), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n1034));
  AND4_X1   g609(.A1(new_n933), .A2(new_n948), .A3(new_n850), .A4(new_n762), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1348), .B1(new_n935), .B2(new_n940), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n1038), .B2(new_n1035), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n619), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1026), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1025), .B(new_n1041), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1042), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1030), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1034), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1038), .A2(new_n1035), .A3(KEYINPUT119), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT60), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1037), .A2(new_n1048), .A3(new_n1039), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n619), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT61), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(KEYINPUT122), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1043), .B2(new_n1029), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(KEYINPUT122), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n951), .B2(G1996), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT58), .B(G1341), .Z(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n965), .B2(new_n932), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n951), .A2(new_n1056), .A3(G1996), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n554), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AND2_X1   g637(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1063));
  NOR2_X1   g638(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1050), .A2(new_n1055), .A3(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT122), .B(new_n1051), .C1(new_n1043), .C2(new_n1029), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n554), .B(new_n1063), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1069));
  OAI211_X1 g644(.A(KEYINPUT60), .B(new_n612), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1044), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(G168), .A2(new_n964), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n995), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n931), .B1(new_n991), .B2(new_n992), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT51), .B1(new_n1077), .B2(new_n1074), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n964), .B1(new_n991), .B2(new_n992), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1076), .A2(new_n1078), .B1(G286), .B2(new_n1079), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n965), .A2(new_n949), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n811), .A2(KEYINPUT53), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n947), .A2(new_n948), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1082), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n988), .A2(new_n1084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(KEYINPUT125), .A3(new_n948), .A4(new_n947), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n947), .A2(new_n950), .A3(new_n811), .A4(new_n948), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT124), .B(KEYINPUT53), .Z(new_n1092));
  AOI21_X1  g667(.A(G171), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1031), .A2(new_n806), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1090), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1083), .A2(new_n948), .A3(new_n1085), .A4(new_n989), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1081), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1080), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n973), .A2(new_n986), .A3(new_n1012), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1088), .A2(new_n1090), .A3(new_n1096), .A4(new_n1094), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1097), .A2(new_n1094), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1093), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1104), .B(KEYINPUT54), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1101), .A2(new_n1006), .A3(new_n1102), .A4(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n998), .B(new_n1017), .C1(new_n1073), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1102), .A2(new_n1006), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT54), .B1(new_n1106), .B2(new_n1105), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(G171), .B2(new_n1103), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1114), .A2(new_n1080), .A3(new_n1100), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1050), .A2(new_n1055), .A3(new_n1066), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1071), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1112), .B(new_n1115), .C1(new_n1117), .C2(new_n1044), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(KEYINPUT126), .A3(new_n998), .A4(new_n1017), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1080), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1099), .B1(new_n1120), .B2(KEYINPUT62), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1112), .B(new_n1121), .C1(KEYINPUT62), .C2(new_n1120), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1111), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1083), .A2(new_n932), .ZN(new_n1124));
  INV_X1    g699(.A(G1996), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n743), .B(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n757), .B(new_n762), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n702), .B(new_n697), .Z(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G290), .B(G1986), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1124), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT46), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1124), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1127), .A2(new_n744), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT47), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n702), .A2(new_n697), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n757), .A2(G2067), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1136), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1136), .A2(G1986), .A3(G290), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(KEYINPUT48), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(KEYINPUT48), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1146), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1141), .A2(new_n1142), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1133), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g728(.A1(new_n916), .A2(new_n920), .ZN(new_n1155));
  NOR4_X1   g729(.A1(G401), .A2(new_n460), .A3(G227), .A4(G229), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n1155), .A2(new_n868), .A3(new_n1156), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


