//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT74), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT74), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n190), .B1(G472), .B2(G902), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G210), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n195), .B(KEYINPUT27), .Z(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G101), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n198), .B(KEYINPUT72), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT70), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G146), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT64), .A2(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT64), .A2(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(new_n209), .B2(G146), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT64), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT64), .A2(G143), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n211), .A2(KEYINPUT66), .A3(G146), .A4(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n203), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT64), .B(G143), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n220), .B2(new_n218), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n203), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  AOI21_X1  g040(.A(G146), .B1(new_n211), .B2(new_n212), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n226), .B(new_n223), .C1(new_n227), .C2(new_n219), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NOR3_X1   g043(.A1(new_n207), .A2(new_n208), .A3(new_n218), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n213), .B1(new_n230), .B2(new_n206), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT67), .A3(new_n203), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT11), .B1(new_n234), .B2(G134), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(KEYINPUT68), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G137), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT11), .A2(G134), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n237), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AOI211_X1 g062(.A(new_n245), .B(new_n246), .C1(new_n237), .C2(new_n242), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n201), .B1(new_n233), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n247), .A2(new_n245), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n246), .B1(new_n237), .B2(new_n242), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(new_n249), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT66), .B1(new_n218), .B2(G143), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n220), .B2(new_n218), .ZN(new_n258));
  AOI211_X1 g072(.A(new_n216), .B(new_n202), .C1(new_n258), .C2(new_n213), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT67), .B1(new_n231), .B2(new_n203), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(new_n261), .A3(KEYINPUT70), .A4(new_n229), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n231), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(G143), .B2(new_n218), .ZN(new_n269));
  OAI22_X1  g083(.A1(new_n227), .A2(new_n219), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(G134), .B1(new_n238), .B2(new_n240), .ZN(new_n272));
  INV_X1    g086(.A(new_n236), .ZN(new_n273));
  OAI21_X1  g087(.A(G131), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g090(.A(KEYINPUT71), .B(G131), .C1(new_n272), .C2(new_n273), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(new_n247), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n263), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT2), .B(G113), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G116), .B(G119), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g098(.A(G116), .B(G119), .Z(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n280), .A2(KEYINPUT73), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n287), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(new_n279), .C1(new_n233), .C2(new_n251), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n291));
  INV_X1    g105(.A(new_n279), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n252), .B2(new_n262), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n289), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT28), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n290), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n200), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n256), .A2(new_n261), .A3(new_n229), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n300), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n287), .B(new_n301), .C1(new_n293), .C2(KEYINPUT30), .ZN(new_n302));
  INV_X1    g116(.A(new_n198), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n290), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT31), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n302), .A2(new_n306), .A3(new_n290), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n192), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT32), .ZN(new_n310));
  INV_X1    g124(.A(new_n298), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n295), .B2(KEYINPUT28), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n305), .B(new_n307), .C1(new_n312), .C2(new_n200), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n192), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n290), .A2(new_n317), .A3(new_n297), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n279), .B1(new_n233), .B2(new_n251), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n287), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n297), .B1(new_n320), .B2(new_n290), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n298), .A2(KEYINPUT75), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n198), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G902), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(KEYINPUT76), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n328));
  AOI211_X1 g142(.A(new_n328), .B(G902), .C1(new_n323), .C2(new_n325), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n296), .A2(new_n298), .A3(new_n200), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n302), .A2(new_n290), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT29), .B1(new_n332), .B2(new_n198), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  AOI211_X1 g148(.A(KEYINPUT77), .B(new_n187), .C1(new_n330), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n336));
  INV_X1    g150(.A(new_n318), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n289), .B1(new_n300), .B2(new_n279), .ZN(new_n338));
  INV_X1    g152(.A(new_n290), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT28), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n317), .B1(new_n290), .B2(new_n297), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n325), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n188), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n328), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n326), .A2(KEYINPUT76), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n311), .B(new_n199), .C1(new_n295), .C2(KEYINPUT28), .ZN(new_n347));
  INV_X1    g161(.A(new_n333), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n345), .B(new_n346), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n336), .B1(new_n349), .B2(G472), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n316), .B1(new_n335), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT78), .B(G217), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(G234), .B2(new_n188), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(G125), .B(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n218), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  INV_X1    g174(.A(G125), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT16), .ZN(new_n363));
  OR3_X1    g177(.A1(new_n361), .A2(KEYINPUT16), .A3(G140), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n364), .A3(G146), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n363), .A2(new_n364), .A3(new_n367), .A4(G146), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n369));
  INV_X1    g183(.A(G119), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n370), .B2(G128), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n268), .A2(KEYINPUT23), .A3(G119), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(new_n372), .C1(G119), .C2(new_n268), .ZN(new_n373));
  XNOR2_X1  g187(.A(G119), .B(G128), .ZN(new_n374));
  XOR2_X1   g188(.A(KEYINPUT24), .B(G110), .Z(new_n375));
  OAI22_X1  g189(.A1(new_n373), .A2(G110), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n358), .A2(new_n366), .A3(new_n368), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n364), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n218), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n365), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n373), .A2(G110), .B1(new_n374), .B2(new_n375), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n384), .B(new_n385), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n382), .A3(new_n386), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n188), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT25), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n388), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n389), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n354), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n389), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n353), .A2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n394), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  INV_X1    g218(.A(G104), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT19), .B1(new_n355), .B2(KEYINPUT91), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT91), .A2(new_n360), .A3(new_n362), .A4(KEYINPUT19), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n218), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n366), .A3(new_n368), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT92), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n193), .A2(new_n194), .A3(G214), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n209), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n193), .A2(new_n194), .A3(G143), .A4(G214), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G131), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n246), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n409), .A2(new_n419), .A3(new_n366), .A4(new_n368), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n411), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  OR2_X1    g235(.A1(new_n355), .A2(new_n218), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n356), .A2(new_n357), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT80), .B1(new_n355), .B2(new_n218), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT18), .A2(G131), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n415), .A2(new_n426), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n425), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n406), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n406), .B(KEYINPUT93), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n418), .A2(KEYINPUT17), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n379), .B(new_n365), .C1(new_n416), .C2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n430), .B(new_n432), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT94), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(G475), .A2(G902), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT94), .ZN(new_n440));
  INV_X1    g254(.A(new_n429), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n441), .A2(new_n427), .B1(new_n358), .B2(new_n422), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n410), .A2(KEYINPUT92), .B1(new_n416), .B2(new_n417), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n420), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n440), .B(new_n436), .C1(new_n444), .C2(new_n406), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n439), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT20), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n448), .B(new_n439), .C1(new_n431), .C2(new_n437), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G475), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n433), .A2(new_n435), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n442), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n436), .B1(new_n453), .B2(new_n406), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n451), .B1(new_n454), .B2(new_n188), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G478), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(KEYINPUT15), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n207), .A2(new_n208), .A3(new_n268), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT95), .B1(new_n461), .B2(KEYINPUT13), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n205), .A2(G128), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n461), .B2(KEYINPUT13), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n211), .A2(G128), .A3(new_n212), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT13), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G134), .ZN(new_n470));
  INV_X1    g284(.A(G134), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n465), .B(new_n471), .C1(G128), .C2(new_n205), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n473));
  INV_X1    g287(.A(G107), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT82), .A2(G107), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G122), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G116), .ZN(new_n479));
  INV_X1    g293(.A(G116), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n477), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n470), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n480), .A2(G122), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n481), .B1(new_n488), .B2(KEYINPUT14), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT96), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n491), .B(new_n481), .C1(new_n488), .C2(KEYINPUT14), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n481), .A2(KEYINPUT14), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G107), .ZN(new_n495));
  OAI21_X1  g309(.A(G134), .B1(new_n461), .B2(new_n463), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n484), .B1(new_n496), .B2(new_n472), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT9), .B(G234), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n352), .A2(new_n499), .A3(G953), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n487), .A2(KEYINPUT97), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n500), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n495), .A2(new_n497), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n485), .B1(new_n469), .B2(G134), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n470), .A2(new_n486), .B1(new_n497), .B2(new_n495), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT97), .B1(new_n507), .B2(new_n500), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n188), .B(new_n460), .C1(new_n506), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT99), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n487), .A2(new_n498), .A3(new_n500), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT97), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n505), .A3(new_n501), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT99), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n188), .A4(new_n460), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n194), .A2(G952), .ZN(new_n518));
  INV_X1    g332(.A(G234), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n518), .B1(new_n519), .B2(new_n193), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n188), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n188), .B1(new_n506), .B2(new_n508), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT98), .B1(new_n526), .B2(new_n459), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n528));
  AOI211_X1 g342(.A(new_n528), .B(new_n460), .C1(new_n514), .C2(new_n188), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n517), .B(new_n525), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT100), .B1(new_n457), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n455), .B1(new_n447), .B2(new_n449), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n459), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n528), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n526), .A2(KEYINPUT98), .A3(new_n459), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n534), .A2(new_n535), .B1(new_n510), .B2(new_n516), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT100), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n532), .A2(new_n536), .A3(new_n537), .A4(new_n525), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT3), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n475), .A2(new_n540), .A3(G104), .A4(new_n476), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n474), .B2(G104), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n474), .A2(G104), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G101), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n544), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n545), .A2(KEYINPUT83), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n546), .A2(KEYINPUT4), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(KEYINPUT4), .A3(new_n548), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n287), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT87), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n546), .A2(KEYINPUT4), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n547), .A2(new_n548), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT87), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n287), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT5), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n370), .A3(G116), .ZN(new_n561));
  OAI211_X1 g375(.A(G113), .B(new_n561), .C1(new_n285), .C2(new_n560), .ZN(new_n562));
  AOI21_X1  g376(.A(G104), .B1(new_n475), .B2(new_n476), .ZN(new_n563));
  INV_X1    g377(.A(new_n543), .ZN(new_n564));
  OAI21_X1  g378(.A(G101), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n565), .A3(new_n284), .A4(new_n546), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT88), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(G110), .B(G122), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n568), .B1(new_n558), .B2(new_n553), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n571), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT6), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n577), .A3(new_n572), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n271), .A2(G125), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(G125), .B2(new_n233), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n194), .A2(G224), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G210), .B1(G237), .B2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT90), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n581), .A2(KEYINPUT7), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n562), .A2(new_n284), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n565), .A2(new_n546), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(KEYINPUT89), .A3(new_n566), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n571), .B(KEYINPUT8), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n593), .B(new_n594), .C1(KEYINPUT89), .C2(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n595), .B1(new_n580), .B2(new_n588), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n597), .B2(new_n575), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n583), .A2(new_n587), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n587), .B1(new_n583), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G214), .B1(G237), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G221), .B1(new_n499), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(G469), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n188), .ZN(new_n608));
  XNOR2_X1  g422(.A(G110), .B(G140), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n194), .A2(G227), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n565), .A2(KEYINPUT10), .A3(new_n546), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n271), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G128), .B1(new_n227), .B2(new_n264), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n258), .A3(new_n213), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n591), .B1(new_n615), .B2(new_n267), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(KEYINPUT10), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT84), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n549), .A2(new_n551), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n233), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n261), .A2(new_n556), .A3(KEYINPUT84), .A4(new_n229), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n256), .B(new_n617), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  INV_X1    g437(.A(new_n617), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n251), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n611), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n623), .A2(new_n251), .A3(new_n624), .ZN(new_n627));
  INV_X1    g441(.A(new_n611), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n267), .A2(new_n591), .A3(new_n270), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n615), .A2(new_n267), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n591), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT12), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(KEYINPUT85), .A3(new_n632), .A4(new_n256), .ZN(new_n633));
  INV_X1    g447(.A(new_n629), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n256), .B1(new_n634), .B2(new_n616), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n627), .A2(new_n628), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n626), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n608), .B1(new_n640), .B2(new_n607), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n638), .A2(new_n633), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n611), .B1(new_n622), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n627), .A2(KEYINPUT86), .A3(new_n628), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n623), .A2(new_n624), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n256), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(KEYINPUT86), .B1(new_n627), .B2(new_n628), .ZN(new_n648));
  OAI211_X1 g462(.A(G469), .B(new_n643), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n606), .B1(new_n641), .B2(new_n649), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n539), .A2(new_n604), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n351), .A2(new_n403), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n583), .A2(new_n584), .A3(new_n598), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n584), .B1(new_n583), .B2(new_n598), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n525), .B(new_n602), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n505), .A2(KEYINPUT33), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n514), .A2(new_n658), .B1(new_n659), .B2(new_n511), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(G478), .A3(new_n188), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n526), .A2(new_n458), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n457), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n654), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n583), .A2(new_n598), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n585), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n583), .A2(new_n584), .A3(new_n598), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n603), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n532), .B1(new_n662), .B2(new_n661), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(KEYINPUT101), .A4(new_n525), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n187), .B1(new_n313), .B2(new_n188), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n628), .B1(new_n646), .B2(new_n627), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n622), .A2(new_n642), .A3(new_n611), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n607), .B(new_n188), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n608), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n649), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n678), .A2(new_n403), .A3(new_n605), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n305), .A2(new_n307), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n289), .B1(new_n263), .B2(new_n279), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n339), .B1(new_n681), .B2(KEYINPUT73), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n297), .B1(new_n682), .B2(new_n294), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n199), .B1(new_n683), .B2(new_n311), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n680), .A2(new_n684), .B1(new_n191), .B2(new_n189), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n673), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n672), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT34), .B(G104), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G6));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n438), .A2(new_n448), .A3(new_n445), .A4(new_n439), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n455), .B1(new_n447), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n517), .B1(new_n527), .B2(new_n529), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n690), .B1(new_n657), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n669), .A2(KEYINPUT102), .A3(new_n525), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n686), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT35), .B(G107), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G9));
  NOR2_X1   g515(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n383), .B(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n397), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n394), .A2(new_n705), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n539), .A2(new_n604), .A3(new_n650), .A4(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n673), .A2(new_n685), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT37), .B(G110), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G12));
  NAND2_X1  g525(.A1(new_n669), .A2(new_n706), .ZN(new_n712));
  INV_X1    g526(.A(G900), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n522), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n520), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n712), .A2(new_n694), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n351), .A2(new_n650), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  INV_X1    g533(.A(new_n650), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n715), .B(new_n721), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n601), .B(KEYINPUT38), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n532), .A2(new_n536), .A3(new_n603), .ZN(new_n726));
  INV_X1    g540(.A(new_n706), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n724), .A2(new_n725), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n199), .B1(new_n338), .B2(new_n339), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n304), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n731), .B2(G902), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n316), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n220), .ZN(G45));
  NAND3_X1  g550(.A1(new_n457), .A2(new_n663), .A3(new_n715), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n712), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n351), .A2(new_n650), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(new_n676), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n640), .A2(new_n607), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n605), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n665), .B2(new_n671), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n351), .A2(new_n403), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(KEYINPUT104), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n746), .B(new_n748), .ZN(G15));
  AOI21_X1  g563(.A(new_n744), .B1(new_n695), .B2(new_n697), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n351), .A2(new_n403), .A3(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G116), .ZN(G18));
  INV_X1    g566(.A(new_n539), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n744), .A3(new_n712), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n351), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n313), .A2(new_n188), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(G472), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n192), .B(KEYINPUT105), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n342), .A2(new_n199), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n305), .A2(KEYINPUT106), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n307), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT106), .B1(new_n305), .B2(new_n760), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n744), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n667), .A2(new_n668), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n726), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n524), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n766), .A2(new_n399), .A3(new_n767), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n738), .A3(new_n767), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  INV_X1    g588(.A(new_n737), .ZN(new_n775));
  INV_X1    g589(.A(new_n600), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n583), .A2(new_n587), .A3(new_n598), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n602), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n720), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n351), .A2(new_n403), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n349), .A2(G472), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT77), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n349), .A2(new_n336), .A3(G472), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n310), .A2(new_n787), .A3(new_n315), .ZN(new_n788));
  INV_X1    g602(.A(new_n315), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n314), .B1(new_n313), .B2(new_n192), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT107), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n720), .A2(new_n778), .A3(new_n737), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n793), .A2(KEYINPUT42), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n792), .A2(new_n794), .A3(new_n399), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n782), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G131), .ZN(G33));
  NOR2_X1   g611(.A1(new_n694), .A2(new_n716), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n351), .A2(new_n403), .A3(new_n798), .A4(new_n779), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NAND2_X1  g614(.A1(new_n532), .A2(new_n663), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT43), .Z(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n708), .A3(new_n727), .ZN(new_n804));
  OR3_X1    g618(.A1(new_n804), .A2(KEYINPUT109), .A3(KEYINPUT44), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n647), .A2(new_n648), .ZN(new_n806));
  INV_X1    g620(.A(new_n643), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n808), .A2(KEYINPUT45), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(KEYINPUT45), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(G469), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT46), .B1(new_n811), .B2(new_n677), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n741), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n606), .B(new_n722), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n804), .B2(KEYINPUT44), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n778), .B(KEYINPUT108), .Z(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n804), .B2(KEYINPUT44), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n805), .A2(new_n815), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  INV_X1    g634(.A(new_n351), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n778), .A2(new_n737), .A3(new_n403), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n813), .A2(new_n814), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT47), .B1(new_n826), .B2(new_n605), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT47), .ZN(new_n828));
  AOI211_X1 g642(.A(new_n828), .B(new_n606), .C1(new_n813), .C2(new_n814), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n824), .B(new_n825), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  NOR2_X1   g645(.A1(new_n827), .A2(new_n829), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n743), .A2(new_n606), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n832), .A2(KEYINPUT117), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n803), .A2(new_n520), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n765), .A2(new_n394), .A3(new_n398), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n817), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT117), .B1(new_n832), .B2(new_n833), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n744), .A2(new_n778), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n803), .A2(new_n520), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n765), .A2(new_n727), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n403), .A2(new_n521), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n733), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n532), .A2(new_n662), .A3(new_n661), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n602), .B1(KEYINPUT116), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n837), .A2(new_n725), .A3(new_n767), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n853));
  OAI221_X1 g667(.A(new_n846), .B1(new_n848), .B2(new_n849), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n832), .A2(KEYINPUT115), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n833), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n832), .A2(KEYINPUT115), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n839), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT51), .B1(new_n860), .B2(new_n855), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n792), .A2(new_n399), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n844), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n863), .B(KEYINPUT48), .Z(new_n864));
  NAND4_X1  g678(.A1(new_n835), .A2(new_n836), .A3(new_n669), .A4(new_n767), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n865), .B(new_n518), .C1(new_n664), .C2(new_n848), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n856), .A2(new_n861), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n718), .A2(new_n773), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n706), .A2(new_n716), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n650), .A2(new_n726), .A3(new_n768), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n316), .B2(new_n732), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n720), .B1(new_n786), .B2(new_n316), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n872), .B2(new_n738), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n868), .A2(new_n873), .A3(KEYINPUT52), .ZN(new_n874));
  INV_X1    g688(.A(new_n871), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n718), .A2(new_n739), .A3(new_n875), .A4(new_n773), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n692), .A2(new_n536), .A3(new_n715), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n601), .A4(new_n602), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT112), .B1(new_n778), .B2(new_n880), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n727), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n351), .A2(new_n650), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n845), .A2(new_n793), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n799), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n746), .A2(new_n751), .A3(new_n771), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n525), .B(new_n602), .C1(new_n599), .C2(new_n600), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n532), .A2(new_n693), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n664), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n707), .A2(new_n708), .B1(new_n686), .B2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n652), .A2(new_n893), .A3(new_n755), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n796), .A2(new_n888), .A3(new_n889), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n799), .A2(new_n886), .A3(new_n887), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n782), .B2(new_n795), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n746), .A2(new_n751), .A3(new_n771), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n652), .A2(new_n893), .A3(new_n755), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT113), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n879), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT52), .B1(new_n868), .B2(new_n873), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n876), .A2(new_n877), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT53), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT114), .B1(new_n910), .B2(new_n895), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n905), .B1(new_n874), .B2(new_n878), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n796), .A2(new_n888), .A3(new_n889), .A4(new_n894), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT114), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT54), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n904), .A2(new_n905), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n867), .A2(new_n907), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(G952), .B2(G953), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n399), .A2(new_n602), .A3(new_n605), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n801), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT49), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n743), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT111), .Z(new_n925));
  INV_X1    g739(.A(new_n733), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n743), .A2(new_n923), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n925), .A2(new_n926), .A3(new_n725), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n920), .A2(new_n928), .ZN(G75));
  AND3_X1   g743(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n914), .B1(new_n912), .B2(new_n913), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n895), .A2(new_n896), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n899), .A2(KEYINPUT113), .A3(new_n902), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n935), .B2(new_n879), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n188), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT56), .B1(new_n938), .B2(G210), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n576), .A2(new_n578), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(new_n582), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT55), .Z(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n194), .A2(G952), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n939), .A2(KEYINPUT118), .A3(new_n943), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT118), .B1(new_n939), .B2(new_n943), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G51));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT54), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n952), .B1(new_n930), .B2(new_n931), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n953), .B2(new_n936), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT119), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT54), .B1(new_n932), .B2(new_n936), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n608), .B(KEYINPUT57), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n626), .A2(new_n639), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT120), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n962), .A3(new_n958), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n937), .A2(new_n188), .A3(new_n811), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n945), .B1(new_n964), .B2(new_n965), .ZN(G54));
  NAND3_X1  g780(.A1(new_n938), .A2(KEYINPUT58), .A3(G475), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n438), .A2(new_n445), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n945), .ZN(G60));
  NAND2_X1  g785(.A1(G478), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT59), .Z(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n907), .B2(new_n918), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n946), .B1(new_n974), .B2(new_n660), .ZN(new_n975));
  INV_X1    g789(.A(new_n973), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n957), .A2(new_n660), .A3(new_n976), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(KEYINPUT121), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G63));
  XNOR2_X1  g794(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n981), .B(new_n982), .Z(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n932), .B2(new_n936), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n945), .B1(new_n984), .B2(new_n395), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n986));
  INV_X1    g800(.A(new_n984), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n703), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n984), .A2(KEYINPUT123), .A3(new_n704), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g806(.A(KEYINPUT61), .B(new_n985), .C1(new_n988), .C2(new_n989), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(G66));
  INV_X1    g808(.A(G224), .ZN(new_n995));
  OAI21_X1  g809(.A(G953), .B1(new_n523), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n902), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n940), .B1(G898), .B2(new_n194), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT124), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n997), .B(new_n999), .ZN(G69));
  OAI21_X1  g814(.A(new_n301), .B1(new_n293), .B2(KEYINPUT30), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n407), .A2(new_n408), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n815), .A2(new_n768), .A3(new_n726), .A4(new_n862), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT126), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n830), .A2(new_n819), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n868), .A2(new_n739), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n1008), .A2(new_n799), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1006), .A2(new_n1007), .A3(new_n796), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1004), .B1(new_n1010), .B2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n735), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT62), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1008), .A2(new_n1014), .A3(new_n735), .ZN(new_n1015));
  INV_X1    g829(.A(new_n723), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n778), .B1(new_n664), .B2(new_n891), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1016), .A2(new_n351), .A3(new_n403), .A4(new_n1017), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1007), .A2(new_n1013), .A3(new_n1015), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(KEYINPUT125), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n830), .A2(new_n819), .A3(new_n1018), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT125), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1021), .A2(new_n1022), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1023));
  AOI21_X1  g837(.A(G953), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1003), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1011), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT127), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1028), .B(new_n1011), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1027), .A2(new_n1031), .A3(new_n1029), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(G72));
  NAND2_X1  g849(.A1(G472), .A2(G902), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1036), .B(KEYINPUT63), .Z(new_n1037));
  NAND2_X1  g851(.A1(new_n332), .A2(new_n198), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n304), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1010), .A2(new_n198), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1040), .A2(new_n1038), .A3(new_n304), .A4(new_n902), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n198), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1042));
  OAI221_X1 g856(.A(new_n946), .B1(new_n1037), .B2(new_n1039), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1039), .A2(new_n1037), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1043), .B1(new_n906), .B2(new_n1044), .ZN(G57));
endmodule


