//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n461), .A2(G2105), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(G101), .ZN(new_n469));
  AND4_X1   g044(.A1(new_n467), .A2(new_n465), .A3(G101), .A4(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n462), .A2(new_n464), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n462), .A2(new_n464), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n476), .A2(new_n465), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  AND3_X1   g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n465), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  AND2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT6), .A2(G651), .ZN(new_n498));
  OAI21_X1  g073(.A(G543), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G50), .ZN(new_n500));
  OR3_X1    g075(.A1(new_n499), .A2(KEYINPUT70), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT70), .B1(new_n499), .B2(new_n500), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n504), .A2(KEYINPUT71), .A3(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(KEYINPUT71), .B1(new_n504), .B2(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n497), .A2(new_n498), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n507), .A2(G62), .A3(new_n509), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n515), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n507), .A2(new_n509), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n511), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT73), .B(G89), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n499), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  AND4_X1   g105(.A1(new_n524), .A2(new_n525), .A3(new_n528), .A4(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n516), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n522), .A2(G81), .B1(G43), .B2(new_n529), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n521), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n541), .A2(new_n542), .A3(G651), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n542), .B1(new_n541), .B2(G651), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n507), .A2(G65), .A3(new_n509), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n516), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n507), .A2(G91), .A3(new_n509), .A4(new_n512), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n529), .B(new_n559), .C1(KEYINPUT75), .C2(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n561), .B(new_n562), .C1(new_n499), .C2(new_n558), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n557), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  NAND4_X1  g142(.A1(new_n524), .A2(new_n525), .A3(new_n528), .A4(new_n530), .ZN(G286));
  AND2_X1   g143(.A1(new_n517), .A2(new_n518), .ZN(new_n569));
  OAI221_X1 g144(.A(new_n503), .B1(new_n513), .B2(new_n514), .C1(new_n516), .C2(new_n569), .ZN(G303));
  OAI21_X1  g145(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n507), .A2(G87), .A3(new_n509), .A4(new_n512), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n529), .A2(G49), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n507), .A2(G61), .A3(new_n509), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n516), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n507), .A2(G86), .A3(new_n509), .A4(new_n512), .ZN(new_n580));
  OAI211_X1 g155(.A(G48), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n581));
  XOR2_X1   g156(.A(new_n581), .B(KEYINPUT76), .Z(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n522), .A2(G85), .B1(G47), .B2(new_n529), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G60), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n521), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n513), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n522), .A2(G92), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n529), .A2(G54), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n516), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n590), .B1(G868), .B2(new_n600), .ZN(G284));
  XNOR2_X1  g176(.A(G284), .B(KEYINPUT78), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n565), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G868), .B2(new_n565), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n600), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n547), .ZN(G323));
  XNOR2_X1  g185(.A(KEYINPUT79), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  NAND2_X1  g187(.A1(new_n477), .A2(G2104), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT80), .B(G2100), .Z(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n477), .A2(G135), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n482), .A2(G123), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n465), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G1341), .B(G1348), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT83), .Z(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT84), .Z(G401));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT85), .Z(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT17), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  INV_X1    g227(.A(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n646), .B2(new_n648), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT86), .Z(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n647), .B2(new_n649), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n652), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT91), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT33), .B(G1976), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n680), .A2(G22), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n680), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G6), .A2(G16), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n582), .A2(new_n580), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(new_n578), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n692), .B1(new_n694), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n686), .A2(new_n687), .A3(new_n691), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n477), .A2(G131), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT88), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n465), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n482), .A2(G119), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G25), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT35), .B(G1991), .Z(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT89), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(G16), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT90), .B(G1986), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n699), .A2(new_n700), .A3(new_n711), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT36), .Z(new_n716));
  NOR2_X1   g291(.A1(G29), .A2(G35), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G162), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n719));
  INV_X1    g294(.A(G2090), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n718), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n680), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n680), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G1961), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n547), .A2(new_n680), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n680), .B2(G19), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n726), .B1(new_n727), .B2(new_n729), .C1(G1961), .C2(new_n724), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n680), .A2(G20), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT23), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n565), .B2(new_n680), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1956), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G4), .A2(G16), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n600), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT92), .B(G1348), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G168), .A2(new_n680), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n680), .B2(G21), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT94), .Z(new_n745));
  NOR2_X1   g320(.A1(G29), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n477), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n482), .A2(G129), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n468), .A2(G105), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  NAND4_X1  g326(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT30), .B(G28), .ZN(new_n758));
  INV_X1    g333(.A(G29), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n623), .B2(new_n759), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n759), .A2(G26), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT28), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n477), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n482), .A2(G128), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n465), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n765), .B1(new_n770), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2067), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n775), .B2(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(KEYINPUT24), .B2(new_n775), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n468), .A2(new_n467), .A3(G101), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(KEYINPUT68), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n473), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n493), .B2(G125), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n466), .B(new_n781), .C1(new_n783), .C2(new_n465), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(new_n759), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n763), .B(new_n773), .C1(new_n774), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n759), .A2(G33), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  AOI22_X1  g364(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(new_n477), .ZN(new_n791));
  INV_X1    g366(.A(G139), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(new_n790), .B2(new_n465), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(new_n759), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n795), .A2(G2072), .B1(new_n774), .B2(new_n785), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G2072), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n757), .A2(new_n786), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G164), .A2(G29), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G27), .B2(G29), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT95), .B(G2078), .Z(new_n801));
  AOI22_X1  g376(.A1(new_n742), .A2(new_n743), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n745), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n731), .A2(new_n736), .A3(new_n740), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n716), .A2(new_n805), .ZN(G311));
  OR2_X1    g381(.A1(new_n716), .A2(new_n805), .ZN(G150));
  NAND4_X1  g382(.A1(new_n507), .A2(G93), .A3(new_n509), .A4(new_n512), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT98), .B(G55), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n499), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n507), .A2(G67), .A3(new_n509), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n516), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G860), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT99), .B1(new_n810), .B2(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(new_n546), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n541), .A2(G651), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT74), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(new_n543), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n825), .A2(new_n538), .A3(new_n819), .A4(new_n820), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n600), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n830));
  XOR2_X1   g405(.A(new_n829), .B(new_n830), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n815), .B1(new_n832), .B2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n817), .B1(new_n833), .B2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n623), .B(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(G162), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n492), .A2(new_n495), .ZN(new_n838));
  INV_X1    g413(.A(new_n490), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n770), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT100), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n770), .B(G164), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n753), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(new_n845), .A3(new_n754), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n793), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n707), .B(new_n614), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n477), .A2(G142), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n482), .A2(G130), .ZN(new_n852));
  OR2_X1    g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n850), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n843), .A2(new_n752), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n843), .A2(new_n752), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n793), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n849), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n847), .A2(new_n848), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n794), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n850), .B(new_n855), .Z(new_n866));
  NAND4_X1  g441(.A1(new_n865), .A2(new_n866), .A3(new_n862), .A4(new_n859), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n856), .B1(new_n849), .B2(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n837), .B1(new_n863), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(KEYINPUT102), .B(new_n837), .C1(new_n863), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n861), .A2(new_n837), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g453(.A(new_n608), .B(KEYINPUT103), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n827), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n600), .A2(new_n565), .ZN(new_n881));
  OAI21_X1  g456(.A(G299), .B1(new_n596), .B2(new_n599), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g460(.A(KEYINPUT41), .B1(new_n881), .B2(new_n882), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n884), .B1(new_n887), .B2(new_n880), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n682), .A2(new_n588), .A3(new_n584), .ZN(new_n889));
  NAND2_X1  g464(.A1(G290), .A2(G288), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G166), .B(G305), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G166), .B(new_n694), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n897), .A2(KEYINPUT104), .A3(new_n890), .A4(new_n889), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT42), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n896), .A2(new_n898), .A3(KEYINPUT105), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT105), .B1(new_n896), .B2(new_n898), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n902), .B2(KEYINPUT42), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n888), .B(new_n903), .Z(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G868), .B2(new_n814), .ZN(G295));
  OAI21_X1  g481(.A(new_n905), .B1(G868), .B2(new_n814), .ZN(G331));
  NAND3_X1  g482(.A1(new_n822), .A2(new_n826), .A3(G301), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(G301), .B1(new_n822), .B2(new_n826), .ZN(new_n910));
  OAI21_X1  g485(.A(G286), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n827), .A2(G171), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(G168), .A3(new_n908), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n913), .A3(new_n883), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT106), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n887), .B1(new_n911), .B2(new_n913), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n902), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n911), .A2(new_n913), .ZN(new_n918));
  INV_X1    g493(.A(new_n887), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n900), .A2(new_n901), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT106), .A4(new_n914), .ZN(new_n922));
  INV_X1    g497(.A(G37), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n917), .A2(new_n922), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n925), .A2(KEYINPUT107), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT43), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT44), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n925), .A2(new_n927), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(KEYINPUT63), .ZN(new_n936));
  NAND3_X1  g511(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n937));
  OAI21_X1  g512(.A(G8), .B1(new_n515), .B2(new_n519), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT55), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT109), .B1(G160), .B2(G40), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n471), .A2(new_n474), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n840), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n840), .A2(new_n950), .A3(new_n947), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n943), .B1(new_n784), .B2(new_n944), .ZN(new_n955));
  NAND3_X1  g530(.A1(G160), .A2(KEYINPUT109), .A3(G40), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n838), .B2(new_n839), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n952), .A2(new_n720), .B1(new_n959), .B2(new_n690), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n941), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n937), .A2(new_n940), .ZN(new_n963));
  INV_X1    g538(.A(new_n959), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(G1971), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n957), .B2(new_n950), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT113), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n946), .A2(new_n967), .A3(new_n951), .A4(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G2090), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n963), .B(G8), .C1(new_n965), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1981), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n579), .A2(new_n972), .A3(new_n580), .A4(new_n582), .ZN(new_n973));
  OAI21_X1  g548(.A(G1981), .B1(new_n693), .B2(new_n578), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT49), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n973), .A2(new_n974), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(KEYINPUT49), .B1(new_n973), .B2(new_n974), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n982), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  NOR2_X1   g561(.A1(G288), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT52), .B1(new_n982), .B2(new_n987), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n962), .A2(new_n971), .A3(new_n984), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT115), .B(G2084), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n994), .A2(new_n967), .A3(new_n968), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(G164), .B2(G1384), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n948), .B2(new_n953), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n955), .A2(new_n956), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n743), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n961), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G168), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n936), .B1(new_n993), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n984), .A2(new_n992), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n965), .B2(new_n970), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n941), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1003), .A2(new_n936), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1005), .A2(new_n971), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n984), .A2(new_n986), .A3(new_n682), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n973), .ZN(new_n1012));
  INV_X1    g587(.A(new_n971), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1012), .A2(new_n985), .B1(new_n1013), .B2(new_n1005), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n952), .A2(G1956), .B1(new_n959), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n564), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n554), .A2(new_n555), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G651), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT57), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(KEYINPUT57), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1022), .B(KEYINPUT57), .C1(new_n556), .C2(new_n564), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1018), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n1029));
  INV_X1    g604(.A(G1956), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n964), .A2(new_n1016), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1027), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT61), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1027), .A2(KEYINPUT118), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1025), .A2(new_n1036), .A3(new_n1026), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n1038), .B2(new_n1031), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1018), .A2(new_n1040), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1033), .A2(KEYINPUT61), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n981), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n959), .B2(G1996), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT120), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n1046), .C1(new_n959), .C2(G1996), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n546), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n969), .A2(KEYINPUT117), .ZN(new_n1054));
  INV_X1    g629(.A(G1348), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n994), .A2(new_n1056), .A3(new_n967), .A4(new_n968), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n946), .A2(new_n772), .A3(new_n957), .ZN(new_n1059));
  AND2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n600), .ZN(new_n1062));
  INV_X1    g637(.A(new_n600), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1058), .A2(new_n1063), .A3(new_n1059), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT60), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1044), .A2(new_n1053), .A3(new_n1062), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1042), .B1(new_n1063), .B2(new_n1060), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1033), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1961), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1054), .A2(new_n1071), .A3(new_n1057), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n959), .B2(G2078), .ZN(new_n1074));
  NOR4_X1   g649(.A1(new_n784), .A2(new_n1073), .A3(new_n944), .A4(G2078), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n954), .A2(new_n958), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(G171), .B(KEYINPUT54), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OR4_X1    g654(.A1(KEYINPUT123), .A2(new_n999), .A3(new_n1000), .A4(G2078), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n1081));
  NOR3_X1   g656(.A1(G164), .A2(G1384), .A3(new_n953), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n946), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT123), .B1(new_n1084), .B2(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(KEYINPUT53), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1079), .B1(new_n1087), .B2(new_n1078), .ZN(new_n1088));
  AND4_X1   g663(.A1(new_n962), .A2(new_n971), .A3(new_n984), .A4(new_n992), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G286), .A2(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n996), .B2(new_n1001), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1091), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1002), .A2(new_n1094), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1097), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n968), .A2(new_n951), .A3(new_n955), .A4(new_n956), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT113), .B1(new_n948), .B2(KEYINPUT50), .ZN(new_n1101));
  INV_X1    g676(.A(new_n995), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1966), .B1(new_n1083), .B2(new_n946), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1099), .B1(new_n1105), .B2(new_n1091), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1093), .B1(new_n1098), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT122), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1091), .A3(new_n1099), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1001), .B1(new_n969), .B2(new_n1102), .ZN(new_n1110));
  OAI211_X1 g685(.A(G8), .B(new_n1097), .C1(new_n1110), .C2(G286), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1093), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1090), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1015), .B1(new_n1070), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1108), .A2(new_n1117), .A3(new_n1114), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1089), .A2(G171), .A3(new_n1087), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(KEYINPUT124), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1113), .B1(new_n1112), .B2(new_n1093), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT122), .B(new_n1092), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT62), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT125), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(KEYINPUT62), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT124), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1116), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1000), .A2(new_n954), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G1996), .A3(new_n752), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1131), .A2(KEYINPUT110), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(KEYINPUT110), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n770), .B(new_n772), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n753), .B2(G1996), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1130), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT111), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n707), .B(new_n709), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT112), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1130), .A3(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(G290), .A2(G1986), .ZN(new_n1144));
  NOR2_X1   g719(.A1(G290), .A2(G1986), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1130), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1129), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1138), .A2(new_n702), .A3(new_n706), .A4(new_n709), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1151), .B1(G2067), .B2(new_n770), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1130), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1134), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1130), .B1(new_n1154), .B2(new_n752), .ZN(new_n1155));
  INV_X1    g730(.A(G1996), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1130), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(KEYINPUT46), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT47), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1145), .A2(new_n1130), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1143), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1153), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1149), .A2(new_n1150), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n1168));
  NOR3_X1   g743(.A1(new_n1121), .A2(new_n1122), .A3(KEYINPUT62), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1089), .A2(G171), .A3(new_n1087), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1171), .A2(new_n1120), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1147), .B1(new_n1172), .B2(new_n1116), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT126), .B1(new_n1173), .B2(new_n1165), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1167), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g750(.A1(G227), .A2(new_n459), .ZN(new_n1177));
  NAND3_X1  g751(.A1(new_n678), .A2(new_n1177), .A3(new_n643), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1178), .B1(new_n874), .B2(new_n876), .ZN(new_n1179));
  AND3_X1   g753(.A1(new_n1179), .A2(new_n932), .A3(KEYINPUT127), .ZN(new_n1180));
  AOI21_X1  g754(.A(KEYINPUT127), .B1(new_n1179), .B2(new_n932), .ZN(new_n1181));
  NOR2_X1   g755(.A1(new_n1180), .A2(new_n1181), .ZN(G308));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n932), .ZN(G225));
endmodule


