

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U551 ( .A1(n682), .A2(n793), .ZN(n727) );
  BUF_X2 U552 ( .A(n877), .Z(n516) );
  XOR2_X1 U553 ( .A(KEYINPUT17), .B(n517), .Z(n877) );
  INV_X1 U554 ( .A(n727), .ZN(n712) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n648) );
  NOR2_X1 U557 ( .A1(n745), .A2(n717), .ZN(n719) );
  NOR2_X1 U558 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U559 ( .A1(G651), .A2(n633), .ZN(n638) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n536), .Z(n639) );
  NAND2_X1 U561 ( .A1(G138), .A2(n516), .ZN(n519) );
  INV_X1 U562 ( .A(G2105), .ZN(n524) );
  AND2_X1 U563 ( .A1(n524), .A2(G2104), .ZN(n878) );
  NAND2_X1 U564 ( .A1(G102), .A2(n878), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n519), .A2(n518), .ZN(n521) );
  INV_X1 U566 ( .A(KEYINPUT90), .ZN(n520) );
  XNOR2_X1 U567 ( .A(n521), .B(n520), .ZN(n523) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U569 ( .A1(n881), .A2(G114), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n523), .A2(n522), .ZN(n527) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n524), .ZN(n882) );
  NAND2_X1 U572 ( .A1(G126), .A2(n882), .ZN(n525) );
  XNOR2_X1 U573 ( .A(KEYINPUT89), .B(n525), .ZN(n526) );
  NOR2_X1 U574 ( .A1(n527), .A2(n526), .ZN(G164) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(KEYINPUT65), .Z(n529) );
  NAND2_X1 U576 ( .A1(G101), .A2(n878), .ZN(n528) );
  XOR2_X1 U577 ( .A(n529), .B(n528), .Z(n677) );
  NAND2_X1 U578 ( .A1(n516), .A2(G137), .ZN(n530) );
  XNOR2_X1 U579 ( .A(n530), .B(KEYINPUT66), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G113), .A2(n881), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U582 ( .A(KEYINPUT67), .B(n533), .ZN(n681) );
  NAND2_X1 U583 ( .A1(G125), .A2(n882), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT64), .ZN(n678) );
  AND2_X1 U585 ( .A1(n681), .A2(n678), .ZN(n535) );
  AND2_X1 U586 ( .A1(n677), .A2(n535), .ZN(G160) );
  XOR2_X1 U587 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U588 ( .A1(G47), .A2(n638), .ZN(n538) );
  INV_X1 U589 ( .A(G651), .ZN(n539) );
  NOR2_X1 U590 ( .A1(G543), .A2(n539), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G60), .A2(n639), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G85), .A2(n648), .ZN(n541) );
  NOR2_X1 U594 ( .A1(n633), .A2(n539), .ZN(n642) );
  NAND2_X1 U595 ( .A1(G72), .A2(n642), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U597 ( .A1(n543), .A2(n542), .ZN(G290) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G69), .ZN(G235) );
  INV_X1 U601 ( .A(G108), .ZN(G238) );
  INV_X1 U602 ( .A(G120), .ZN(G236) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(G88), .A2(n648), .ZN(n545) );
  NAND2_X1 U605 ( .A1(G75), .A2(n642), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G50), .A2(n638), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G62), .A2(n639), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U610 ( .A1(n549), .A2(n548), .ZN(G166) );
  NAND2_X1 U611 ( .A1(G52), .A2(n638), .ZN(n551) );
  NAND2_X1 U612 ( .A1(G64), .A2(n639), .ZN(n550) );
  NAND2_X1 U613 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U614 ( .A(KEYINPUT68), .B(n552), .ZN(n558) );
  NAND2_X1 U615 ( .A1(n642), .A2(G77), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT69), .B(n553), .Z(n555) );
  NAND2_X1 U617 ( .A1(n648), .A2(G90), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U620 ( .A1(n558), .A2(n557), .ZN(G171) );
  INV_X1 U621 ( .A(G166), .ZN(G303) );
  NAND2_X1 U622 ( .A1(G51), .A2(n638), .ZN(n560) );
  NAND2_X1 U623 ( .A1(G63), .A2(n639), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(KEYINPUT6), .B(n561), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n648), .A2(G89), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G76), .A2(n642), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(n565), .B(KEYINPUT5), .Z(n566) );
  NOR2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U632 ( .A(KEYINPUT7), .B(n568), .Z(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT77), .B(n569), .Z(G168) );
  XOR2_X1 U634 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U637 ( .A(G223), .ZN(n828) );
  NAND2_X1 U638 ( .A1(n828), .A2(G567), .ZN(n571) );
  XOR2_X1 U639 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U640 ( .A1(n639), .A2(G56), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT14), .B(n572), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G81), .A2(n648), .ZN(n573) );
  XNOR2_X1 U643 ( .A(n573), .B(KEYINPUT12), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT72), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G68), .A2(n642), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(n577), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT73), .ZN(n582) );
  NAND2_X1 U650 ( .A1(G43), .A2(n638), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n1008) );
  INV_X1 U652 ( .A(G860), .ZN(n603) );
  OR2_X1 U653 ( .A1(n1008), .A2(n603), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G301), .A2(G868), .ZN(n583) );
  XNOR2_X1 U656 ( .A(n583), .B(KEYINPUT74), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G54), .A2(n638), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(KEYINPUT76), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G92), .A2(n648), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G79), .A2(n642), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G66), .A2(n639), .ZN(n587) );
  XNOR2_X1 U663 ( .A(KEYINPUT75), .B(n587), .ZN(n588) );
  NOR2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U665 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X2 U666 ( .A(KEYINPUT15), .B(n592), .ZN(n992) );
  OR2_X1 U667 ( .A1(G868), .A2(n992), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G53), .A2(n638), .ZN(n596) );
  NAND2_X1 U670 ( .A1(G65), .A2(n639), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G91), .A2(n648), .ZN(n598) );
  NAND2_X1 U673 ( .A1(G78), .A2(n642), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n600), .A2(n599), .ZN(n996) );
  XOR2_X1 U676 ( .A(n996), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U677 ( .A1(G299), .A2(G868), .ZN(n602) );
  INV_X1 U678 ( .A(G868), .ZN(n659) );
  NOR2_X1 U679 ( .A1(G286), .A2(n659), .ZN(n601) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(G297) );
  NAND2_X1 U681 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n604), .A2(n992), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U684 ( .A1(G868), .A2(n1008), .ZN(n608) );
  NAND2_X1 U685 ( .A1(G868), .A2(n992), .ZN(n606) );
  NOR2_X1 U686 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G111), .A2(n881), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G99), .A2(n878), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U691 ( .A(KEYINPUT78), .B(n611), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G123), .A2(n882), .ZN(n612) );
  XNOR2_X1 U693 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n516), .A2(G135), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n972) );
  XNOR2_X1 U697 ( .A(n972), .B(G2096), .ZN(n618) );
  INV_X1 U698 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U700 ( .A1(G55), .A2(n638), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G67), .A2(n639), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n642), .A2(G80), .ZN(n621) );
  XOR2_X1 U704 ( .A(KEYINPUT80), .B(n621), .Z(n622) );
  NOR2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n648), .A2(G93), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n660) );
  XNOR2_X1 U708 ( .A(n1008), .B(KEYINPUT79), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n992), .A2(G559), .ZN(n626) );
  XOR2_X1 U710 ( .A(n627), .B(n626), .Z(n657) );
  NOR2_X1 U711 ( .A1(n657), .A2(G860), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n628), .B(KEYINPUT81), .ZN(n629) );
  XNOR2_X1 U713 ( .A(n660), .B(n629), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G49), .A2(n638), .ZN(n631) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U716 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U717 ( .A(KEYINPUT82), .B(n632), .Z(n635) );
  NAND2_X1 U718 ( .A1(n633), .A2(G87), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U720 ( .A1(n636), .A2(n639), .ZN(n637) );
  XNOR2_X1 U721 ( .A(n637), .B(KEYINPUT83), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G48), .A2(n638), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n647) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(KEYINPUT85), .Z(n644) );
  NAND2_X1 U726 ( .A1(G73), .A2(n642), .ZN(n643) );
  XNOR2_X1 U727 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U728 ( .A(KEYINPUT84), .B(n645), .Z(n646) );
  NOR2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n648), .A2(G86), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G305) );
  XNOR2_X1 U732 ( .A(G299), .B(G288), .ZN(n651) );
  XNOR2_X1 U733 ( .A(n651), .B(n660), .ZN(n652) );
  XOR2_X1 U734 ( .A(n652), .B(KEYINPUT86), .Z(n654) );
  XNOR2_X1 U735 ( .A(G166), .B(KEYINPUT19), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U737 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(G305), .ZN(n895) );
  XOR2_X1 U739 ( .A(n657), .B(n895), .Z(n658) );
  NAND2_X1 U740 ( .A1(n658), .A2(G868), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U742 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(KEYINPUT87), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n664), .B(KEYINPUT20), .ZN(n665) );
  NAND2_X1 U746 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U750 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U753 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G96), .A2(n670), .ZN(n915) );
  NAND2_X1 U755 ( .A1(n915), .A2(G2106), .ZN(n675) );
  NOR2_X1 U756 ( .A1(G236), .A2(G238), .ZN(n672) );
  NOR2_X1 U757 ( .A1(G235), .A2(G237), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U759 ( .A(KEYINPUT88), .B(n673), .ZN(n916) );
  NAND2_X1 U760 ( .A1(n916), .A2(G567), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n832) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U763 ( .A1(n832), .A2(n676), .ZN(n831) );
  NAND2_X1 U764 ( .A1(n831), .A2(G36), .ZN(G176) );
  XOR2_X1 U765 ( .A(G1981), .B(G305), .Z(n1011) );
  AND2_X1 U766 ( .A1(n677), .A2(G40), .ZN(n679) );
  AND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n792) );
  INV_X1 U769 ( .A(n792), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n793) );
  NAND2_X1 U771 ( .A1(G8), .A2(n727), .ZN(n768) );
  NOR2_X1 U772 ( .A1(G288), .A2(G1976), .ZN(n683) );
  XNOR2_X1 U773 ( .A(n683), .B(KEYINPUT103), .ZN(n1003) );
  NOR2_X1 U774 ( .A1(n768), .A2(n1003), .ZN(n684) );
  NAND2_X1 U775 ( .A1(KEYINPUT33), .A2(n684), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n1011), .A2(n685), .ZN(n762) );
  INV_X1 U777 ( .A(n1008), .ZN(n696) );
  AND2_X1 U778 ( .A1(n696), .A2(n992), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n712), .ZN(n686) );
  XNOR2_X1 U780 ( .A(n686), .B(KEYINPUT26), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n727), .A2(G1341), .ZN(n687) );
  XNOR2_X1 U782 ( .A(n687), .B(KEYINPUT96), .ZN(n688) );
  AND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n697) );
  NAND2_X1 U784 ( .A1(n690), .A2(n697), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n712), .A2(G1348), .ZN(n692) );
  NOR2_X1 U786 ( .A1(G2067), .A2(n727), .ZN(n691) );
  NOR2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U788 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n695), .B(KEYINPUT97), .ZN(n700) );
  AND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U791 ( .A1(n992), .A2(n698), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n706) );
  NAND2_X1 U793 ( .A1(n712), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n701), .B(KEYINPUT27), .ZN(n703) );
  INV_X1 U795 ( .A(G1956), .ZN(n939) );
  NOR2_X1 U796 ( .A1(n712), .A2(n939), .ZN(n702) );
  NOR2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n996), .A2(n707), .ZN(n704) );
  XOR2_X1 U799 ( .A(KEYINPUT98), .B(n704), .Z(n705) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U801 ( .A1(n996), .A2(n707), .ZN(n708) );
  XNOR2_X1 U802 ( .A(n708), .B(KEYINPUT28), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n711), .B(KEYINPUT29), .ZN(n740) );
  NAND2_X1 U805 ( .A1(G1961), .A2(n727), .ZN(n714) );
  XOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .Z(n918) );
  NAND2_X1 U807 ( .A1(n712), .A2(n918), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n721) );
  OR2_X1 U809 ( .A1(n721), .A2(G301), .ZN(n739) );
  AND2_X1 U810 ( .A1(n739), .A2(G286), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n740), .A2(n715), .ZN(n736) );
  INV_X1 U812 ( .A(G286), .ZN(n726) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n768), .ZN(n745) );
  NOR2_X1 U814 ( .A1(n727), .A2(G2084), .ZN(n716) );
  XNOR2_X1 U815 ( .A(n716), .B(KEYINPUT95), .ZN(n743) );
  NAND2_X1 U816 ( .A1(G8), .A2(n743), .ZN(n717) );
  XNOR2_X1 U817 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n718) );
  XNOR2_X1 U818 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U819 ( .A1(n720), .A2(G168), .ZN(n724) );
  NAND2_X1 U820 ( .A1(G301), .A2(n721), .ZN(n722) );
  XOR2_X1 U821 ( .A(KEYINPUT100), .B(n722), .Z(n723) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n725), .Z(n741) );
  NOR2_X1 U823 ( .A1(n726), .A2(n741), .ZN(n734) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n727), .ZN(n728) );
  XOR2_X1 U825 ( .A(KEYINPUT101), .B(n728), .Z(n730) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n768), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U828 ( .A(n731), .B(KEYINPUT102), .ZN(n732) );
  AND2_X1 U829 ( .A1(n732), .A2(G303), .ZN(n733) );
  NOR2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U832 ( .A1(n737), .A2(G8), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n742) );
  AND2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n748) );
  INV_X1 U836 ( .A(n743), .ZN(n744) );
  AND2_X1 U837 ( .A1(G8), .A2(n744), .ZN(n746) );
  OR2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n765) );
  INV_X1 U841 ( .A(n1003), .ZN(n753) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n751) );
  XNOR2_X1 U843 ( .A(KEYINPUT104), .B(n751), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n755) );
  INV_X1 U845 ( .A(KEYINPUT33), .ZN(n754) );
  AND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n765), .A2(n756), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  INV_X1 U849 ( .A(n1002), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n757), .A2(n768), .ZN(n758) );
  OR2_X1 U851 ( .A1(KEYINPUT33), .A2(n758), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n774) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U855 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n766), .A2(n768), .ZN(n772) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XNOR2_X1 U859 ( .A(KEYINPUT24), .B(n767), .ZN(n770) );
  INV_X1 U860 ( .A(n768), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U862 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U864 ( .A(n775), .B(KEYINPUT105), .ZN(n808) );
  NAND2_X1 U865 ( .A1(G107), .A2(n881), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G95), .A2(n878), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G131), .A2(n516), .ZN(n779) );
  NAND2_X1 U869 ( .A1(G119), .A2(n882), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n864) );
  NAND2_X1 U872 ( .A1(n864), .A2(G1991), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G117), .A2(n881), .ZN(n783) );
  NAND2_X1 U874 ( .A1(G129), .A2(n882), .ZN(n782) );
  NAND2_X1 U875 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n878), .A2(G105), .ZN(n784) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n516), .A2(G141), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n861) );
  NAND2_X1 U881 ( .A1(G1996), .A2(n861), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U883 ( .A(n791), .B(KEYINPUT93), .ZN(n968) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n823) );
  XOR2_X1 U885 ( .A(n823), .B(KEYINPUT94), .Z(n794) );
  NOR2_X1 U886 ( .A1(n968), .A2(n794), .ZN(n815) );
  NAND2_X1 U887 ( .A1(G140), .A2(n516), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G104), .A2(n878), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT34), .B(n797), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G116), .A2(n881), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G128), .A2(n882), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U894 ( .A(n800), .B(KEYINPUT35), .Z(n801) );
  NOR2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U896 ( .A(KEYINPUT36), .B(n803), .Z(n804) );
  XNOR2_X1 U897 ( .A(KEYINPUT91), .B(n804), .ZN(n891) );
  XNOR2_X1 U898 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NOR2_X1 U899 ( .A1(n891), .A2(n821), .ZN(n805) );
  XNOR2_X1 U900 ( .A(n805), .B(KEYINPUT92), .ZN(n971) );
  NAND2_X1 U901 ( .A1(n823), .A2(n971), .ZN(n818) );
  INV_X1 U902 ( .A(n818), .ZN(n806) );
  NOR2_X1 U903 ( .A1(n815), .A2(n806), .ZN(n807) );
  AND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U905 ( .A(n809), .B(KEYINPUT106), .ZN(n811) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U907 ( .A1(n998), .A2(n823), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n861), .ZN(n812) );
  XOR2_X1 U910 ( .A(KEYINPUT107), .B(n812), .Z(n978) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n864), .ZN(n973) );
  NOR2_X1 U913 ( .A1(n813), .A2(n973), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n978), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT108), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n821), .A2(n891), .ZN(n988) );
  NAND2_X1 U920 ( .A1(n822), .A2(n988), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U929 ( .A(n832), .ZN(G319) );
  XOR2_X1 U930 ( .A(G2474), .B(G1981), .Z(n834) );
  XNOR2_X1 U931 ( .A(G1986), .B(G1971), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n835), .B(KEYINPUT112), .Z(n837) );
  XNOR2_X1 U934 ( .A(G1991), .B(G1996), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U936 ( .A(G1976), .B(G1956), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1966), .B(G1961), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G229) );
  XOR2_X1 U942 ( .A(KEYINPUT43), .B(G2678), .Z(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U945 ( .A(KEYINPUT42), .B(G2090), .Z(n847) );
  XNOR2_X1 U946 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U948 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2096), .B(G2100), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n853) );
  XOR2_X1 U951 ( .A(G2078), .B(G2084), .Z(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G227) );
  NAND2_X1 U953 ( .A1(G124), .A2(n882), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n881), .A2(G112), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U957 ( .A1(G136), .A2(n516), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G100), .A2(n878), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U960 ( .A1(n860), .A2(n859), .ZN(G162) );
  XNOR2_X1 U961 ( .A(n861), .B(G162), .ZN(n863) );
  XNOR2_X1 U962 ( .A(G160), .B(G164), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n893) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT115), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n876) );
  NAND2_X1 U967 ( .A1(G118), .A2(n881), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G130), .A2(n882), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n874) );
  NAND2_X1 U970 ( .A1(G142), .A2(n516), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G106), .A2(n878), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U973 ( .A(KEYINPUT45), .B(n871), .Z(n872) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(n872), .ZN(n873) );
  NOR2_X1 U975 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n876), .B(n875), .Z(n889) );
  NAND2_X1 U977 ( .A1(G139), .A2(n516), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n982) );
  XNOR2_X1 U985 ( .A(n972), .B(n982), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U989 ( .A1(G37), .A2(n894), .ZN(G395) );
  XOR2_X1 U990 ( .A(n895), .B(G286), .Z(n897) );
  XNOR2_X1 U991 ( .A(G171), .B(n992), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U993 ( .A(n898), .B(n1008), .Z(n899) );
  NOR2_X1 U994 ( .A1(G37), .A2(n899), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2430), .B(G2451), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2446), .B(G2427), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U998 ( .A(G2438), .B(KEYINPUT109), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2443), .B(G2454), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1001 ( .A(n904), .B(G2435), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G1341), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n909), .A2(G14), .ZN(n917) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n917), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  XOR2_X1 U1012 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(G325) );
  INV_X1 U1016 ( .A(G325), .ZN(G261) );
  INV_X1 U1017 ( .A(n917), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G2090), .B(G35), .Z(n932) );
  XNOR2_X1 U1019 ( .A(G1996), .B(G32), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(n918), .B(G27), .ZN(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(n921), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(G2067), .B(G26), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1025 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1027 ( .A(G1991), .B(G25), .Z(n926) );
  NAND2_X1 U1028 ( .A1(n926), .A2(G28), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n929), .B(KEYINPUT53), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n930), .B(KEYINPUT119), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(G34), .B(G2084), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(n936), .B(KEYINPUT120), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(G29), .A2(n937), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(KEYINPUT55), .B(n938), .ZN(n1023) );
  XOR2_X1 U1039 ( .A(G1961), .B(G5), .Z(n950) );
  XNOR2_X1 U1040 ( .A(G20), .B(n939), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1042 ( .A(n940), .B(G4), .ZN(n941) );
  NAND2_X1 U1043 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1046 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(n945), .B(KEYINPUT123), .ZN(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n948), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(G1966), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(G21), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT125), .B(n954), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(n955), .B(KEYINPUT58), .ZN(n961) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n959) );
  XNOR2_X1 U1058 ( .A(G1971), .B(G22), .ZN(n957) );
  XNOR2_X1 U1059 ( .A(G23), .B(G1976), .ZN(n956) );
  NOR2_X1 U1060 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1061 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1062 ( .A(n961), .B(n960), .Z(n962) );
  NOR2_X1 U1063 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1064 ( .A(KEYINPUT61), .B(n964), .ZN(n966) );
  INV_X1 U1065 ( .A(G16), .ZN(n965) );
  NAND2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(n967), .A2(G11), .ZN(n1021) );
  XNOR2_X1 U1068 ( .A(G160), .B(G2084), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT117), .B(n976), .ZN(n981) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT51), .B(n979), .Z(n980) );
  NAND2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1078 ( .A(G2072), .B(n982), .Z(n984) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n985), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(n990), .B(KEYINPUT52), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n991), .A2(G29), .ZN(n1019) );
  XNOR2_X1 U1086 ( .A(G16), .B(KEYINPUT56), .ZN(n1017) );
  XOR2_X1 U1087 ( .A(n992), .B(G1348), .Z(n994) );
  XOR2_X1 U1088 ( .A(G171), .B(G1961), .Z(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G166), .ZN(n995) );
  XNOR2_X1 U1091 ( .A(n995), .B(KEYINPUT122), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n996), .B(G1956), .ZN(n997) );
  XNOR2_X1 U1093 ( .A(n997), .B(KEYINPUT121), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(G1341), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G168), .ZN(n1012) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(n1013), .B(KEYINPUT57), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

